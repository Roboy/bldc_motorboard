// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Sep 18 2019 23:28:45

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    output USBPU;
    output PIN_9;
    input PIN_8;
    input PIN_7;
    inout PIN_6;
    inout PIN_5;
    inout PIN_4;
    output PIN_3;
    output PIN_24;
    output PIN_23;
    output PIN_22;
    input PIN_21;
    input PIN_20;
    output PIN_2;
    input PIN_19;
    input PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    input PIN_13;
    input PIN_12;
    inout PIN_11;
    inout PIN_10;
    output PIN_1;
    output LED;
    input CLK;

    wire N__70064;
    wire N__70063;
    wire N__70062;
    wire N__70055;
    wire N__70054;
    wire N__70053;
    wire N__70046;
    wire N__70045;
    wire N__70044;
    wire N__70037;
    wire N__70036;
    wire N__70035;
    wire N__70028;
    wire N__70027;
    wire N__70026;
    wire N__70019;
    wire N__70018;
    wire N__70017;
    wire N__70010;
    wire N__70009;
    wire N__70008;
    wire N__70001;
    wire N__70000;
    wire N__69999;
    wire N__69992;
    wire N__69991;
    wire N__69990;
    wire N__69983;
    wire N__69982;
    wire N__69981;
    wire N__69974;
    wire N__69973;
    wire N__69972;
    wire N__69965;
    wire N__69964;
    wire N__69963;
    wire N__69956;
    wire N__69955;
    wire N__69954;
    wire N__69947;
    wire N__69946;
    wire N__69945;
    wire N__69938;
    wire N__69937;
    wire N__69936;
    wire N__69929;
    wire N__69928;
    wire N__69927;
    wire N__69920;
    wire N__69919;
    wire N__69918;
    wire N__69911;
    wire N__69910;
    wire N__69909;
    wire N__69902;
    wire N__69901;
    wire N__69900;
    wire N__69883;
    wire N__69882;
    wire N__69881;
    wire N__69880;
    wire N__69879;
    wire N__69878;
    wire N__69877;
    wire N__69876;
    wire N__69873;
    wire N__69872;
    wire N__69871;
    wire N__69868;
    wire N__69867;
    wire N__69866;
    wire N__69865;
    wire N__69864;
    wire N__69861;
    wire N__69860;
    wire N__69857;
    wire N__69854;
    wire N__69851;
    wire N__69848;
    wire N__69847;
    wire N__69846;
    wire N__69845;
    wire N__69844;
    wire N__69841;
    wire N__69840;
    wire N__69839;
    wire N__69836;
    wire N__69833;
    wire N__69830;
    wire N__69827;
    wire N__69824;
    wire N__69821;
    wire N__69818;
    wire N__69815;
    wire N__69810;
    wire N__69807;
    wire N__69806;
    wire N__69803;
    wire N__69802;
    wire N__69801;
    wire N__69798;
    wire N__69795;
    wire N__69794;
    wire N__69791;
    wire N__69784;
    wire N__69781;
    wire N__69778;
    wire N__69777;
    wire N__69774;
    wire N__69771;
    wire N__69766;
    wire N__69761;
    wire N__69758;
    wire N__69751;
    wire N__69750;
    wire N__69747;
    wire N__69744;
    wire N__69741;
    wire N__69736;
    wire N__69731;
    wire N__69730;
    wire N__69727;
    wire N__69720;
    wire N__69717;
    wire N__69716;
    wire N__69713;
    wire N__69710;
    wire N__69703;
    wire N__69698;
    wire N__69697;
    wire N__69696;
    wire N__69695;
    wire N__69692;
    wire N__69687;
    wire N__69680;
    wire N__69677;
    wire N__69674;
    wire N__69669;
    wire N__69666;
    wire N__69663;
    wire N__69656;
    wire N__69649;
    wire N__69646;
    wire N__69641;
    wire N__69638;
    wire N__69633;
    wire N__69630;
    wire N__69625;
    wire N__69616;
    wire N__69613;
    wire N__69608;
    wire N__69605;
    wire N__69602;
    wire N__69595;
    wire N__69594;
    wire N__69591;
    wire N__69588;
    wire N__69585;
    wire N__69584;
    wire N__69581;
    wire N__69578;
    wire N__69575;
    wire N__69568;
    wire N__69567;
    wire N__69566;
    wire N__69565;
    wire N__69564;
    wire N__69563;
    wire N__69562;
    wire N__69561;
    wire N__69560;
    wire N__69559;
    wire N__69558;
    wire N__69557;
    wire N__69556;
    wire N__69555;
    wire N__69552;
    wire N__69549;
    wire N__69548;
    wire N__69545;
    wire N__69542;
    wire N__69539;
    wire N__69538;
    wire N__69537;
    wire N__69534;
    wire N__69529;
    wire N__69526;
    wire N__69521;
    wire N__69518;
    wire N__69513;
    wire N__69510;
    wire N__69507;
    wire N__69504;
    wire N__69503;
    wire N__69502;
    wire N__69497;
    wire N__69494;
    wire N__69493;
    wire N__69492;
    wire N__69491;
    wire N__69488;
    wire N__69487;
    wire N__69486;
    wire N__69483;
    wire N__69482;
    wire N__69481;
    wire N__69480;
    wire N__69477;
    wire N__69474;
    wire N__69471;
    wire N__69468;
    wire N__69465;
    wire N__69456;
    wire N__69453;
    wire N__69452;
    wire N__69451;
    wire N__69450;
    wire N__69447;
    wire N__69442;
    wire N__69439;
    wire N__69436;
    wire N__69433;
    wire N__69430;
    wire N__69427;
    wire N__69424;
    wire N__69421;
    wire N__69418;
    wire N__69413;
    wire N__69410;
    wire N__69405;
    wire N__69400;
    wire N__69397;
    wire N__69394;
    wire N__69391;
    wire N__69388;
    wire N__69385;
    wire N__69376;
    wire N__69375;
    wire N__69374;
    wire N__69371;
    wire N__69368;
    wire N__69365;
    wire N__69360;
    wire N__69355;
    wire N__69352;
    wire N__69349;
    wire N__69344;
    wire N__69341;
    wire N__69338;
    wire N__69335;
    wire N__69330;
    wire N__69327;
    wire N__69324;
    wire N__69319;
    wire N__69314;
    wire N__69309;
    wire N__69304;
    wire N__69295;
    wire N__69280;
    wire N__69279;
    wire N__69276;
    wire N__69273;
    wire N__69270;
    wire N__69269;
    wire N__69266;
    wire N__69263;
    wire N__69260;
    wire N__69253;
    wire N__69250;
    wire N__69249;
    wire N__69246;
    wire N__69245;
    wire N__69244;
    wire N__69241;
    wire N__69238;
    wire N__69235;
    wire N__69234;
    wire N__69233;
    wire N__69232;
    wire N__69231;
    wire N__69228;
    wire N__69227;
    wire N__69226;
    wire N__69223;
    wire N__69220;
    wire N__69217;
    wire N__69214;
    wire N__69213;
    wire N__69212;
    wire N__69211;
    wire N__69210;
    wire N__69207;
    wire N__69206;
    wire N__69205;
    wire N__69204;
    wire N__69203;
    wire N__69200;
    wire N__69199;
    wire N__69198;
    wire N__69197;
    wire N__69194;
    wire N__69193;
    wire N__69192;
    wire N__69191;
    wire N__69184;
    wire N__69177;
    wire N__69174;
    wire N__69169;
    wire N__69168;
    wire N__69165;
    wire N__69162;
    wire N__69155;
    wire N__69152;
    wire N__69151;
    wire N__69148;
    wire N__69143;
    wire N__69138;
    wire N__69135;
    wire N__69132;
    wire N__69129;
    wire N__69126;
    wire N__69125;
    wire N__69124;
    wire N__69119;
    wire N__69116;
    wire N__69113;
    wire N__69110;
    wire N__69107;
    wire N__69100;
    wire N__69097;
    wire N__69094;
    wire N__69089;
    wire N__69086;
    wire N__69081;
    wire N__69078;
    wire N__69075;
    wire N__69072;
    wire N__69069;
    wire N__69066;
    wire N__69065;
    wire N__69064;
    wire N__69063;
    wire N__69062;
    wire N__69059;
    wire N__69056;
    wire N__69053;
    wire N__69050;
    wire N__69043;
    wire N__69034;
    wire N__69027;
    wire N__69018;
    wire N__69015;
    wire N__69008;
    wire N__69005;
    wire N__69000;
    wire N__68989;
    wire N__68988;
    wire N__68987;
    wire N__68984;
    wire N__68981;
    wire N__68980;
    wire N__68979;
    wire N__68976;
    wire N__68975;
    wire N__68974;
    wire N__68973;
    wire N__68972;
    wire N__68971;
    wire N__68970;
    wire N__68965;
    wire N__68962;
    wire N__68959;
    wire N__68958;
    wire N__68957;
    wire N__68956;
    wire N__68955;
    wire N__68954;
    wire N__68951;
    wire N__68948;
    wire N__68945;
    wire N__68944;
    wire N__68941;
    wire N__68940;
    wire N__68939;
    wire N__68938;
    wire N__68935;
    wire N__68932;
    wire N__68929;
    wire N__68926;
    wire N__68921;
    wire N__68916;
    wire N__68913;
    wire N__68910;
    wire N__68909;
    wire N__68908;
    wire N__68905;
    wire N__68900;
    wire N__68897;
    wire N__68894;
    wire N__68889;
    wire N__68884;
    wire N__68883;
    wire N__68882;
    wire N__68881;
    wire N__68880;
    wire N__68877;
    wire N__68876;
    wire N__68873;
    wire N__68868;
    wire N__68867;
    wire N__68866;
    wire N__68865;
    wire N__68862;
    wire N__68855;
    wire N__68852;
    wire N__68849;
    wire N__68846;
    wire N__68837;
    wire N__68834;
    wire N__68831;
    wire N__68826;
    wire N__68823;
    wire N__68820;
    wire N__68817;
    wire N__68812;
    wire N__68809;
    wire N__68806;
    wire N__68803;
    wire N__68800;
    wire N__68797;
    wire N__68792;
    wire N__68789;
    wire N__68786;
    wire N__68785;
    wire N__68784;
    wire N__68781;
    wire N__68776;
    wire N__68771;
    wire N__68766;
    wire N__68763;
    wire N__68756;
    wire N__68753;
    wire N__68746;
    wire N__68743;
    wire N__68740;
    wire N__68731;
    wire N__68722;
    wire N__68713;
    wire N__68712;
    wire N__68709;
    wire N__68706;
    wire N__68705;
    wire N__68702;
    wire N__68699;
    wire N__68696;
    wire N__68695;
    wire N__68690;
    wire N__68685;
    wire N__68680;
    wire N__68679;
    wire N__68678;
    wire N__68675;
    wire N__68674;
    wire N__68673;
    wire N__68672;
    wire N__68671;
    wire N__68670;
    wire N__68669;
    wire N__68666;
    wire N__68663;
    wire N__68660;
    wire N__68659;
    wire N__68658;
    wire N__68655;
    wire N__68650;
    wire N__68647;
    wire N__68644;
    wire N__68639;
    wire N__68638;
    wire N__68633;
    wire N__68632;
    wire N__68629;
    wire N__68628;
    wire N__68625;
    wire N__68620;
    wire N__68617;
    wire N__68614;
    wire N__68611;
    wire N__68608;
    wire N__68605;
    wire N__68602;
    wire N__68601;
    wire N__68600;
    wire N__68595;
    wire N__68592;
    wire N__68591;
    wire N__68590;
    wire N__68589;
    wire N__68584;
    wire N__68579;
    wire N__68576;
    wire N__68571;
    wire N__68570;
    wire N__68569;
    wire N__68568;
    wire N__68565;
    wire N__68562;
    wire N__68557;
    wire N__68554;
    wire N__68553;
    wire N__68552;
    wire N__68549;
    wire N__68546;
    wire N__68545;
    wire N__68542;
    wire N__68539;
    wire N__68536;
    wire N__68533;
    wire N__68530;
    wire N__68527;
    wire N__68524;
    wire N__68517;
    wire N__68516;
    wire N__68513;
    wire N__68506;
    wire N__68503;
    wire N__68500;
    wire N__68493;
    wire N__68488;
    wire N__68485;
    wire N__68480;
    wire N__68477;
    wire N__68468;
    wire N__68463;
    wire N__68460;
    wire N__68457;
    wire N__68450;
    wire N__68443;
    wire N__68442;
    wire N__68441;
    wire N__68438;
    wire N__68437;
    wire N__68436;
    wire N__68435;
    wire N__68434;
    wire N__68433;
    wire N__68430;
    wire N__68427;
    wire N__68426;
    wire N__68423;
    wire N__68420;
    wire N__68419;
    wire N__68418;
    wire N__68417;
    wire N__68416;
    wire N__68413;
    wire N__68412;
    wire N__68411;
    wire N__68410;
    wire N__68407;
    wire N__68404;
    wire N__68399;
    wire N__68396;
    wire N__68395;
    wire N__68394;
    wire N__68393;
    wire N__68390;
    wire N__68385;
    wire N__68378;
    wire N__68377;
    wire N__68374;
    wire N__68373;
    wire N__68370;
    wire N__68369;
    wire N__68366;
    wire N__68363;
    wire N__68360;
    wire N__68359;
    wire N__68358;
    wire N__68357;
    wire N__68356;
    wire N__68355;
    wire N__68354;
    wire N__68353;
    wire N__68352;
    wire N__68349;
    wire N__68346;
    wire N__68341;
    wire N__68338;
    wire N__68333;
    wire N__68330;
    wire N__68325;
    wire N__68322;
    wire N__68319;
    wire N__68316;
    wire N__68313;
    wire N__68310;
    wire N__68307;
    wire N__68304;
    wire N__68301;
    wire N__68296;
    wire N__68293;
    wire N__68290;
    wire N__68289;
    wire N__68288;
    wire N__68285;
    wire N__68280;
    wire N__68277;
    wire N__68274;
    wire N__68269;
    wire N__68262;
    wire N__68259;
    wire N__68256;
    wire N__68251;
    wire N__68248;
    wire N__68243;
    wire N__68238;
    wire N__68235;
    wire N__68230;
    wire N__68227;
    wire N__68224;
    wire N__68219;
    wire N__68216;
    wire N__68211;
    wire N__68208;
    wire N__68205;
    wire N__68196;
    wire N__68189;
    wire N__68178;
    wire N__68167;
    wire N__68166;
    wire N__68165;
    wire N__68164;
    wire N__68163;
    wire N__68162;
    wire N__68161;
    wire N__68160;
    wire N__68159;
    wire N__68158;
    wire N__68157;
    wire N__68156;
    wire N__68155;
    wire N__68152;
    wire N__68149;
    wire N__68148;
    wire N__68147;
    wire N__68146;
    wire N__68145;
    wire N__68144;
    wire N__68143;
    wire N__68142;
    wire N__68141;
    wire N__68140;
    wire N__68139;
    wire N__68138;
    wire N__68137;
    wire N__68136;
    wire N__68135;
    wire N__68132;
    wire N__68129;
    wire N__68122;
    wire N__68117;
    wire N__68112;
    wire N__68111;
    wire N__68110;
    wire N__68109;
    wire N__68104;
    wire N__68101;
    wire N__68098;
    wire N__68097;
    wire N__68096;
    wire N__68095;
    wire N__68094;
    wire N__68093;
    wire N__68092;
    wire N__68091;
    wire N__68088;
    wire N__68087;
    wire N__68086;
    wire N__68083;
    wire N__68078;
    wire N__68071;
    wire N__68070;
    wire N__68069;
    wire N__68068;
    wire N__68067;
    wire N__68066;
    wire N__68065;
    wire N__68062;
    wire N__68057;
    wire N__68048;
    wire N__68045;
    wire N__68044;
    wire N__68043;
    wire N__68042;
    wire N__68039;
    wire N__68036;
    wire N__68033;
    wire N__68030;
    wire N__68023;
    wire N__68020;
    wire N__68019;
    wire N__68018;
    wire N__68017;
    wire N__68012;
    wire N__68009;
    wire N__68008;
    wire N__68007;
    wire N__68006;
    wire N__68003;
    wire N__68000;
    wire N__67995;
    wire N__67990;
    wire N__67987;
    wire N__67984;
    wire N__67979;
    wire N__67974;
    wire N__67971;
    wire N__67966;
    wire N__67959;
    wire N__67954;
    wire N__67949;
    wire N__67946;
    wire N__67941;
    wire N__67938;
    wire N__67933;
    wire N__67926;
    wire N__67919;
    wire N__67916;
    wire N__67913;
    wire N__67912;
    wire N__67911;
    wire N__67904;
    wire N__67901;
    wire N__67892;
    wire N__67885;
    wire N__67874;
    wire N__67871;
    wire N__67866;
    wire N__67861;
    wire N__67854;
    wire N__67849;
    wire N__67838;
    wire N__67831;
    wire N__67828;
    wire N__67819;
    wire N__67818;
    wire N__67815;
    wire N__67812;
    wire N__67811;
    wire N__67808;
    wire N__67805;
    wire N__67802;
    wire N__67795;
    wire N__67794;
    wire N__67793;
    wire N__67792;
    wire N__67791;
    wire N__67784;
    wire N__67779;
    wire N__67778;
    wire N__67777;
    wire N__67776;
    wire N__67775;
    wire N__67770;
    wire N__67765;
    wire N__67764;
    wire N__67763;
    wire N__67762;
    wire N__67761;
    wire N__67760;
    wire N__67759;
    wire N__67758;
    wire N__67757;
    wire N__67756;
    wire N__67753;
    wire N__67752;
    wire N__67751;
    wire N__67750;
    wire N__67749;
    wire N__67748;
    wire N__67745;
    wire N__67744;
    wire N__67739;
    wire N__67734;
    wire N__67733;
    wire N__67732;
    wire N__67731;
    wire N__67724;
    wire N__67721;
    wire N__67718;
    wire N__67715;
    wire N__67712;
    wire N__67709;
    wire N__67708;
    wire N__67707;
    wire N__67706;
    wire N__67705;
    wire N__67702;
    wire N__67699;
    wire N__67692;
    wire N__67689;
    wire N__67686;
    wire N__67685;
    wire N__67682;
    wire N__67679;
    wire N__67678;
    wire N__67677;
    wire N__67676;
    wire N__67675;
    wire N__67674;
    wire N__67673;
    wire N__67672;
    wire N__67665;
    wire N__67662;
    wire N__67659;
    wire N__67656;
    wire N__67649;
    wire N__67646;
    wire N__67643;
    wire N__67638;
    wire N__67633;
    wire N__67630;
    wire N__67625;
    wire N__67624;
    wire N__67623;
    wire N__67622;
    wire N__67621;
    wire N__67620;
    wire N__67617;
    wire N__67612;
    wire N__67611;
    wire N__67610;
    wire N__67609;
    wire N__67606;
    wire N__67603;
    wire N__67600;
    wire N__67597;
    wire N__67592;
    wire N__67589;
    wire N__67586;
    wire N__67583;
    wire N__67576;
    wire N__67573;
    wire N__67564;
    wire N__67561;
    wire N__67556;
    wire N__67553;
    wire N__67548;
    wire N__67545;
    wire N__67542;
    wire N__67539;
    wire N__67536;
    wire N__67533;
    wire N__67522;
    wire N__67513;
    wire N__67506;
    wire N__67495;
    wire N__67480;
    wire N__67479;
    wire N__67478;
    wire N__67477;
    wire N__67476;
    wire N__67475;
    wire N__67472;
    wire N__67471;
    wire N__67470;
    wire N__67469;
    wire N__67466;
    wire N__67463;
    wire N__67462;
    wire N__67461;
    wire N__67460;
    wire N__67459;
    wire N__67458;
    wire N__67457;
    wire N__67454;
    wire N__67453;
    wire N__67452;
    wire N__67451;
    wire N__67446;
    wire N__67445;
    wire N__67440;
    wire N__67437;
    wire N__67434;
    wire N__67425;
    wire N__67418;
    wire N__67415;
    wire N__67412;
    wire N__67409;
    wire N__67408;
    wire N__67407;
    wire N__67404;
    wire N__67403;
    wire N__67402;
    wire N__67399;
    wire N__67396;
    wire N__67393;
    wire N__67392;
    wire N__67391;
    wire N__67386;
    wire N__67383;
    wire N__67380;
    wire N__67379;
    wire N__67376;
    wire N__67373;
    wire N__67368;
    wire N__67365;
    wire N__67364;
    wire N__67363;
    wire N__67362;
    wire N__67361;
    wire N__67358;
    wire N__67355;
    wire N__67352;
    wire N__67349;
    wire N__67348;
    wire N__67345;
    wire N__67340;
    wire N__67339;
    wire N__67334;
    wire N__67331;
    wire N__67326;
    wire N__67323;
    wire N__67320;
    wire N__67317;
    wire N__67312;
    wire N__67307;
    wire N__67304;
    wire N__67301;
    wire N__67296;
    wire N__67293;
    wire N__67290;
    wire N__67287;
    wire N__67282;
    wire N__67279;
    wire N__67272;
    wire N__67269;
    wire N__67262;
    wire N__67251;
    wire N__67240;
    wire N__67237;
    wire N__67234;
    wire N__67231;
    wire N__67228;
    wire N__67219;
    wire N__67218;
    wire N__67217;
    wire N__67216;
    wire N__67215;
    wire N__67214;
    wire N__67211;
    wire N__67210;
    wire N__67209;
    wire N__67208;
    wire N__67207;
    wire N__67206;
    wire N__67203;
    wire N__67202;
    wire N__67201;
    wire N__67196;
    wire N__67193;
    wire N__67190;
    wire N__67187;
    wire N__67186;
    wire N__67183;
    wire N__67180;
    wire N__67177;
    wire N__67172;
    wire N__67171;
    wire N__67170;
    wire N__67167;
    wire N__67164;
    wire N__67163;
    wire N__67162;
    wire N__67161;
    wire N__67158;
    wire N__67157;
    wire N__67154;
    wire N__67149;
    wire N__67146;
    wire N__67143;
    wire N__67142;
    wire N__67139;
    wire N__67134;
    wire N__67131;
    wire N__67128;
    wire N__67125;
    wire N__67124;
    wire N__67123;
    wire N__67122;
    wire N__67117;
    wire N__67114;
    wire N__67111;
    wire N__67108;
    wire N__67105;
    wire N__67104;
    wire N__67103;
    wire N__67100;
    wire N__67097;
    wire N__67094;
    wire N__67089;
    wire N__67086;
    wire N__67083;
    wire N__67080;
    wire N__67079;
    wire N__67076;
    wire N__67071;
    wire N__67070;
    wire N__67067;
    wire N__67064;
    wire N__67063;
    wire N__67060;
    wire N__67057;
    wire N__67054;
    wire N__67051;
    wire N__67046;
    wire N__67043;
    wire N__67040;
    wire N__67033;
    wire N__67030;
    wire N__67027;
    wire N__67022;
    wire N__67019;
    wire N__67014;
    wire N__67011;
    wire N__67006;
    wire N__67005;
    wire N__67002;
    wire N__66991;
    wire N__66982;
    wire N__66979;
    wire N__66976;
    wire N__66975;
    wire N__66974;
    wire N__66971;
    wire N__66968;
    wire N__66963;
    wire N__66960;
    wire N__66953;
    wire N__66948;
    wire N__66945;
    wire N__66942;
    wire N__66939;
    wire N__66934;
    wire N__66929;
    wire N__66926;
    wire N__66913;
    wire N__66912;
    wire N__66909;
    wire N__66908;
    wire N__66905;
    wire N__66902;
    wire N__66899;
    wire N__66896;
    wire N__66893;
    wire N__66890;
    wire N__66883;
    wire N__66880;
    wire N__66877;
    wire N__66876;
    wire N__66875;
    wire N__66872;
    wire N__66871;
    wire N__66870;
    wire N__66869;
    wire N__66868;
    wire N__66867;
    wire N__66866;
    wire N__66865;
    wire N__66864;
    wire N__66863;
    wire N__66862;
    wire N__66861;
    wire N__66860;
    wire N__66859;
    wire N__66858;
    wire N__66857;
    wire N__66856;
    wire N__66855;
    wire N__66854;
    wire N__66853;
    wire N__66852;
    wire N__66851;
    wire N__66850;
    wire N__66849;
    wire N__66848;
    wire N__66847;
    wire N__66846;
    wire N__66845;
    wire N__66844;
    wire N__66843;
    wire N__66842;
    wire N__66841;
    wire N__66840;
    wire N__66839;
    wire N__66838;
    wire N__66837;
    wire N__66836;
    wire N__66835;
    wire N__66834;
    wire N__66833;
    wire N__66832;
    wire N__66831;
    wire N__66830;
    wire N__66829;
    wire N__66828;
    wire N__66827;
    wire N__66826;
    wire N__66825;
    wire N__66824;
    wire N__66823;
    wire N__66822;
    wire N__66821;
    wire N__66820;
    wire N__66819;
    wire N__66818;
    wire N__66817;
    wire N__66816;
    wire N__66815;
    wire N__66814;
    wire N__66813;
    wire N__66812;
    wire N__66811;
    wire N__66810;
    wire N__66809;
    wire N__66808;
    wire N__66807;
    wire N__66806;
    wire N__66805;
    wire N__66804;
    wire N__66803;
    wire N__66802;
    wire N__66801;
    wire N__66800;
    wire N__66799;
    wire N__66798;
    wire N__66797;
    wire N__66796;
    wire N__66795;
    wire N__66794;
    wire N__66793;
    wire N__66792;
    wire N__66791;
    wire N__66790;
    wire N__66789;
    wire N__66788;
    wire N__66787;
    wire N__66786;
    wire N__66785;
    wire N__66784;
    wire N__66783;
    wire N__66782;
    wire N__66781;
    wire N__66780;
    wire N__66779;
    wire N__66778;
    wire N__66777;
    wire N__66776;
    wire N__66775;
    wire N__66774;
    wire N__66773;
    wire N__66772;
    wire N__66771;
    wire N__66770;
    wire N__66769;
    wire N__66768;
    wire N__66767;
    wire N__66766;
    wire N__66765;
    wire N__66764;
    wire N__66763;
    wire N__66762;
    wire N__66761;
    wire N__66760;
    wire N__66759;
    wire N__66758;
    wire N__66757;
    wire N__66756;
    wire N__66755;
    wire N__66754;
    wire N__66753;
    wire N__66752;
    wire N__66751;
    wire N__66750;
    wire N__66749;
    wire N__66748;
    wire N__66747;
    wire N__66746;
    wire N__66745;
    wire N__66744;
    wire N__66743;
    wire N__66742;
    wire N__66741;
    wire N__66740;
    wire N__66739;
    wire N__66738;
    wire N__66737;
    wire N__66736;
    wire N__66735;
    wire N__66734;
    wire N__66733;
    wire N__66732;
    wire N__66731;
    wire N__66730;
    wire N__66729;
    wire N__66728;
    wire N__66727;
    wire N__66726;
    wire N__66725;
    wire N__66724;
    wire N__66723;
    wire N__66722;
    wire N__66721;
    wire N__66720;
    wire N__66719;
    wire N__66718;
    wire N__66717;
    wire N__66716;
    wire N__66715;
    wire N__66714;
    wire N__66713;
    wire N__66712;
    wire N__66711;
    wire N__66710;
    wire N__66709;
    wire N__66708;
    wire N__66707;
    wire N__66706;
    wire N__66705;
    wire N__66704;
    wire N__66703;
    wire N__66702;
    wire N__66701;
    wire N__66700;
    wire N__66699;
    wire N__66698;
    wire N__66697;
    wire N__66696;
    wire N__66695;
    wire N__66694;
    wire N__66693;
    wire N__66692;
    wire N__66691;
    wire N__66690;
    wire N__66689;
    wire N__66688;
    wire N__66687;
    wire N__66686;
    wire N__66685;
    wire N__66684;
    wire N__66683;
    wire N__66682;
    wire N__66681;
    wire N__66680;
    wire N__66679;
    wire N__66678;
    wire N__66677;
    wire N__66676;
    wire N__66675;
    wire N__66674;
    wire N__66673;
    wire N__66672;
    wire N__66671;
    wire N__66670;
    wire N__66669;
    wire N__66668;
    wire N__66667;
    wire N__66666;
    wire N__66665;
    wire N__66664;
    wire N__66663;
    wire N__66662;
    wire N__66661;
    wire N__66660;
    wire N__66659;
    wire N__66658;
    wire N__66657;
    wire N__66656;
    wire N__66655;
    wire N__66654;
    wire N__66653;
    wire N__66652;
    wire N__66651;
    wire N__66650;
    wire N__66649;
    wire N__66648;
    wire N__66647;
    wire N__66646;
    wire N__66645;
    wire N__66644;
    wire N__66643;
    wire N__66642;
    wire N__66641;
    wire N__66640;
    wire N__66639;
    wire N__66638;
    wire N__66637;
    wire N__66636;
    wire N__66635;
    wire N__66634;
    wire N__66633;
    wire N__66632;
    wire N__66631;
    wire N__66630;
    wire N__66139;
    wire N__66136;
    wire N__66135;
    wire N__66132;
    wire N__66129;
    wire N__66128;
    wire N__66125;
    wire N__66124;
    wire N__66121;
    wire N__66118;
    wire N__66115;
    wire N__66112;
    wire N__66107;
    wire N__66104;
    wire N__66097;
    wire N__66096;
    wire N__66095;
    wire N__66092;
    wire N__66089;
    wire N__66086;
    wire N__66083;
    wire N__66080;
    wire N__66077;
    wire N__66072;
    wire N__66067;
    wire N__66066;
    wire N__66065;
    wire N__66060;
    wire N__66057;
    wire N__66054;
    wire N__66049;
    wire N__66048;
    wire N__66045;
    wire N__66042;
    wire N__66039;
    wire N__66034;
    wire N__66031;
    wire N__66030;
    wire N__66029;
    wire N__66028;
    wire N__66025;
    wire N__66022;
    wire N__66021;
    wire N__66020;
    wire N__66019;
    wire N__66016;
    wire N__66015;
    wire N__66014;
    wire N__66013;
    wire N__66012;
    wire N__66009;
    wire N__66008;
    wire N__66007;
    wire N__66004;
    wire N__66003;
    wire N__66002;
    wire N__66001;
    wire N__65998;
    wire N__65993;
    wire N__65992;
    wire N__65991;
    wire N__65988;
    wire N__65985;
    wire N__65982;
    wire N__65977;
    wire N__65974;
    wire N__65973;
    wire N__65972;
    wire N__65971;
    wire N__65970;
    wire N__65969;
    wire N__65964;
    wire N__65961;
    wire N__65958;
    wire N__65953;
    wire N__65950;
    wire N__65949;
    wire N__65944;
    wire N__65941;
    wire N__65940;
    wire N__65939;
    wire N__65938;
    wire N__65937;
    wire N__65936;
    wire N__65933;
    wire N__65932;
    wire N__65929;
    wire N__65926;
    wire N__65923;
    wire N__65920;
    wire N__65917;
    wire N__65908;
    wire N__65905;
    wire N__65900;
    wire N__65899;
    wire N__65894;
    wire N__65891;
    wire N__65888;
    wire N__65885;
    wire N__65882;
    wire N__65879;
    wire N__65876;
    wire N__65869;
    wire N__65866;
    wire N__65865;
    wire N__65862;
    wire N__65859;
    wire N__65850;
    wire N__65847;
    wire N__65842;
    wire N__65839;
    wire N__65834;
    wire N__65825;
    wire N__65822;
    wire N__65819;
    wire N__65816;
    wire N__65813;
    wire N__65806;
    wire N__65801;
    wire N__65798;
    wire N__65793;
    wire N__65788;
    wire N__65785;
    wire N__65780;
    wire N__65777;
    wire N__65772;
    wire N__65761;
    wire N__65760;
    wire N__65759;
    wire N__65756;
    wire N__65751;
    wire N__65750;
    wire N__65747;
    wire N__65744;
    wire N__65741;
    wire N__65738;
    wire N__65735;
    wire N__65732;
    wire N__65729;
    wire N__65726;
    wire N__65719;
    wire N__65718;
    wire N__65715;
    wire N__65712;
    wire N__65709;
    wire N__65706;
    wire N__65703;
    wire N__65698;
    wire N__65697;
    wire N__65696;
    wire N__65693;
    wire N__65690;
    wire N__65689;
    wire N__65686;
    wire N__65681;
    wire N__65678;
    wire N__65675;
    wire N__65674;
    wire N__65673;
    wire N__65672;
    wire N__65671;
    wire N__65670;
    wire N__65667;
    wire N__65662;
    wire N__65661;
    wire N__65658;
    wire N__65655;
    wire N__65650;
    wire N__65649;
    wire N__65648;
    wire N__65647;
    wire N__65644;
    wire N__65639;
    wire N__65636;
    wire N__65631;
    wire N__65628;
    wire N__65625;
    wire N__65624;
    wire N__65623;
    wire N__65620;
    wire N__65617;
    wire N__65604;
    wire N__65601;
    wire N__65598;
    wire N__65595;
    wire N__65592;
    wire N__65591;
    wire N__65588;
    wire N__65583;
    wire N__65582;
    wire N__65577;
    wire N__65576;
    wire N__65575;
    wire N__65574;
    wire N__65573;
    wire N__65572;
    wire N__65571;
    wire N__65570;
    wire N__65569;
    wire N__65568;
    wire N__65567;
    wire N__65564;
    wire N__65563;
    wire N__65562;
    wire N__65557;
    wire N__65554;
    wire N__65551;
    wire N__65548;
    wire N__65545;
    wire N__65542;
    wire N__65537;
    wire N__65532;
    wire N__65529;
    wire N__65524;
    wire N__65521;
    wire N__65518;
    wire N__65515;
    wire N__65512;
    wire N__65509;
    wire N__65504;
    wire N__65503;
    wire N__65502;
    wire N__65501;
    wire N__65498;
    wire N__65495;
    wire N__65492;
    wire N__65489;
    wire N__65486;
    wire N__65481;
    wire N__65470;
    wire N__65465;
    wire N__65462;
    wire N__65459;
    wire N__65454;
    wire N__65451;
    wire N__65446;
    wire N__65443;
    wire N__65428;
    wire N__65425;
    wire N__65424;
    wire N__65421;
    wire N__65418;
    wire N__65417;
    wire N__65414;
    wire N__65409;
    wire N__65404;
    wire N__65401;
    wire N__65400;
    wire N__65397;
    wire N__65394;
    wire N__65391;
    wire N__65388;
    wire N__65385;
    wire N__65380;
    wire N__65379;
    wire N__65378;
    wire N__65375;
    wire N__65370;
    wire N__65365;
    wire N__65364;
    wire N__65361;
    wire N__65358;
    wire N__65357;
    wire N__65356;
    wire N__65355;
    wire N__65352;
    wire N__65349;
    wire N__65344;
    wire N__65341;
    wire N__65338;
    wire N__65335;
    wire N__65326;
    wire N__65323;
    wire N__65322;
    wire N__65319;
    wire N__65316;
    wire N__65311;
    wire N__65308;
    wire N__65305;
    wire N__65304;
    wire N__65301;
    wire N__65298;
    wire N__65297;
    wire N__65292;
    wire N__65289;
    wire N__65286;
    wire N__65283;
    wire N__65280;
    wire N__65275;
    wire N__65272;
    wire N__65269;
    wire N__65266;
    wire N__65265;
    wire N__65262;
    wire N__65259;
    wire N__65256;
    wire N__65253;
    wire N__65248;
    wire N__65247;
    wire N__65246;
    wire N__65245;
    wire N__65242;
    wire N__65239;
    wire N__65234;
    wire N__65231;
    wire N__65230;
    wire N__65227;
    wire N__65224;
    wire N__65221;
    wire N__65218;
    wire N__65213;
    wire N__65206;
    wire N__65203;
    wire N__65200;
    wire N__65197;
    wire N__65194;
    wire N__65193;
    wire N__65192;
    wire N__65189;
    wire N__65186;
    wire N__65183;
    wire N__65180;
    wire N__65179;
    wire N__65176;
    wire N__65173;
    wire N__65170;
    wire N__65167;
    wire N__65164;
    wire N__65155;
    wire N__65154;
    wire N__65153;
    wire N__65150;
    wire N__65147;
    wire N__65146;
    wire N__65143;
    wire N__65140;
    wire N__65137;
    wire N__65134;
    wire N__65131;
    wire N__65128;
    wire N__65123;
    wire N__65120;
    wire N__65113;
    wire N__65110;
    wire N__65107;
    wire N__65104;
    wire N__65103;
    wire N__65100;
    wire N__65097;
    wire N__65094;
    wire N__65091;
    wire N__65086;
    wire N__65083;
    wire N__65080;
    wire N__65077;
    wire N__65074;
    wire N__65073;
    wire N__65070;
    wire N__65067;
    wire N__65062;
    wire N__65061;
    wire N__65060;
    wire N__65059;
    wire N__65054;
    wire N__65053;
    wire N__65050;
    wire N__65047;
    wire N__65044;
    wire N__65041;
    wire N__65038;
    wire N__65035;
    wire N__65032;
    wire N__65029;
    wire N__65020;
    wire N__65017;
    wire N__65016;
    wire N__65013;
    wire N__65010;
    wire N__65007;
    wire N__65004;
    wire N__65001;
    wire N__64998;
    wire N__64995;
    wire N__64990;
    wire N__64989;
    wire N__64986;
    wire N__64983;
    wire N__64980;
    wire N__64975;
    wire N__64972;
    wire N__64969;
    wire N__64966;
    wire N__64963;
    wire N__64962;
    wire N__64957;
    wire N__64954;
    wire N__64951;
    wire N__64948;
    wire N__64947;
    wire N__64944;
    wire N__64941;
    wire N__64938;
    wire N__64933;
    wire N__64932;
    wire N__64929;
    wire N__64926;
    wire N__64923;
    wire N__64920;
    wire N__64917;
    wire N__64912;
    wire N__64911;
    wire N__64908;
    wire N__64905;
    wire N__64900;
    wire N__64897;
    wire N__64894;
    wire N__64893;
    wire N__64892;
    wire N__64889;
    wire N__64888;
    wire N__64887;
    wire N__64886;
    wire N__64885;
    wire N__64884;
    wire N__64883;
    wire N__64880;
    wire N__64879;
    wire N__64876;
    wire N__64875;
    wire N__64874;
    wire N__64873;
    wire N__64872;
    wire N__64871;
    wire N__64868;
    wire N__64865;
    wire N__64864;
    wire N__64863;
    wire N__64862;
    wire N__64859;
    wire N__64854;
    wire N__64853;
    wire N__64852;
    wire N__64851;
    wire N__64846;
    wire N__64843;
    wire N__64840;
    wire N__64837;
    wire N__64836;
    wire N__64833;
    wire N__64830;
    wire N__64827;
    wire N__64826;
    wire N__64825;
    wire N__64824;
    wire N__64823;
    wire N__64820;
    wire N__64819;
    wire N__64818;
    wire N__64815;
    wire N__64812;
    wire N__64809;
    wire N__64806;
    wire N__64803;
    wire N__64800;
    wire N__64797;
    wire N__64794;
    wire N__64789;
    wire N__64786;
    wire N__64781;
    wire N__64778;
    wire N__64775;
    wire N__64772;
    wire N__64767;
    wire N__64764;
    wire N__64761;
    wire N__64758;
    wire N__64755;
    wire N__64752;
    wire N__64749;
    wire N__64748;
    wire N__64745;
    wire N__64742;
    wire N__64739;
    wire N__64734;
    wire N__64731;
    wire N__64726;
    wire N__64721;
    wire N__64718;
    wire N__64715;
    wire N__64706;
    wire N__64701;
    wire N__64700;
    wire N__64699;
    wire N__64698;
    wire N__64695;
    wire N__64692;
    wire N__64689;
    wire N__64686;
    wire N__64683;
    wire N__64678;
    wire N__64671;
    wire N__64668;
    wire N__64665;
    wire N__64660;
    wire N__64653;
    wire N__64650;
    wire N__64645;
    wire N__64642;
    wire N__64633;
    wire N__64626;
    wire N__64621;
    wire N__64618;
    wire N__64603;
    wire N__64600;
    wire N__64599;
    wire N__64596;
    wire N__64593;
    wire N__64588;
    wire N__64587;
    wire N__64584;
    wire N__64581;
    wire N__64578;
    wire N__64575;
    wire N__64572;
    wire N__64567;
    wire N__64566;
    wire N__64565;
    wire N__64562;
    wire N__64561;
    wire N__64560;
    wire N__64557;
    wire N__64556;
    wire N__64553;
    wire N__64552;
    wire N__64551;
    wire N__64550;
    wire N__64549;
    wire N__64546;
    wire N__64543;
    wire N__64540;
    wire N__64537;
    wire N__64536;
    wire N__64535;
    wire N__64534;
    wire N__64533;
    wire N__64532;
    wire N__64531;
    wire N__64528;
    wire N__64527;
    wire N__64524;
    wire N__64523;
    wire N__64520;
    wire N__64519;
    wire N__64518;
    wire N__64517;
    wire N__64514;
    wire N__64513;
    wire N__64512;
    wire N__64511;
    wire N__64508;
    wire N__64505;
    wire N__64502;
    wire N__64499;
    wire N__64498;
    wire N__64495;
    wire N__64492;
    wire N__64487;
    wire N__64482;
    wire N__64481;
    wire N__64478;
    wire N__64473;
    wire N__64470;
    wire N__64467;
    wire N__64464;
    wire N__64459;
    wire N__64458;
    wire N__64455;
    wire N__64452;
    wire N__64451;
    wire N__64448;
    wire N__64441;
    wire N__64438;
    wire N__64435;
    wire N__64430;
    wire N__64427;
    wire N__64420;
    wire N__64417;
    wire N__64414;
    wire N__64411;
    wire N__64404;
    wire N__64399;
    wire N__64396;
    wire N__64391;
    wire N__64388;
    wire N__64385;
    wire N__64382;
    wire N__64375;
    wire N__64372;
    wire N__64365;
    wire N__64358;
    wire N__64357;
    wire N__64356;
    wire N__64353;
    wire N__64350;
    wire N__64347;
    wire N__64346;
    wire N__64345;
    wire N__64342;
    wire N__64339;
    wire N__64336;
    wire N__64333;
    wire N__64328;
    wire N__64323;
    wire N__64316;
    wire N__64313;
    wire N__64310;
    wire N__64305;
    wire N__64302;
    wire N__64299;
    wire N__64296;
    wire N__64291;
    wire N__64276;
    wire N__64275;
    wire N__64272;
    wire N__64269;
    wire N__64266;
    wire N__64263;
    wire N__64258;
    wire N__64257;
    wire N__64254;
    wire N__64251;
    wire N__64248;
    wire N__64245;
    wire N__64244;
    wire N__64239;
    wire N__64236;
    wire N__64231;
    wire N__64228;
    wire N__64225;
    wire N__64224;
    wire N__64221;
    wire N__64220;
    wire N__64219;
    wire N__64216;
    wire N__64213;
    wire N__64208;
    wire N__64207;
    wire N__64204;
    wire N__64199;
    wire N__64196;
    wire N__64189;
    wire N__64186;
    wire N__64183;
    wire N__64180;
    wire N__64177;
    wire N__64174;
    wire N__64173;
    wire N__64170;
    wire N__64167;
    wire N__64164;
    wire N__64161;
    wire N__64156;
    wire N__64153;
    wire N__64152;
    wire N__64149;
    wire N__64146;
    wire N__64141;
    wire N__64138;
    wire N__64135;
    wire N__64132;
    wire N__64129;
    wire N__64126;
    wire N__64123;
    wire N__64122;
    wire N__64119;
    wire N__64116;
    wire N__64111;
    wire N__64110;
    wire N__64109;
    wire N__64106;
    wire N__64101;
    wire N__64098;
    wire N__64095;
    wire N__64092;
    wire N__64089;
    wire N__64084;
    wire N__64081;
    wire N__64078;
    wire N__64075;
    wire N__64072;
    wire N__64069;
    wire N__64066;
    wire N__64065;
    wire N__64062;
    wire N__64059;
    wire N__64054;
    wire N__64051;
    wire N__64048;
    wire N__64045;
    wire N__64042;
    wire N__64039;
    wire N__64036;
    wire N__64035;
    wire N__64034;
    wire N__64031;
    wire N__64030;
    wire N__64027;
    wire N__64024;
    wire N__64021;
    wire N__64018;
    wire N__64017;
    wire N__64014;
    wire N__64011;
    wire N__64008;
    wire N__64003;
    wire N__63994;
    wire N__63991;
    wire N__63988;
    wire N__63985;
    wire N__63982;
    wire N__63979;
    wire N__63976;
    wire N__63973;
    wire N__63970;
    wire N__63969;
    wire N__63966;
    wire N__63963;
    wire N__63958;
    wire N__63957;
    wire N__63956;
    wire N__63953;
    wire N__63950;
    wire N__63947;
    wire N__63944;
    wire N__63941;
    wire N__63938;
    wire N__63935;
    wire N__63932;
    wire N__63929;
    wire N__63922;
    wire N__63919;
    wire N__63918;
    wire N__63917;
    wire N__63914;
    wire N__63911;
    wire N__63908;
    wire N__63905;
    wire N__63902;
    wire N__63901;
    wire N__63900;
    wire N__63897;
    wire N__63894;
    wire N__63891;
    wire N__63886;
    wire N__63877;
    wire N__63876;
    wire N__63873;
    wire N__63870;
    wire N__63865;
    wire N__63864;
    wire N__63863;
    wire N__63862;
    wire N__63861;
    wire N__63860;
    wire N__63859;
    wire N__63856;
    wire N__63855;
    wire N__63854;
    wire N__63853;
    wire N__63852;
    wire N__63851;
    wire N__63850;
    wire N__63849;
    wire N__63846;
    wire N__63843;
    wire N__63840;
    wire N__63835;
    wire N__63832;
    wire N__63831;
    wire N__63830;
    wire N__63827;
    wire N__63826;
    wire N__63825;
    wire N__63820;
    wire N__63817;
    wire N__63816;
    wire N__63815;
    wire N__63814;
    wire N__63813;
    wire N__63810;
    wire N__63807;
    wire N__63804;
    wire N__63801;
    wire N__63800;
    wire N__63797;
    wire N__63794;
    wire N__63793;
    wire N__63790;
    wire N__63785;
    wire N__63782;
    wire N__63781;
    wire N__63780;
    wire N__63779;
    wire N__63776;
    wire N__63773;
    wire N__63770;
    wire N__63769;
    wire N__63768;
    wire N__63765;
    wire N__63764;
    wire N__63761;
    wire N__63758;
    wire N__63753;
    wire N__63750;
    wire N__63747;
    wire N__63744;
    wire N__63741;
    wire N__63738;
    wire N__63735;
    wire N__63732;
    wire N__63727;
    wire N__63724;
    wire N__63717;
    wire N__63716;
    wire N__63713;
    wire N__63710;
    wire N__63707;
    wire N__63700;
    wire N__63695;
    wire N__63692;
    wire N__63689;
    wire N__63686;
    wire N__63679;
    wire N__63672;
    wire N__63665;
    wire N__63660;
    wire N__63657;
    wire N__63654;
    wire N__63651;
    wire N__63644;
    wire N__63643;
    wire N__63638;
    wire N__63633;
    wire N__63626;
    wire N__63623;
    wire N__63620;
    wire N__63617;
    wire N__63612;
    wire N__63609;
    wire N__63606;
    wire N__63603;
    wire N__63600;
    wire N__63597;
    wire N__63592;
    wire N__63589;
    wire N__63574;
    wire N__63573;
    wire N__63570;
    wire N__63567;
    wire N__63564;
    wire N__63561;
    wire N__63560;
    wire N__63555;
    wire N__63552;
    wire N__63547;
    wire N__63546;
    wire N__63543;
    wire N__63540;
    wire N__63539;
    wire N__63538;
    wire N__63535;
    wire N__63532;
    wire N__63529;
    wire N__63526;
    wire N__63523;
    wire N__63520;
    wire N__63517;
    wire N__63510;
    wire N__63505;
    wire N__63502;
    wire N__63501;
    wire N__63498;
    wire N__63495;
    wire N__63490;
    wire N__63487;
    wire N__63486;
    wire N__63485;
    wire N__63482;
    wire N__63479;
    wire N__63476;
    wire N__63475;
    wire N__63470;
    wire N__63467;
    wire N__63464;
    wire N__63459;
    wire N__63456;
    wire N__63455;
    wire N__63450;
    wire N__63447;
    wire N__63444;
    wire N__63439;
    wire N__63436;
    wire N__63433;
    wire N__63432;
    wire N__63429;
    wire N__63426;
    wire N__63421;
    wire N__63418;
    wire N__63417;
    wire N__63416;
    wire N__63413;
    wire N__63410;
    wire N__63407;
    wire N__63404;
    wire N__63401;
    wire N__63398;
    wire N__63395;
    wire N__63388;
    wire N__63387;
    wire N__63384;
    wire N__63381;
    wire N__63378;
    wire N__63375;
    wire N__63372;
    wire N__63369;
    wire N__63364;
    wire N__63361;
    wire N__63358;
    wire N__63357;
    wire N__63356;
    wire N__63355;
    wire N__63352;
    wire N__63351;
    wire N__63348;
    wire N__63345;
    wire N__63342;
    wire N__63339;
    wire N__63336;
    wire N__63331;
    wire N__63328;
    wire N__63321;
    wire N__63316;
    wire N__63313;
    wire N__63310;
    wire N__63309;
    wire N__63308;
    wire N__63305;
    wire N__63304;
    wire N__63301;
    wire N__63296;
    wire N__63295;
    wire N__63292;
    wire N__63289;
    wire N__63286;
    wire N__63283;
    wire N__63280;
    wire N__63275;
    wire N__63268;
    wire N__63267;
    wire N__63264;
    wire N__63261;
    wire N__63258;
    wire N__63257;
    wire N__63254;
    wire N__63251;
    wire N__63248;
    wire N__63245;
    wire N__63238;
    wire N__63235;
    wire N__63232;
    wire N__63229;
    wire N__63226;
    wire N__63225;
    wire N__63222;
    wire N__63219;
    wire N__63218;
    wire N__63217;
    wire N__63216;
    wire N__63213;
    wire N__63210;
    wire N__63207;
    wire N__63206;
    wire N__63205;
    wire N__63204;
    wire N__63201;
    wire N__63198;
    wire N__63195;
    wire N__63192;
    wire N__63189;
    wire N__63188;
    wire N__63185;
    wire N__63182;
    wire N__63179;
    wire N__63178;
    wire N__63177;
    wire N__63176;
    wire N__63175;
    wire N__63174;
    wire N__63173;
    wire N__63172;
    wire N__63171;
    wire N__63170;
    wire N__63165;
    wire N__63162;
    wire N__63161;
    wire N__63156;
    wire N__63153;
    wire N__63150;
    wire N__63147;
    wire N__63146;
    wire N__63145;
    wire N__63144;
    wire N__63143;
    wire N__63140;
    wire N__63139;
    wire N__63136;
    wire N__63133;
    wire N__63130;
    wire N__63125;
    wire N__63124;
    wire N__63123;
    wire N__63120;
    wire N__63117;
    wire N__63114;
    wire N__63111;
    wire N__63108;
    wire N__63107;
    wire N__63106;
    wire N__63103;
    wire N__63100;
    wire N__63093;
    wire N__63092;
    wire N__63089;
    wire N__63086;
    wire N__63083;
    wire N__63078;
    wire N__63075;
    wire N__63072;
    wire N__63069;
    wire N__63062;
    wire N__63059;
    wire N__63058;
    wire N__63055;
    wire N__63052;
    wire N__63049;
    wire N__63046;
    wire N__63041;
    wire N__63038;
    wire N__63035;
    wire N__63030;
    wire N__63027;
    wire N__63024;
    wire N__63021;
    wire N__63018;
    wire N__63015;
    wire N__63010;
    wire N__63001;
    wire N__63000;
    wire N__62997;
    wire N__62990;
    wire N__62985;
    wire N__62982;
    wire N__62979;
    wire N__62976;
    wire N__62975;
    wire N__62972;
    wire N__62967;
    wire N__62964;
    wire N__62961;
    wire N__62956;
    wire N__62953;
    wire N__62944;
    wire N__62941;
    wire N__62938;
    wire N__62935;
    wire N__62932;
    wire N__62929;
    wire N__62922;
    wire N__62913;
    wire N__62902;
    wire N__62901;
    wire N__62900;
    wire N__62897;
    wire N__62894;
    wire N__62893;
    wire N__62890;
    wire N__62887;
    wire N__62884;
    wire N__62881;
    wire N__62874;
    wire N__62869;
    wire N__62866;
    wire N__62863;
    wire N__62860;
    wire N__62857;
    wire N__62854;
    wire N__62851;
    wire N__62850;
    wire N__62847;
    wire N__62844;
    wire N__62839;
    wire N__62836;
    wire N__62833;
    wire N__62830;
    wire N__62827;
    wire N__62826;
    wire N__62823;
    wire N__62822;
    wire N__62819;
    wire N__62816;
    wire N__62815;
    wire N__62812;
    wire N__62807;
    wire N__62804;
    wire N__62801;
    wire N__62798;
    wire N__62791;
    wire N__62788;
    wire N__62787;
    wire N__62784;
    wire N__62781;
    wire N__62778;
    wire N__62775;
    wire N__62770;
    wire N__62767;
    wire N__62766;
    wire N__62765;
    wire N__62762;
    wire N__62757;
    wire N__62752;
    wire N__62751;
    wire N__62748;
    wire N__62745;
    wire N__62742;
    wire N__62739;
    wire N__62736;
    wire N__62733;
    wire N__62730;
    wire N__62729;
    wire N__62726;
    wire N__62723;
    wire N__62720;
    wire N__62717;
    wire N__62714;
    wire N__62707;
    wire N__62706;
    wire N__62703;
    wire N__62702;
    wire N__62699;
    wire N__62698;
    wire N__62695;
    wire N__62690;
    wire N__62687;
    wire N__62682;
    wire N__62677;
    wire N__62676;
    wire N__62673;
    wire N__62672;
    wire N__62671;
    wire N__62668;
    wire N__62665;
    wire N__62662;
    wire N__62661;
    wire N__62658;
    wire N__62655;
    wire N__62650;
    wire N__62647;
    wire N__62644;
    wire N__62635;
    wire N__62632;
    wire N__62631;
    wire N__62630;
    wire N__62627;
    wire N__62624;
    wire N__62621;
    wire N__62618;
    wire N__62615;
    wire N__62612;
    wire N__62609;
    wire N__62606;
    wire N__62599;
    wire N__62598;
    wire N__62595;
    wire N__62592;
    wire N__62591;
    wire N__62590;
    wire N__62587;
    wire N__62584;
    wire N__62581;
    wire N__62578;
    wire N__62573;
    wire N__62570;
    wire N__62567;
    wire N__62564;
    wire N__62557;
    wire N__62556;
    wire N__62555;
    wire N__62554;
    wire N__62551;
    wire N__62546;
    wire N__62545;
    wire N__62544;
    wire N__62543;
    wire N__62542;
    wire N__62541;
    wire N__62540;
    wire N__62539;
    wire N__62538;
    wire N__62535;
    wire N__62532;
    wire N__62531;
    wire N__62530;
    wire N__62529;
    wire N__62528;
    wire N__62527;
    wire N__62526;
    wire N__62525;
    wire N__62524;
    wire N__62523;
    wire N__62522;
    wire N__62519;
    wire N__62514;
    wire N__62511;
    wire N__62510;
    wire N__62509;
    wire N__62508;
    wire N__62507;
    wire N__62506;
    wire N__62505;
    wire N__62504;
    wire N__62503;
    wire N__62502;
    wire N__62501;
    wire N__62500;
    wire N__62499;
    wire N__62498;
    wire N__62497;
    wire N__62496;
    wire N__62495;
    wire N__62494;
    wire N__62493;
    wire N__62492;
    wire N__62491;
    wire N__62490;
    wire N__62487;
    wire N__62484;
    wire N__62477;
    wire N__62472;
    wire N__62465;
    wire N__62458;
    wire N__62449;
    wire N__62444;
    wire N__62441;
    wire N__62436;
    wire N__62433;
    wire N__62432;
    wire N__62431;
    wire N__62430;
    wire N__62429;
    wire N__62428;
    wire N__62427;
    wire N__62422;
    wire N__62417;
    wire N__62412;
    wire N__62409;
    wire N__62406;
    wire N__62397;
    wire N__62396;
    wire N__62383;
    wire N__62380;
    wire N__62379;
    wire N__62378;
    wire N__62377;
    wire N__62376;
    wire N__62375;
    wire N__62374;
    wire N__62365;
    wire N__62360;
    wire N__62357;
    wire N__62352;
    wire N__62351;
    wire N__62348;
    wire N__62343;
    wire N__62340;
    wire N__62333;
    wire N__62330;
    wire N__62327;
    wire N__62324;
    wire N__62317;
    wire N__62314;
    wire N__62311;
    wire N__62308;
    wire N__62305;
    wire N__62302;
    wire N__62299;
    wire N__62292;
    wire N__62289;
    wire N__62282;
    wire N__62279;
    wire N__62276;
    wire N__62273;
    wire N__62260;
    wire N__62257;
    wire N__62252;
    wire N__62249;
    wire N__62236;
    wire N__62233;
    wire N__62230;
    wire N__62227;
    wire N__62222;
    wire N__62217;
    wire N__62206;
    wire N__62205;
    wire N__62204;
    wire N__62203;
    wire N__62202;
    wire N__62199;
    wire N__62198;
    wire N__62197;
    wire N__62194;
    wire N__62191;
    wire N__62190;
    wire N__62189;
    wire N__62188;
    wire N__62187;
    wire N__62186;
    wire N__62185;
    wire N__62184;
    wire N__62183;
    wire N__62182;
    wire N__62181;
    wire N__62178;
    wire N__62177;
    wire N__62174;
    wire N__62171;
    wire N__62168;
    wire N__62167;
    wire N__62166;
    wire N__62161;
    wire N__62160;
    wire N__62157;
    wire N__62154;
    wire N__62151;
    wire N__62150;
    wire N__62149;
    wire N__62148;
    wire N__62145;
    wire N__62142;
    wire N__62137;
    wire N__62132;
    wire N__62125;
    wire N__62122;
    wire N__62121;
    wire N__62120;
    wire N__62117;
    wire N__62112;
    wire N__62107;
    wire N__62104;
    wire N__62101;
    wire N__62098;
    wire N__62095;
    wire N__62092;
    wire N__62089;
    wire N__62088;
    wire N__62087;
    wire N__62086;
    wire N__62083;
    wire N__62080;
    wire N__62077;
    wire N__62074;
    wire N__62071;
    wire N__62068;
    wire N__62065;
    wire N__62062;
    wire N__62059;
    wire N__62058;
    wire N__62055;
    wire N__62052;
    wire N__62049;
    wire N__62046;
    wire N__62043;
    wire N__62038;
    wire N__62033;
    wire N__62030;
    wire N__62027;
    wire N__62024;
    wire N__62021;
    wire N__62018;
    wire N__62015;
    wire N__62010;
    wire N__62007;
    wire N__62004;
    wire N__62001;
    wire N__61998;
    wire N__61995;
    wire N__61992;
    wire N__61989;
    wire N__61982;
    wire N__61977;
    wire N__61974;
    wire N__61971;
    wire N__61970;
    wire N__61969;
    wire N__61966;
    wire N__61961;
    wire N__61950;
    wire N__61945;
    wire N__61934;
    wire N__61929;
    wire N__61924;
    wire N__61921;
    wire N__61918;
    wire N__61915;
    wire N__61910;
    wire N__61907;
    wire N__61894;
    wire N__61891;
    wire N__61888;
    wire N__61887;
    wire N__61886;
    wire N__61885;
    wire N__61884;
    wire N__61881;
    wire N__61878;
    wire N__61875;
    wire N__61872;
    wire N__61869;
    wire N__61866;
    wire N__61861;
    wire N__61852;
    wire N__61849;
    wire N__61848;
    wire N__61845;
    wire N__61842;
    wire N__61839;
    wire N__61836;
    wire N__61833;
    wire N__61828;
    wire N__61825;
    wire N__61824;
    wire N__61823;
    wire N__61820;
    wire N__61817;
    wire N__61814;
    wire N__61813;
    wire N__61808;
    wire N__61807;
    wire N__61804;
    wire N__61801;
    wire N__61798;
    wire N__61795;
    wire N__61786;
    wire N__61783;
    wire N__61780;
    wire N__61777;
    wire N__61774;
    wire N__61773;
    wire N__61770;
    wire N__61767;
    wire N__61764;
    wire N__61763;
    wire N__61760;
    wire N__61757;
    wire N__61754;
    wire N__61747;
    wire N__61746;
    wire N__61745;
    wire N__61742;
    wire N__61741;
    wire N__61738;
    wire N__61737;
    wire N__61734;
    wire N__61731;
    wire N__61728;
    wire N__61725;
    wire N__61722;
    wire N__61715;
    wire N__61708;
    wire N__61705;
    wire N__61702;
    wire N__61699;
    wire N__61696;
    wire N__61695;
    wire N__61694;
    wire N__61691;
    wire N__61688;
    wire N__61685;
    wire N__61682;
    wire N__61679;
    wire N__61672;
    wire N__61669;
    wire N__61668;
    wire N__61667;
    wire N__61666;
    wire N__61663;
    wire N__61660;
    wire N__61655;
    wire N__61652;
    wire N__61647;
    wire N__61642;
    wire N__61641;
    wire N__61638;
    wire N__61635;
    wire N__61632;
    wire N__61629;
    wire N__61626;
    wire N__61623;
    wire N__61618;
    wire N__61617;
    wire N__61616;
    wire N__61615;
    wire N__61612;
    wire N__61609;
    wire N__61604;
    wire N__61603;
    wire N__61600;
    wire N__61597;
    wire N__61594;
    wire N__61591;
    wire N__61588;
    wire N__61579;
    wire N__61578;
    wire N__61575;
    wire N__61572;
    wire N__61569;
    wire N__61566;
    wire N__61561;
    wire N__61558;
    wire N__61555;
    wire N__61552;
    wire N__61549;
    wire N__61546;
    wire N__61543;
    wire N__61542;
    wire N__61539;
    wire N__61536;
    wire N__61533;
    wire N__61530;
    wire N__61525;
    wire N__61522;
    wire N__61519;
    wire N__61518;
    wire N__61517;
    wire N__61514;
    wire N__61511;
    wire N__61508;
    wire N__61501;
    wire N__61500;
    wire N__61497;
    wire N__61496;
    wire N__61493;
    wire N__61488;
    wire N__61485;
    wire N__61482;
    wire N__61481;
    wire N__61476;
    wire N__61473;
    wire N__61468;
    wire N__61467;
    wire N__61464;
    wire N__61461;
    wire N__61458;
    wire N__61455;
    wire N__61452;
    wire N__61449;
    wire N__61448;
    wire N__61443;
    wire N__61440;
    wire N__61435;
    wire N__61434;
    wire N__61431;
    wire N__61430;
    wire N__61427;
    wire N__61424;
    wire N__61421;
    wire N__61420;
    wire N__61417;
    wire N__61416;
    wire N__61415;
    wire N__61410;
    wire N__61407;
    wire N__61404;
    wire N__61399;
    wire N__61390;
    wire N__61389;
    wire N__61386;
    wire N__61383;
    wire N__61382;
    wire N__61379;
    wire N__61376;
    wire N__61373;
    wire N__61370;
    wire N__61367;
    wire N__61360;
    wire N__61359;
    wire N__61356;
    wire N__61353;
    wire N__61350;
    wire N__61347;
    wire N__61344;
    wire N__61343;
    wire N__61338;
    wire N__61335;
    wire N__61330;
    wire N__61329;
    wire N__61326;
    wire N__61323;
    wire N__61322;
    wire N__61319;
    wire N__61316;
    wire N__61313;
    wire N__61312;
    wire N__61307;
    wire N__61304;
    wire N__61301;
    wire N__61294;
    wire N__61291;
    wire N__61290;
    wire N__61289;
    wire N__61286;
    wire N__61285;
    wire N__61284;
    wire N__61281;
    wire N__61278;
    wire N__61275;
    wire N__61268;
    wire N__61261;
    wire N__61258;
    wire N__61255;
    wire N__61254;
    wire N__61251;
    wire N__61248;
    wire N__61243;
    wire N__61242;
    wire N__61239;
    wire N__61236;
    wire N__61235;
    wire N__61232;
    wire N__61229;
    wire N__61226;
    wire N__61219;
    wire N__61216;
    wire N__61213;
    wire N__61210;
    wire N__61209;
    wire N__61206;
    wire N__61203;
    wire N__61202;
    wire N__61199;
    wire N__61196;
    wire N__61193;
    wire N__61188;
    wire N__61185;
    wire N__61182;
    wire N__61177;
    wire N__61176;
    wire N__61173;
    wire N__61172;
    wire N__61169;
    wire N__61166;
    wire N__61163;
    wire N__61156;
    wire N__61153;
    wire N__61150;
    wire N__61149;
    wire N__61146;
    wire N__61143;
    wire N__61138;
    wire N__61135;
    wire N__61132;
    wire N__61131;
    wire N__61128;
    wire N__61125;
    wire N__61124;
    wire N__61119;
    wire N__61116;
    wire N__61111;
    wire N__61108;
    wire N__61107;
    wire N__61104;
    wire N__61103;
    wire N__61100;
    wire N__61097;
    wire N__61094;
    wire N__61093;
    wire N__61092;
    wire N__61089;
    wire N__61084;
    wire N__61079;
    wire N__61072;
    wire N__61069;
    wire N__61066;
    wire N__61063;
    wire N__61062;
    wire N__61059;
    wire N__61056;
    wire N__61051;
    wire N__61048;
    wire N__61045;
    wire N__61044;
    wire N__61041;
    wire N__61040;
    wire N__61037;
    wire N__61032;
    wire N__61027;
    wire N__61024;
    wire N__61023;
    wire N__61020;
    wire N__61017;
    wire N__61014;
    wire N__61011;
    wire N__61008;
    wire N__61003;
    wire N__61000;
    wire N__60997;
    wire N__60996;
    wire N__60993;
    wire N__60990;
    wire N__60989;
    wire N__60986;
    wire N__60983;
    wire N__60980;
    wire N__60973;
    wire N__60972;
    wire N__60969;
    wire N__60966;
    wire N__60963;
    wire N__60958;
    wire N__60955;
    wire N__60952;
    wire N__60949;
    wire N__60948;
    wire N__60947;
    wire N__60944;
    wire N__60941;
    wire N__60938;
    wire N__60937;
    wire N__60934;
    wire N__60931;
    wire N__60928;
    wire N__60925;
    wire N__60922;
    wire N__60915;
    wire N__60912;
    wire N__60907;
    wire N__60904;
    wire N__60901;
    wire N__60898;
    wire N__60897;
    wire N__60896;
    wire N__60895;
    wire N__60894;
    wire N__60893;
    wire N__60892;
    wire N__60891;
    wire N__60890;
    wire N__60889;
    wire N__60888;
    wire N__60887;
    wire N__60884;
    wire N__60883;
    wire N__60882;
    wire N__60881;
    wire N__60878;
    wire N__60871;
    wire N__60870;
    wire N__60869;
    wire N__60868;
    wire N__60867;
    wire N__60864;
    wire N__60863;
    wire N__60856;
    wire N__60853;
    wire N__60852;
    wire N__60851;
    wire N__60850;
    wire N__60849;
    wire N__60848;
    wire N__60847;
    wire N__60846;
    wire N__60845;
    wire N__60844;
    wire N__60843;
    wire N__60842;
    wire N__60839;
    wire N__60836;
    wire N__60835;
    wire N__60834;
    wire N__60831;
    wire N__60824;
    wire N__60823;
    wire N__60820;
    wire N__60817;
    wire N__60808;
    wire N__60807;
    wire N__60806;
    wire N__60803;
    wire N__60800;
    wire N__60795;
    wire N__60784;
    wire N__60777;
    wire N__60770;
    wire N__60767;
    wire N__60766;
    wire N__60765;
    wire N__60764;
    wire N__60763;
    wire N__60762;
    wire N__60761;
    wire N__60760;
    wire N__60759;
    wire N__60758;
    wire N__60757;
    wire N__60756;
    wire N__60755;
    wire N__60752;
    wire N__60747;
    wire N__60742;
    wire N__60739;
    wire N__60734;
    wire N__60731;
    wire N__60728;
    wire N__60727;
    wire N__60724;
    wire N__60719;
    wire N__60716;
    wire N__60715;
    wire N__60714;
    wire N__60713;
    wire N__60708;
    wire N__60703;
    wire N__60688;
    wire N__60685;
    wire N__60676;
    wire N__60673;
    wire N__60668;
    wire N__60661;
    wire N__60658;
    wire N__60655;
    wire N__60652;
    wire N__60649;
    wire N__60646;
    wire N__60645;
    wire N__60644;
    wire N__60643;
    wire N__60642;
    wire N__60639;
    wire N__60634;
    wire N__60629;
    wire N__60624;
    wire N__60617;
    wire N__60614;
    wire N__60611;
    wire N__60602;
    wire N__60593;
    wire N__60574;
    wire N__60571;
    wire N__60568;
    wire N__60567;
    wire N__60566;
    wire N__60563;
    wire N__60558;
    wire N__60553;
    wire N__60550;
    wire N__60547;
    wire N__60546;
    wire N__60543;
    wire N__60540;
    wire N__60535;
    wire N__60532;
    wire N__60531;
    wire N__60528;
    wire N__60525;
    wire N__60520;
    wire N__60519;
    wire N__60516;
    wire N__60513;
    wire N__60512;
    wire N__60511;
    wire N__60508;
    wire N__60503;
    wire N__60500;
    wire N__60497;
    wire N__60490;
    wire N__60489;
    wire N__60486;
    wire N__60483;
    wire N__60482;
    wire N__60479;
    wire N__60476;
    wire N__60473;
    wire N__60470;
    wire N__60467;
    wire N__60464;
    wire N__60461;
    wire N__60458;
    wire N__60451;
    wire N__60450;
    wire N__60447;
    wire N__60444;
    wire N__60441;
    wire N__60436;
    wire N__60435;
    wire N__60432;
    wire N__60429;
    wire N__60426;
    wire N__60421;
    wire N__60418;
    wire N__60415;
    wire N__60412;
    wire N__60409;
    wire N__60406;
    wire N__60403;
    wire N__60400;
    wire N__60399;
    wire N__60398;
    wire N__60395;
    wire N__60392;
    wire N__60389;
    wire N__60384;
    wire N__60383;
    wire N__60380;
    wire N__60377;
    wire N__60374;
    wire N__60367;
    wire N__60364;
    wire N__60363;
    wire N__60360;
    wire N__60357;
    wire N__60356;
    wire N__60351;
    wire N__60348;
    wire N__60345;
    wire N__60340;
    wire N__60337;
    wire N__60334;
    wire N__60333;
    wire N__60330;
    wire N__60329;
    wire N__60326;
    wire N__60323;
    wire N__60320;
    wire N__60313;
    wire N__60312;
    wire N__60311;
    wire N__60310;
    wire N__60305;
    wire N__60302;
    wire N__60299;
    wire N__60296;
    wire N__60293;
    wire N__60290;
    wire N__60287;
    wire N__60284;
    wire N__60277;
    wire N__60274;
    wire N__60271;
    wire N__60268;
    wire N__60265;
    wire N__60262;
    wire N__60259;
    wire N__60256;
    wire N__60255;
    wire N__60254;
    wire N__60253;
    wire N__60250;
    wire N__60245;
    wire N__60242;
    wire N__60235;
    wire N__60234;
    wire N__60233;
    wire N__60232;
    wire N__60229;
    wire N__60226;
    wire N__60223;
    wire N__60220;
    wire N__60211;
    wire N__60208;
    wire N__60207;
    wire N__60204;
    wire N__60201;
    wire N__60196;
    wire N__60195;
    wire N__60192;
    wire N__60191;
    wire N__60188;
    wire N__60185;
    wire N__60182;
    wire N__60179;
    wire N__60176;
    wire N__60173;
    wire N__60172;
    wire N__60169;
    wire N__60164;
    wire N__60161;
    wire N__60154;
    wire N__60151;
    wire N__60150;
    wire N__60147;
    wire N__60144;
    wire N__60143;
    wire N__60140;
    wire N__60139;
    wire N__60134;
    wire N__60131;
    wire N__60128;
    wire N__60121;
    wire N__60118;
    wire N__60117;
    wire N__60114;
    wire N__60111;
    wire N__60108;
    wire N__60103;
    wire N__60102;
    wire N__60101;
    wire N__60098;
    wire N__60095;
    wire N__60094;
    wire N__60091;
    wire N__60088;
    wire N__60085;
    wire N__60082;
    wire N__60081;
    wire N__60078;
    wire N__60073;
    wire N__60068;
    wire N__60061;
    wire N__60058;
    wire N__60055;
    wire N__60054;
    wire N__60051;
    wire N__60048;
    wire N__60045;
    wire N__60042;
    wire N__60037;
    wire N__60034;
    wire N__60031;
    wire N__60030;
    wire N__60027;
    wire N__60024;
    wire N__60021;
    wire N__60018;
    wire N__60015;
    wire N__60012;
    wire N__60007;
    wire N__60004;
    wire N__60003;
    wire N__60002;
    wire N__59999;
    wire N__59996;
    wire N__59993;
    wire N__59990;
    wire N__59983;
    wire N__59980;
    wire N__59977;
    wire N__59976;
    wire N__59973;
    wire N__59970;
    wire N__59965;
    wire N__59962;
    wire N__59959;
    wire N__59958;
    wire N__59957;
    wire N__59954;
    wire N__59949;
    wire N__59944;
    wire N__59941;
    wire N__59940;
    wire N__59939;
    wire N__59936;
    wire N__59933;
    wire N__59930;
    wire N__59925;
    wire N__59922;
    wire N__59919;
    wire N__59914;
    wire N__59911;
    wire N__59910;
    wire N__59907;
    wire N__59904;
    wire N__59899;
    wire N__59898;
    wire N__59897;
    wire N__59894;
    wire N__59889;
    wire N__59884;
    wire N__59883;
    wire N__59880;
    wire N__59877;
    wire N__59874;
    wire N__59869;
    wire N__59868;
    wire N__59865;
    wire N__59864;
    wire N__59863;
    wire N__59860;
    wire N__59859;
    wire N__59856;
    wire N__59853;
    wire N__59850;
    wire N__59845;
    wire N__59842;
    wire N__59833;
    wire N__59832;
    wire N__59829;
    wire N__59826;
    wire N__59823;
    wire N__59820;
    wire N__59817;
    wire N__59812;
    wire N__59811;
    wire N__59808;
    wire N__59805;
    wire N__59802;
    wire N__59797;
    wire N__59794;
    wire N__59791;
    wire N__59788;
    wire N__59787;
    wire N__59784;
    wire N__59781;
    wire N__59778;
    wire N__59775;
    wire N__59770;
    wire N__59767;
    wire N__59764;
    wire N__59761;
    wire N__59758;
    wire N__59757;
    wire N__59756;
    wire N__59753;
    wire N__59752;
    wire N__59751;
    wire N__59750;
    wire N__59749;
    wire N__59748;
    wire N__59747;
    wire N__59740;
    wire N__59733;
    wire N__59728;
    wire N__59725;
    wire N__59716;
    wire N__59715;
    wire N__59712;
    wire N__59711;
    wire N__59710;
    wire N__59709;
    wire N__59708;
    wire N__59705;
    wire N__59700;
    wire N__59699;
    wire N__59698;
    wire N__59695;
    wire N__59694;
    wire N__59691;
    wire N__59690;
    wire N__59685;
    wire N__59682;
    wire N__59677;
    wire N__59672;
    wire N__59669;
    wire N__59666;
    wire N__59659;
    wire N__59656;
    wire N__59655;
    wire N__59654;
    wire N__59653;
    wire N__59650;
    wire N__59647;
    wire N__59644;
    wire N__59641;
    wire N__59634;
    wire N__59631;
    wire N__59628;
    wire N__59625;
    wire N__59620;
    wire N__59617;
    wire N__59610;
    wire N__59607;
    wire N__59604;
    wire N__59601;
    wire N__59598;
    wire N__59593;
    wire N__59592;
    wire N__59589;
    wire N__59584;
    wire N__59581;
    wire N__59580;
    wire N__59579;
    wire N__59578;
    wire N__59575;
    wire N__59572;
    wire N__59569;
    wire N__59566;
    wire N__59563;
    wire N__59558;
    wire N__59555;
    wire N__59552;
    wire N__59549;
    wire N__59542;
    wire N__59541;
    wire N__59538;
    wire N__59535;
    wire N__59534;
    wire N__59533;
    wire N__59528;
    wire N__59523;
    wire N__59522;
    wire N__59517;
    wire N__59514;
    wire N__59511;
    wire N__59508;
    wire N__59505;
    wire N__59500;
    wire N__59499;
    wire N__59496;
    wire N__59493;
    wire N__59490;
    wire N__59489;
    wire N__59488;
    wire N__59485;
    wire N__59482;
    wire N__59477;
    wire N__59470;
    wire N__59467;
    wire N__59464;
    wire N__59461;
    wire N__59458;
    wire N__59455;
    wire N__59452;
    wire N__59449;
    wire N__59446;
    wire N__59445;
    wire N__59440;
    wire N__59439;
    wire N__59436;
    wire N__59433;
    wire N__59430;
    wire N__59427;
    wire N__59424;
    wire N__59419;
    wire N__59416;
    wire N__59413;
    wire N__59410;
    wire N__59409;
    wire N__59408;
    wire N__59407;
    wire N__59402;
    wire N__59401;
    wire N__59400;
    wire N__59397;
    wire N__59394;
    wire N__59393;
    wire N__59390;
    wire N__59385;
    wire N__59382;
    wire N__59377;
    wire N__59372;
    wire N__59365;
    wire N__59362;
    wire N__59359;
    wire N__59356;
    wire N__59353;
    wire N__59352;
    wire N__59349;
    wire N__59346;
    wire N__59343;
    wire N__59340;
    wire N__59337;
    wire N__59336;
    wire N__59335;
    wire N__59332;
    wire N__59329;
    wire N__59324;
    wire N__59317;
    wire N__59314;
    wire N__59311;
    wire N__59310;
    wire N__59307;
    wire N__59306;
    wire N__59303;
    wire N__59300;
    wire N__59297;
    wire N__59290;
    wire N__59289;
    wire N__59286;
    wire N__59283;
    wire N__59280;
    wire N__59279;
    wire N__59278;
    wire N__59275;
    wire N__59272;
    wire N__59269;
    wire N__59266;
    wire N__59257;
    wire N__59256;
    wire N__59253;
    wire N__59250;
    wire N__59245;
    wire N__59244;
    wire N__59241;
    wire N__59238;
    wire N__59235;
    wire N__59232;
    wire N__59227;
    wire N__59226;
    wire N__59223;
    wire N__59220;
    wire N__59217;
    wire N__59212;
    wire N__59211;
    wire N__59210;
    wire N__59207;
    wire N__59204;
    wire N__59201;
    wire N__59200;
    wire N__59199;
    wire N__59198;
    wire N__59195;
    wire N__59190;
    wire N__59187;
    wire N__59184;
    wire N__59181;
    wire N__59178;
    wire N__59173;
    wire N__59170;
    wire N__59169;
    wire N__59168;
    wire N__59165;
    wire N__59162;
    wire N__59157;
    wire N__59154;
    wire N__59151;
    wire N__59148;
    wire N__59141;
    wire N__59138;
    wire N__59135;
    wire N__59130;
    wire N__59125;
    wire N__59122;
    wire N__59119;
    wire N__59118;
    wire N__59117;
    wire N__59114;
    wire N__59109;
    wire N__59104;
    wire N__59101;
    wire N__59098;
    wire N__59095;
    wire N__59092;
    wire N__59089;
    wire N__59086;
    wire N__59083;
    wire N__59080;
    wire N__59079;
    wire N__59074;
    wire N__59071;
    wire N__59068;
    wire N__59067;
    wire N__59066;
    wire N__59065;
    wire N__59062;
    wire N__59059;
    wire N__59054;
    wire N__59047;
    wire N__59044;
    wire N__59043;
    wire N__59038;
    wire N__59035;
    wire N__59032;
    wire N__59031;
    wire N__59026;
    wire N__59023;
    wire N__59020;
    wire N__59019;
    wire N__59016;
    wire N__59013;
    wire N__59008;
    wire N__59007;
    wire N__59006;
    wire N__59003;
    wire N__59000;
    wire N__58997;
    wire N__58996;
    wire N__58993;
    wire N__58990;
    wire N__58987;
    wire N__58984;
    wire N__58979;
    wire N__58972;
    wire N__58969;
    wire N__58966;
    wire N__58963;
    wire N__58960;
    wire N__58957;
    wire N__58954;
    wire N__58953;
    wire N__58952;
    wire N__58949;
    wire N__58944;
    wire N__58939;
    wire N__58938;
    wire N__58935;
    wire N__58932;
    wire N__58929;
    wire N__58926;
    wire N__58923;
    wire N__58918;
    wire N__58915;
    wire N__58912;
    wire N__58909;
    wire N__58906;
    wire N__58903;
    wire N__58900;
    wire N__58899;
    wire N__58898;
    wire N__58897;
    wire N__58896;
    wire N__58893;
    wire N__58890;
    wire N__58885;
    wire N__58882;
    wire N__58873;
    wire N__58870;
    wire N__58867;
    wire N__58866;
    wire N__58861;
    wire N__58858;
    wire N__58855;
    wire N__58852;
    wire N__58849;
    wire N__58846;
    wire N__58845;
    wire N__58842;
    wire N__58839;
    wire N__58838;
    wire N__58837;
    wire N__58836;
    wire N__58835;
    wire N__58832;
    wire N__58829;
    wire N__58826;
    wire N__58823;
    wire N__58822;
    wire N__58819;
    wire N__58816;
    wire N__58813;
    wire N__58810;
    wire N__58807;
    wire N__58804;
    wire N__58799;
    wire N__58796;
    wire N__58793;
    wire N__58788;
    wire N__58783;
    wire N__58774;
    wire N__58771;
    wire N__58770;
    wire N__58767;
    wire N__58766;
    wire N__58763;
    wire N__58760;
    wire N__58757;
    wire N__58754;
    wire N__58751;
    wire N__58746;
    wire N__58741;
    wire N__58740;
    wire N__58737;
    wire N__58734;
    wire N__58729;
    wire N__58726;
    wire N__58723;
    wire N__58720;
    wire N__58717;
    wire N__58714;
    wire N__58713;
    wire N__58712;
    wire N__58709;
    wire N__58706;
    wire N__58703;
    wire N__58696;
    wire N__58693;
    wire N__58692;
    wire N__58691;
    wire N__58688;
    wire N__58685;
    wire N__58682;
    wire N__58675;
    wire N__58672;
    wire N__58669;
    wire N__58666;
    wire N__58663;
    wire N__58660;
    wire N__58657;
    wire N__58654;
    wire N__58651;
    wire N__58648;
    wire N__58645;
    wire N__58644;
    wire N__58643;
    wire N__58638;
    wire N__58637;
    wire N__58634;
    wire N__58631;
    wire N__58628;
    wire N__58623;
    wire N__58618;
    wire N__58615;
    wire N__58614;
    wire N__58611;
    wire N__58610;
    wire N__58609;
    wire N__58606;
    wire N__58603;
    wire N__58600;
    wire N__58597;
    wire N__58594;
    wire N__58591;
    wire N__58588;
    wire N__58583;
    wire N__58580;
    wire N__58573;
    wire N__58570;
    wire N__58567;
    wire N__58564;
    wire N__58561;
    wire N__58560;
    wire N__58557;
    wire N__58554;
    wire N__58551;
    wire N__58548;
    wire N__58543;
    wire N__58542;
    wire N__58541;
    wire N__58536;
    wire N__58533;
    wire N__58528;
    wire N__58525;
    wire N__58522;
    wire N__58519;
    wire N__58516;
    wire N__58513;
    wire N__58510;
    wire N__58507;
    wire N__58504;
    wire N__58501;
    wire N__58498;
    wire N__58497;
    wire N__58494;
    wire N__58491;
    wire N__58490;
    wire N__58487;
    wire N__58484;
    wire N__58483;
    wire N__58480;
    wire N__58475;
    wire N__58472;
    wire N__58469;
    wire N__58466;
    wire N__58459;
    wire N__58458;
    wire N__58455;
    wire N__58452;
    wire N__58447;
    wire N__58446;
    wire N__58441;
    wire N__58438;
    wire N__58435;
    wire N__58432;
    wire N__58429;
    wire N__58428;
    wire N__58427;
    wire N__58426;
    wire N__58423;
    wire N__58420;
    wire N__58417;
    wire N__58414;
    wire N__58409;
    wire N__58404;
    wire N__58401;
    wire N__58396;
    wire N__58393;
    wire N__58390;
    wire N__58387;
    wire N__58384;
    wire N__58381;
    wire N__58378;
    wire N__58377;
    wire N__58374;
    wire N__58371;
    wire N__58368;
    wire N__58365;
    wire N__58362;
    wire N__58357;
    wire N__58354;
    wire N__58351;
    wire N__58348;
    wire N__58345;
    wire N__58342;
    wire N__58341;
    wire N__58338;
    wire N__58337;
    wire N__58334;
    wire N__58331;
    wire N__58328;
    wire N__58327;
    wire N__58324;
    wire N__58321;
    wire N__58318;
    wire N__58315;
    wire N__58312;
    wire N__58309;
    wire N__58300;
    wire N__58297;
    wire N__58294;
    wire N__58291;
    wire N__58288;
    wire N__58285;
    wire N__58282;
    wire N__58279;
    wire N__58278;
    wire N__58275;
    wire N__58272;
    wire N__58269;
    wire N__58266;
    wire N__58261;
    wire N__58258;
    wire N__58257;
    wire N__58256;
    wire N__58253;
    wire N__58248;
    wire N__58243;
    wire N__58240;
    wire N__58237;
    wire N__58236;
    wire N__58233;
    wire N__58230;
    wire N__58227;
    wire N__58224;
    wire N__58221;
    wire N__58216;
    wire N__58213;
    wire N__58212;
    wire N__58209;
    wire N__58206;
    wire N__58205;
    wire N__58200;
    wire N__58197;
    wire N__58194;
    wire N__58189;
    wire N__58186;
    wire N__58185;
    wire N__58182;
    wire N__58179;
    wire N__58174;
    wire N__58173;
    wire N__58172;
    wire N__58169;
    wire N__58166;
    wire N__58163;
    wire N__58162;
    wire N__58159;
    wire N__58156;
    wire N__58153;
    wire N__58150;
    wire N__58141;
    wire N__58138;
    wire N__58137;
    wire N__58134;
    wire N__58131;
    wire N__58130;
    wire N__58127;
    wire N__58124;
    wire N__58121;
    wire N__58118;
    wire N__58115;
    wire N__58112;
    wire N__58109;
    wire N__58106;
    wire N__58099;
    wire N__58098;
    wire N__58095;
    wire N__58094;
    wire N__58091;
    wire N__58088;
    wire N__58085;
    wire N__58082;
    wire N__58075;
    wire N__58072;
    wire N__58069;
    wire N__58068;
    wire N__58067;
    wire N__58064;
    wire N__58063;
    wire N__58062;
    wire N__58061;
    wire N__58056;
    wire N__58051;
    wire N__58046;
    wire N__58043;
    wire N__58036;
    wire N__58033;
    wire N__58030;
    wire N__58029;
    wire N__58028;
    wire N__58025;
    wire N__58022;
    wire N__58019;
    wire N__58018;
    wire N__58013;
    wire N__58010;
    wire N__58007;
    wire N__58004;
    wire N__57997;
    wire N__57994;
    wire N__57991;
    wire N__57988;
    wire N__57987;
    wire N__57984;
    wire N__57981;
    wire N__57978;
    wire N__57973;
    wire N__57972;
    wire N__57969;
    wire N__57966;
    wire N__57963;
    wire N__57960;
    wire N__57955;
    wire N__57952;
    wire N__57949;
    wire N__57946;
    wire N__57943;
    wire N__57940;
    wire N__57937;
    wire N__57936;
    wire N__57933;
    wire N__57930;
    wire N__57925;
    wire N__57924;
    wire N__57921;
    wire N__57918;
    wire N__57915;
    wire N__57910;
    wire N__57909;
    wire N__57908;
    wire N__57905;
    wire N__57902;
    wire N__57899;
    wire N__57896;
    wire N__57893;
    wire N__57890;
    wire N__57889;
    wire N__57882;
    wire N__57879;
    wire N__57874;
    wire N__57871;
    wire N__57870;
    wire N__57869;
    wire N__57866;
    wire N__57863;
    wire N__57860;
    wire N__57857;
    wire N__57850;
    wire N__57849;
    wire N__57844;
    wire N__57843;
    wire N__57842;
    wire N__57839;
    wire N__57834;
    wire N__57829;
    wire N__57826;
    wire N__57823;
    wire N__57820;
    wire N__57817;
    wire N__57814;
    wire N__57811;
    wire N__57810;
    wire N__57809;
    wire N__57806;
    wire N__57801;
    wire N__57796;
    wire N__57795;
    wire N__57792;
    wire N__57789;
    wire N__57786;
    wire N__57783;
    wire N__57778;
    wire N__57775;
    wire N__57772;
    wire N__57769;
    wire N__57766;
    wire N__57763;
    wire N__57760;
    wire N__57757;
    wire N__57756;
    wire N__57753;
    wire N__57750;
    wire N__57747;
    wire N__57742;
    wire N__57739;
    wire N__57736;
    wire N__57733;
    wire N__57732;
    wire N__57731;
    wire N__57730;
    wire N__57727;
    wire N__57724;
    wire N__57721;
    wire N__57718;
    wire N__57713;
    wire N__57712;
    wire N__57709;
    wire N__57706;
    wire N__57703;
    wire N__57700;
    wire N__57691;
    wire N__57688;
    wire N__57685;
    wire N__57682;
    wire N__57679;
    wire N__57676;
    wire N__57675;
    wire N__57674;
    wire N__57671;
    wire N__57668;
    wire N__57665;
    wire N__57658;
    wire N__57655;
    wire N__57652;
    wire N__57649;
    wire N__57646;
    wire N__57643;
    wire N__57640;
    wire N__57639;
    wire N__57636;
    wire N__57633;
    wire N__57632;
    wire N__57629;
    wire N__57624;
    wire N__57619;
    wire N__57616;
    wire N__57615;
    wire N__57614;
    wire N__57609;
    wire N__57606;
    wire N__57605;
    wire N__57602;
    wire N__57597;
    wire N__57592;
    wire N__57589;
    wire N__57586;
    wire N__57585;
    wire N__57584;
    wire N__57583;
    wire N__57582;
    wire N__57581;
    wire N__57578;
    wire N__57573;
    wire N__57570;
    wire N__57567;
    wire N__57564;
    wire N__57553;
    wire N__57550;
    wire N__57547;
    wire N__57544;
    wire N__57541;
    wire N__57540;
    wire N__57537;
    wire N__57534;
    wire N__57529;
    wire N__57526;
    wire N__57523;
    wire N__57520;
    wire N__57517;
    wire N__57514;
    wire N__57511;
    wire N__57508;
    wire N__57505;
    wire N__57502;
    wire N__57499;
    wire N__57498;
    wire N__57493;
    wire N__57490;
    wire N__57489;
    wire N__57486;
    wire N__57483;
    wire N__57480;
    wire N__57477;
    wire N__57472;
    wire N__57469;
    wire N__57468;
    wire N__57465;
    wire N__57462;
    wire N__57459;
    wire N__57456;
    wire N__57451;
    wire N__57448;
    wire N__57447;
    wire N__57446;
    wire N__57445;
    wire N__57444;
    wire N__57441;
    wire N__57438;
    wire N__57433;
    wire N__57430;
    wire N__57425;
    wire N__57422;
    wire N__57419;
    wire N__57416;
    wire N__57413;
    wire N__57406;
    wire N__57403;
    wire N__57400;
    wire N__57397;
    wire N__57396;
    wire N__57395;
    wire N__57392;
    wire N__57387;
    wire N__57382;
    wire N__57379;
    wire N__57376;
    wire N__57373;
    wire N__57370;
    wire N__57369;
    wire N__57366;
    wire N__57365;
    wire N__57362;
    wire N__57359;
    wire N__57356;
    wire N__57353;
    wire N__57346;
    wire N__57345;
    wire N__57342;
    wire N__57339;
    wire N__57336;
    wire N__57333;
    wire N__57330;
    wire N__57325;
    wire N__57324;
    wire N__57321;
    wire N__57318;
    wire N__57315;
    wire N__57314;
    wire N__57313;
    wire N__57310;
    wire N__57307;
    wire N__57304;
    wire N__57301;
    wire N__57292;
    wire N__57291;
    wire N__57286;
    wire N__57285;
    wire N__57284;
    wire N__57283;
    wire N__57280;
    wire N__57277;
    wire N__57274;
    wire N__57271;
    wire N__57266;
    wire N__57263;
    wire N__57258;
    wire N__57253;
    wire N__57250;
    wire N__57247;
    wire N__57244;
    wire N__57241;
    wire N__57238;
    wire N__57235;
    wire N__57234;
    wire N__57231;
    wire N__57228;
    wire N__57225;
    wire N__57220;
    wire N__57217;
    wire N__57216;
    wire N__57213;
    wire N__57210;
    wire N__57207;
    wire N__57204;
    wire N__57199;
    wire N__57196;
    wire N__57193;
    wire N__57190;
    wire N__57187;
    wire N__57186;
    wire N__57183;
    wire N__57178;
    wire N__57175;
    wire N__57172;
    wire N__57169;
    wire N__57166;
    wire N__57163;
    wire N__57160;
    wire N__57159;
    wire N__57158;
    wire N__57157;
    wire N__57156;
    wire N__57155;
    wire N__57154;
    wire N__57151;
    wire N__57146;
    wire N__57143;
    wire N__57136;
    wire N__57127;
    wire N__57126;
    wire N__57123;
    wire N__57120;
    wire N__57115;
    wire N__57112;
    wire N__57109;
    wire N__57106;
    wire N__57105;
    wire N__57102;
    wire N__57101;
    wire N__57098;
    wire N__57095;
    wire N__57092;
    wire N__57091;
    wire N__57090;
    wire N__57085;
    wire N__57082;
    wire N__57079;
    wire N__57076;
    wire N__57073;
    wire N__57064;
    wire N__57061;
    wire N__57060;
    wire N__57059;
    wire N__57058;
    wire N__57055;
    wire N__57054;
    wire N__57051;
    wire N__57048;
    wire N__57045;
    wire N__57042;
    wire N__57039;
    wire N__57028;
    wire N__57027;
    wire N__57024;
    wire N__57021;
    wire N__57018;
    wire N__57015;
    wire N__57012;
    wire N__57009;
    wire N__57008;
    wire N__57007;
    wire N__57004;
    wire N__57003;
    wire N__57002;
    wire N__56999;
    wire N__56994;
    wire N__56993;
    wire N__56992;
    wire N__56991;
    wire N__56988;
    wire N__56985;
    wire N__56982;
    wire N__56979;
    wire N__56976;
    wire N__56973;
    wire N__56970;
    wire N__56967;
    wire N__56950;
    wire N__56947;
    wire N__56946;
    wire N__56943;
    wire N__56940;
    wire N__56939;
    wire N__56938;
    wire N__56935;
    wire N__56934;
    wire N__56929;
    wire N__56928;
    wire N__56927;
    wire N__56924;
    wire N__56921;
    wire N__56918;
    wire N__56915;
    wire N__56914;
    wire N__56911;
    wire N__56910;
    wire N__56905;
    wire N__56902;
    wire N__56899;
    wire N__56898;
    wire N__56895;
    wire N__56890;
    wire N__56889;
    wire N__56886;
    wire N__56883;
    wire N__56878;
    wire N__56875;
    wire N__56870;
    wire N__56867;
    wire N__56864;
    wire N__56861;
    wire N__56858;
    wire N__56845;
    wire N__56842;
    wire N__56839;
    wire N__56836;
    wire N__56835;
    wire N__56832;
    wire N__56829;
    wire N__56828;
    wire N__56827;
    wire N__56826;
    wire N__56823;
    wire N__56822;
    wire N__56819;
    wire N__56818;
    wire N__56811;
    wire N__56810;
    wire N__56809;
    wire N__56808;
    wire N__56805;
    wire N__56802;
    wire N__56799;
    wire N__56796;
    wire N__56793;
    wire N__56788;
    wire N__56785;
    wire N__56770;
    wire N__56767;
    wire N__56764;
    wire N__56763;
    wire N__56760;
    wire N__56757;
    wire N__56754;
    wire N__56749;
    wire N__56748;
    wire N__56745;
    wire N__56744;
    wire N__56743;
    wire N__56742;
    wire N__56739;
    wire N__56736;
    wire N__56733;
    wire N__56730;
    wire N__56729;
    wire N__56726;
    wire N__56723;
    wire N__56720;
    wire N__56719;
    wire N__56718;
    wire N__56715;
    wire N__56712;
    wire N__56709;
    wire N__56708;
    wire N__56705;
    wire N__56700;
    wire N__56699;
    wire N__56696;
    wire N__56693;
    wire N__56692;
    wire N__56691;
    wire N__56688;
    wire N__56683;
    wire N__56680;
    wire N__56675;
    wire N__56672;
    wire N__56669;
    wire N__56666;
    wire N__56661;
    wire N__56658;
    wire N__56653;
    wire N__56648;
    wire N__56645;
    wire N__56642;
    wire N__56639;
    wire N__56636;
    wire N__56631;
    wire N__56630;
    wire N__56625;
    wire N__56620;
    wire N__56617;
    wire N__56614;
    wire N__56605;
    wire N__56602;
    wire N__56601;
    wire N__56600;
    wire N__56599;
    wire N__56598;
    wire N__56597;
    wire N__56596;
    wire N__56593;
    wire N__56590;
    wire N__56589;
    wire N__56586;
    wire N__56583;
    wire N__56582;
    wire N__56579;
    wire N__56574;
    wire N__56573;
    wire N__56570;
    wire N__56569;
    wire N__56568;
    wire N__56565;
    wire N__56562;
    wire N__56557;
    wire N__56554;
    wire N__56551;
    wire N__56548;
    wire N__56545;
    wire N__56544;
    wire N__56541;
    wire N__56538;
    wire N__56535;
    wire N__56530;
    wire N__56527;
    wire N__56520;
    wire N__56517;
    wire N__56514;
    wire N__56507;
    wire N__56504;
    wire N__56501;
    wire N__56496;
    wire N__56495;
    wire N__56492;
    wire N__56487;
    wire N__56484;
    wire N__56481;
    wire N__56478;
    wire N__56467;
    wire N__56466;
    wire N__56465;
    wire N__56462;
    wire N__56459;
    wire N__56458;
    wire N__56457;
    wire N__56456;
    wire N__56455;
    wire N__56452;
    wire N__56449;
    wire N__56446;
    wire N__56443;
    wire N__56440;
    wire N__56439;
    wire N__56436;
    wire N__56435;
    wire N__56434;
    wire N__56431;
    wire N__56428;
    wire N__56423;
    wire N__56420;
    wire N__56419;
    wire N__56416;
    wire N__56413;
    wire N__56410;
    wire N__56407;
    wire N__56404;
    wire N__56403;
    wire N__56400;
    wire N__56395;
    wire N__56394;
    wire N__56391;
    wire N__56388;
    wire N__56383;
    wire N__56376;
    wire N__56373;
    wire N__56370;
    wire N__56367;
    wire N__56364;
    wire N__56357;
    wire N__56354;
    wire N__56353;
    wire N__56350;
    wire N__56345;
    wire N__56338;
    wire N__56335;
    wire N__56326;
    wire N__56323;
    wire N__56322;
    wire N__56319;
    wire N__56316;
    wire N__56311;
    wire N__56308;
    wire N__56305;
    wire N__56304;
    wire N__56301;
    wire N__56298;
    wire N__56293;
    wire N__56290;
    wire N__56287;
    wire N__56284;
    wire N__56283;
    wire N__56280;
    wire N__56279;
    wire N__56278;
    wire N__56275;
    wire N__56272;
    wire N__56269;
    wire N__56266;
    wire N__56263;
    wire N__56258;
    wire N__56253;
    wire N__56248;
    wire N__56245;
    wire N__56242;
    wire N__56239;
    wire N__56236;
    wire N__56233;
    wire N__56230;
    wire N__56227;
    wire N__56224;
    wire N__56221;
    wire N__56220;
    wire N__56217;
    wire N__56214;
    wire N__56211;
    wire N__56208;
    wire N__56207;
    wire N__56204;
    wire N__56201;
    wire N__56198;
    wire N__56195;
    wire N__56188;
    wire N__56187;
    wire N__56186;
    wire N__56181;
    wire N__56178;
    wire N__56175;
    wire N__56172;
    wire N__56169;
    wire N__56164;
    wire N__56161;
    wire N__56160;
    wire N__56157;
    wire N__56154;
    wire N__56149;
    wire N__56146;
    wire N__56143;
    wire N__56142;
    wire N__56139;
    wire N__56138;
    wire N__56135;
    wire N__56132;
    wire N__56129;
    wire N__56126;
    wire N__56123;
    wire N__56120;
    wire N__56117;
    wire N__56114;
    wire N__56107;
    wire N__56104;
    wire N__56101;
    wire N__56098;
    wire N__56095;
    wire N__56092;
    wire N__56089;
    wire N__56086;
    wire N__56083;
    wire N__56080;
    wire N__56077;
    wire N__56074;
    wire N__56071;
    wire N__56068;
    wire N__56065;
    wire N__56062;
    wire N__56059;
    wire N__56058;
    wire N__56057;
    wire N__56054;
    wire N__56053;
    wire N__56050;
    wire N__56047;
    wire N__56044;
    wire N__56041;
    wire N__56038;
    wire N__56035;
    wire N__56032;
    wire N__56029;
    wire N__56020;
    wire N__56017;
    wire N__56014;
    wire N__56011;
    wire N__56010;
    wire N__56007;
    wire N__56006;
    wire N__56003;
    wire N__56000;
    wire N__55999;
    wire N__55996;
    wire N__55993;
    wire N__55990;
    wire N__55987;
    wire N__55984;
    wire N__55981;
    wire N__55978;
    wire N__55975;
    wire N__55966;
    wire N__55965;
    wire N__55964;
    wire N__55959;
    wire N__55956;
    wire N__55953;
    wire N__55948;
    wire N__55945;
    wire N__55942;
    wire N__55939;
    wire N__55938;
    wire N__55935;
    wire N__55932;
    wire N__55929;
    wire N__55924;
    wire N__55921;
    wire N__55920;
    wire N__55919;
    wire N__55916;
    wire N__55911;
    wire N__55908;
    wire N__55905;
    wire N__55900;
    wire N__55897;
    wire N__55896;
    wire N__55895;
    wire N__55894;
    wire N__55891;
    wire N__55890;
    wire N__55887;
    wire N__55884;
    wire N__55877;
    wire N__55876;
    wire N__55873;
    wire N__55870;
    wire N__55867;
    wire N__55864;
    wire N__55861;
    wire N__55858;
    wire N__55855;
    wire N__55846;
    wire N__55843;
    wire N__55840;
    wire N__55839;
    wire N__55836;
    wire N__55833;
    wire N__55830;
    wire N__55829;
    wire N__55826;
    wire N__55823;
    wire N__55820;
    wire N__55815;
    wire N__55810;
    wire N__55807;
    wire N__55804;
    wire N__55801;
    wire N__55798;
    wire N__55795;
    wire N__55794;
    wire N__55791;
    wire N__55788;
    wire N__55783;
    wire N__55780;
    wire N__55777;
    wire N__55774;
    wire N__55771;
    wire N__55768;
    wire N__55765;
    wire N__55762;
    wire N__55759;
    wire N__55756;
    wire N__55753;
    wire N__55750;
    wire N__55749;
    wire N__55746;
    wire N__55743;
    wire N__55738;
    wire N__55735;
    wire N__55732;
    wire N__55729;
    wire N__55728;
    wire N__55725;
    wire N__55724;
    wire N__55721;
    wire N__55718;
    wire N__55715;
    wire N__55712;
    wire N__55709;
    wire N__55706;
    wire N__55703;
    wire N__55700;
    wire N__55697;
    wire N__55690;
    wire N__55687;
    wire N__55684;
    wire N__55681;
    wire N__55678;
    wire N__55675;
    wire N__55672;
    wire N__55669;
    wire N__55668;
    wire N__55665;
    wire N__55662;
    wire N__55659;
    wire N__55656;
    wire N__55653;
    wire N__55650;
    wire N__55645;
    wire N__55642;
    wire N__55641;
    wire N__55638;
    wire N__55635;
    wire N__55630;
    wire N__55627;
    wire N__55626;
    wire N__55625;
    wire N__55624;
    wire N__55623;
    wire N__55620;
    wire N__55617;
    wire N__55614;
    wire N__55609;
    wire N__55606;
    wire N__55603;
    wire N__55600;
    wire N__55597;
    wire N__55594;
    wire N__55591;
    wire N__55588;
    wire N__55585;
    wire N__55576;
    wire N__55573;
    wire N__55570;
    wire N__55567;
    wire N__55564;
    wire N__55563;
    wire N__55558;
    wire N__55557;
    wire N__55554;
    wire N__55551;
    wire N__55548;
    wire N__55543;
    wire N__55540;
    wire N__55539;
    wire N__55536;
    wire N__55535;
    wire N__55534;
    wire N__55531;
    wire N__55528;
    wire N__55525;
    wire N__55522;
    wire N__55513;
    wire N__55510;
    wire N__55509;
    wire N__55506;
    wire N__55503;
    wire N__55498;
    wire N__55497;
    wire N__55494;
    wire N__55491;
    wire N__55486;
    wire N__55485;
    wire N__55482;
    wire N__55479;
    wire N__55476;
    wire N__55471;
    wire N__55468;
    wire N__55465;
    wire N__55462;
    wire N__55459;
    wire N__55456;
    wire N__55453;
    wire N__55450;
    wire N__55447;
    wire N__55444;
    wire N__55441;
    wire N__55438;
    wire N__55435;
    wire N__55432;
    wire N__55431;
    wire N__55430;
    wire N__55429;
    wire N__55426;
    wire N__55421;
    wire N__55418;
    wire N__55417;
    wire N__55412;
    wire N__55409;
    wire N__55406;
    wire N__55403;
    wire N__55396;
    wire N__55395;
    wire N__55394;
    wire N__55389;
    wire N__55386;
    wire N__55385;
    wire N__55382;
    wire N__55379;
    wire N__55376;
    wire N__55375;
    wire N__55372;
    wire N__55367;
    wire N__55364;
    wire N__55361;
    wire N__55358;
    wire N__55351;
    wire N__55350;
    wire N__55345;
    wire N__55342;
    wire N__55339;
    wire N__55338;
    wire N__55335;
    wire N__55332;
    wire N__55329;
    wire N__55328;
    wire N__55327;
    wire N__55326;
    wire N__55323;
    wire N__55320;
    wire N__55317;
    wire N__55312;
    wire N__55303;
    wire N__55302;
    wire N__55299;
    wire N__55296;
    wire N__55293;
    wire N__55290;
    wire N__55287;
    wire N__55282;
    wire N__55279;
    wire N__55276;
    wire N__55273;
    wire N__55270;
    wire N__55267;
    wire N__55264;
    wire N__55261;
    wire N__55258;
    wire N__55255;
    wire N__55252;
    wire N__55249;
    wire N__55246;
    wire N__55243;
    wire N__55240;
    wire N__55237;
    wire N__55234;
    wire N__55231;
    wire N__55228;
    wire N__55225;
    wire N__55222;
    wire N__55219;
    wire N__55218;
    wire N__55217;
    wire N__55214;
    wire N__55211;
    wire N__55210;
    wire N__55207;
    wire N__55204;
    wire N__55201;
    wire N__55198;
    wire N__55195;
    wire N__55192;
    wire N__55183;
    wire N__55180;
    wire N__55177;
    wire N__55174;
    wire N__55171;
    wire N__55168;
    wire N__55165;
    wire N__55162;
    wire N__55159;
    wire N__55156;
    wire N__55155;
    wire N__55152;
    wire N__55149;
    wire N__55144;
    wire N__55141;
    wire N__55138;
    wire N__55137;
    wire N__55134;
    wire N__55131;
    wire N__55126;
    wire N__55123;
    wire N__55120;
    wire N__55119;
    wire N__55118;
    wire N__55115;
    wire N__55112;
    wire N__55109;
    wire N__55102;
    wire N__55101;
    wire N__55098;
    wire N__55097;
    wire N__55096;
    wire N__55095;
    wire N__55092;
    wire N__55089;
    wire N__55084;
    wire N__55081;
    wire N__55078;
    wire N__55073;
    wire N__55066;
    wire N__55065;
    wire N__55064;
    wire N__55061;
    wire N__55058;
    wire N__55057;
    wire N__55054;
    wire N__55051;
    wire N__55048;
    wire N__55047;
    wire N__55044;
    wire N__55037;
    wire N__55034;
    wire N__55027;
    wire N__55024;
    wire N__55021;
    wire N__55018;
    wire N__55015;
    wire N__55012;
    wire N__55011;
    wire N__55008;
    wire N__55005;
    wire N__55000;
    wire N__54999;
    wire N__54996;
    wire N__54993;
    wire N__54988;
    wire N__54985;
    wire N__54982;
    wire N__54979;
    wire N__54976;
    wire N__54973;
    wire N__54970;
    wire N__54967;
    wire N__54964;
    wire N__54961;
    wire N__54958;
    wire N__54955;
    wire N__54952;
    wire N__54951;
    wire N__54948;
    wire N__54945;
    wire N__54942;
    wire N__54937;
    wire N__54936;
    wire N__54931;
    wire N__54928;
    wire N__54927;
    wire N__54924;
    wire N__54921;
    wire N__54916;
    wire N__54913;
    wire N__54910;
    wire N__54907;
    wire N__54906;
    wire N__54903;
    wire N__54900;
    wire N__54895;
    wire N__54894;
    wire N__54893;
    wire N__54890;
    wire N__54889;
    wire N__54886;
    wire N__54883;
    wire N__54880;
    wire N__54877;
    wire N__54874;
    wire N__54871;
    wire N__54866;
    wire N__54859;
    wire N__54856;
    wire N__54853;
    wire N__54850;
    wire N__54847;
    wire N__54844;
    wire N__54841;
    wire N__54838;
    wire N__54835;
    wire N__54832;
    wire N__54829;
    wire N__54828;
    wire N__54825;
    wire N__54822;
    wire N__54819;
    wire N__54816;
    wire N__54815;
    wire N__54812;
    wire N__54809;
    wire N__54806;
    wire N__54799;
    wire N__54796;
    wire N__54795;
    wire N__54792;
    wire N__54789;
    wire N__54784;
    wire N__54781;
    wire N__54778;
    wire N__54777;
    wire N__54776;
    wire N__54773;
    wire N__54768;
    wire N__54767;
    wire N__54766;
    wire N__54761;
    wire N__54756;
    wire N__54751;
    wire N__54748;
    wire N__54747;
    wire N__54746;
    wire N__54743;
    wire N__54740;
    wire N__54737;
    wire N__54734;
    wire N__54731;
    wire N__54726;
    wire N__54723;
    wire N__54718;
    wire N__54715;
    wire N__54714;
    wire N__54711;
    wire N__54710;
    wire N__54709;
    wire N__54706;
    wire N__54703;
    wire N__54700;
    wire N__54697;
    wire N__54688;
    wire N__54685;
    wire N__54684;
    wire N__54683;
    wire N__54682;
    wire N__54679;
    wire N__54676;
    wire N__54673;
    wire N__54670;
    wire N__54667;
    wire N__54664;
    wire N__54663;
    wire N__54660;
    wire N__54657;
    wire N__54654;
    wire N__54651;
    wire N__54648;
    wire N__54643;
    wire N__54634;
    wire N__54633;
    wire N__54630;
    wire N__54627;
    wire N__54626;
    wire N__54623;
    wire N__54618;
    wire N__54613;
    wire N__54610;
    wire N__54607;
    wire N__54604;
    wire N__54601;
    wire N__54600;
    wire N__54595;
    wire N__54592;
    wire N__54589;
    wire N__54588;
    wire N__54587;
    wire N__54584;
    wire N__54581;
    wire N__54578;
    wire N__54571;
    wire N__54568;
    wire N__54565;
    wire N__54562;
    wire N__54561;
    wire N__54558;
    wire N__54555;
    wire N__54552;
    wire N__54549;
    wire N__54544;
    wire N__54541;
    wire N__54538;
    wire N__54535;
    wire N__54532;
    wire N__54529;
    wire N__54528;
    wire N__54525;
    wire N__54522;
    wire N__54519;
    wire N__54514;
    wire N__54511;
    wire N__54508;
    wire N__54507;
    wire N__54504;
    wire N__54501;
    wire N__54500;
    wire N__54497;
    wire N__54494;
    wire N__54491;
    wire N__54488;
    wire N__54481;
    wire N__54478;
    wire N__54477;
    wire N__54474;
    wire N__54471;
    wire N__54468;
    wire N__54467;
    wire N__54464;
    wire N__54461;
    wire N__54458;
    wire N__54453;
    wire N__54448;
    wire N__54447;
    wire N__54444;
    wire N__54441;
    wire N__54436;
    wire N__54433;
    wire N__54432;
    wire N__54429;
    wire N__54426;
    wire N__54421;
    wire N__54420;
    wire N__54417;
    wire N__54414;
    wire N__54411;
    wire N__54408;
    wire N__54407;
    wire N__54404;
    wire N__54401;
    wire N__54400;
    wire N__54399;
    wire N__54396;
    wire N__54395;
    wire N__54390;
    wire N__54387;
    wire N__54384;
    wire N__54379;
    wire N__54374;
    wire N__54367;
    wire N__54364;
    wire N__54363;
    wire N__54360;
    wire N__54357;
    wire N__54352;
    wire N__54349;
    wire N__54346;
    wire N__54343;
    wire N__54340;
    wire N__54337;
    wire N__54334;
    wire N__54331;
    wire N__54328;
    wire N__54325;
    wire N__54322;
    wire N__54321;
    wire N__54320;
    wire N__54319;
    wire N__54316;
    wire N__54313;
    wire N__54308;
    wire N__54301;
    wire N__54300;
    wire N__54297;
    wire N__54294;
    wire N__54289;
    wire N__54286;
    wire N__54285;
    wire N__54284;
    wire N__54283;
    wire N__54280;
    wire N__54277;
    wire N__54274;
    wire N__54271;
    wire N__54262;
    wire N__54261;
    wire N__54258;
    wire N__54255;
    wire N__54250;
    wire N__54247;
    wire N__54244;
    wire N__54241;
    wire N__54238;
    wire N__54235;
    wire N__54232;
    wire N__54229;
    wire N__54226;
    wire N__54223;
    wire N__54220;
    wire N__54217;
    wire N__54214;
    wire N__54213;
    wire N__54210;
    wire N__54207;
    wire N__54204;
    wire N__54201;
    wire N__54198;
    wire N__54193;
    wire N__54190;
    wire N__54189;
    wire N__54188;
    wire N__54185;
    wire N__54180;
    wire N__54175;
    wire N__54174;
    wire N__54171;
    wire N__54168;
    wire N__54165;
    wire N__54164;
    wire N__54161;
    wire N__54158;
    wire N__54155;
    wire N__54148;
    wire N__54145;
    wire N__54142;
    wire N__54139;
    wire N__54136;
    wire N__54135;
    wire N__54132;
    wire N__54131;
    wire N__54130;
    wire N__54127;
    wire N__54124;
    wire N__54119;
    wire N__54112;
    wire N__54111;
    wire N__54108;
    wire N__54105;
    wire N__54100;
    wire N__54097;
    wire N__54094;
    wire N__54093;
    wire N__54090;
    wire N__54087;
    wire N__54084;
    wire N__54079;
    wire N__54076;
    wire N__54073;
    wire N__54070;
    wire N__54067;
    wire N__54064;
    wire N__54061;
    wire N__54058;
    wire N__54055;
    wire N__54054;
    wire N__54051;
    wire N__54048;
    wire N__54043;
    wire N__54042;
    wire N__54039;
    wire N__54036;
    wire N__54031;
    wire N__54030;
    wire N__54027;
    wire N__54024;
    wire N__54019;
    wire N__54016;
    wire N__54015;
    wire N__54012;
    wire N__54009;
    wire N__54008;
    wire N__54007;
    wire N__54004;
    wire N__54001;
    wire N__53998;
    wire N__53995;
    wire N__53986;
    wire N__53983;
    wire N__53980;
    wire N__53979;
    wire N__53976;
    wire N__53973;
    wire N__53968;
    wire N__53965;
    wire N__53962;
    wire N__53959;
    wire N__53956;
    wire N__53953;
    wire N__53950;
    wire N__53947;
    wire N__53944;
    wire N__53941;
    wire N__53940;
    wire N__53937;
    wire N__53934;
    wire N__53931;
    wire N__53928;
    wire N__53925;
    wire N__53920;
    wire N__53917;
    wire N__53916;
    wire N__53913;
    wire N__53910;
    wire N__53905;
    wire N__53902;
    wire N__53901;
    wire N__53898;
    wire N__53895;
    wire N__53892;
    wire N__53889;
    wire N__53886;
    wire N__53883;
    wire N__53880;
    wire N__53877;
    wire N__53874;
    wire N__53871;
    wire N__53866;
    wire N__53863;
    wire N__53862;
    wire N__53859;
    wire N__53856;
    wire N__53851;
    wire N__53848;
    wire N__53845;
    wire N__53842;
    wire N__53839;
    wire N__53836;
    wire N__53833;
    wire N__53830;
    wire N__53827;
    wire N__53824;
    wire N__53821;
    wire N__53818;
    wire N__53817;
    wire N__53814;
    wire N__53811;
    wire N__53810;
    wire N__53809;
    wire N__53806;
    wire N__53803;
    wire N__53800;
    wire N__53797;
    wire N__53788;
    wire N__53787;
    wire N__53786;
    wire N__53783;
    wire N__53780;
    wire N__53777;
    wire N__53770;
    wire N__53767;
    wire N__53766;
    wire N__53763;
    wire N__53762;
    wire N__53759;
    wire N__53756;
    wire N__53751;
    wire N__53746;
    wire N__53743;
    wire N__53740;
    wire N__53737;
    wire N__53734;
    wire N__53731;
    wire N__53728;
    wire N__53727;
    wire N__53724;
    wire N__53721;
    wire N__53720;
    wire N__53719;
    wire N__53716;
    wire N__53713;
    wire N__53710;
    wire N__53707;
    wire N__53700;
    wire N__53695;
    wire N__53694;
    wire N__53691;
    wire N__53690;
    wire N__53689;
    wire N__53686;
    wire N__53683;
    wire N__53678;
    wire N__53675;
    wire N__53672;
    wire N__53669;
    wire N__53664;
    wire N__53661;
    wire N__53656;
    wire N__53655;
    wire N__53654;
    wire N__53651;
    wire N__53650;
    wire N__53647;
    wire N__53644;
    wire N__53641;
    wire N__53636;
    wire N__53633;
    wire N__53630;
    wire N__53627;
    wire N__53626;
    wire N__53623;
    wire N__53618;
    wire N__53615;
    wire N__53612;
    wire N__53609;
    wire N__53602;
    wire N__53601;
    wire N__53600;
    wire N__53599;
    wire N__53598;
    wire N__53595;
    wire N__53590;
    wire N__53587;
    wire N__53584;
    wire N__53581;
    wire N__53576;
    wire N__53573;
    wire N__53570;
    wire N__53567;
    wire N__53560;
    wire N__53557;
    wire N__53554;
    wire N__53551;
    wire N__53548;
    wire N__53545;
    wire N__53542;
    wire N__53539;
    wire N__53536;
    wire N__53533;
    wire N__53532;
    wire N__53529;
    wire N__53524;
    wire N__53521;
    wire N__53518;
    wire N__53515;
    wire N__53512;
    wire N__53509;
    wire N__53506;
    wire N__53503;
    wire N__53502;
    wire N__53499;
    wire N__53496;
    wire N__53493;
    wire N__53490;
    wire N__53487;
    wire N__53482;
    wire N__53479;
    wire N__53476;
    wire N__53475;
    wire N__53472;
    wire N__53469;
    wire N__53466;
    wire N__53465;
    wire N__53464;
    wire N__53461;
    wire N__53458;
    wire N__53457;
    wire N__53452;
    wire N__53449;
    wire N__53448;
    wire N__53445;
    wire N__53442;
    wire N__53437;
    wire N__53436;
    wire N__53433;
    wire N__53426;
    wire N__53423;
    wire N__53416;
    wire N__53413;
    wire N__53410;
    wire N__53409;
    wire N__53406;
    wire N__53403;
    wire N__53400;
    wire N__53397;
    wire N__53392;
    wire N__53389;
    wire N__53388;
    wire N__53387;
    wire N__53386;
    wire N__53383;
    wire N__53380;
    wire N__53375;
    wire N__53372;
    wire N__53369;
    wire N__53368;
    wire N__53365;
    wire N__53360;
    wire N__53357;
    wire N__53354;
    wire N__53351;
    wire N__53346;
    wire N__53343;
    wire N__53340;
    wire N__53335;
    wire N__53332;
    wire N__53329;
    wire N__53328;
    wire N__53325;
    wire N__53322;
    wire N__53321;
    wire N__53318;
    wire N__53315;
    wire N__53312;
    wire N__53307;
    wire N__53302;
    wire N__53299;
    wire N__53296;
    wire N__53293;
    wire N__53292;
    wire N__53287;
    wire N__53286;
    wire N__53283;
    wire N__53280;
    wire N__53279;
    wire N__53274;
    wire N__53271;
    wire N__53268;
    wire N__53265;
    wire N__53262;
    wire N__53257;
    wire N__53256;
    wire N__53251;
    wire N__53248;
    wire N__53245;
    wire N__53242;
    wire N__53241;
    wire N__53238;
    wire N__53235;
    wire N__53232;
    wire N__53227;
    wire N__53224;
    wire N__53221;
    wire N__53218;
    wire N__53217;
    wire N__53214;
    wire N__53211;
    wire N__53206;
    wire N__53203;
    wire N__53200;
    wire N__53197;
    wire N__53196;
    wire N__53195;
    wire N__53194;
    wire N__53193;
    wire N__53190;
    wire N__53189;
    wire N__53188;
    wire N__53185;
    wire N__53182;
    wire N__53181;
    wire N__53178;
    wire N__53177;
    wire N__53176;
    wire N__53175;
    wire N__53174;
    wire N__53171;
    wire N__53170;
    wire N__53169;
    wire N__53168;
    wire N__53165;
    wire N__53162;
    wire N__53159;
    wire N__53156;
    wire N__53153;
    wire N__53150;
    wire N__53147;
    wire N__53144;
    wire N__53141;
    wire N__53138;
    wire N__53137;
    wire N__53136;
    wire N__53135;
    wire N__53132;
    wire N__53131;
    wire N__53130;
    wire N__53129;
    wire N__53128;
    wire N__53125;
    wire N__53120;
    wire N__53117;
    wire N__53116;
    wire N__53115;
    wire N__53110;
    wire N__53105;
    wire N__53098;
    wire N__53093;
    wire N__53090;
    wire N__53087;
    wire N__53084;
    wire N__53077;
    wire N__53070;
    wire N__53065;
    wire N__53058;
    wire N__53053;
    wire N__53046;
    wire N__53029;
    wire N__53028;
    wire N__53027;
    wire N__53026;
    wire N__53023;
    wire N__53022;
    wire N__53021;
    wire N__53020;
    wire N__53019;
    wire N__53016;
    wire N__53013;
    wire N__53012;
    wire N__53011;
    wire N__53010;
    wire N__53009;
    wire N__53006;
    wire N__53003;
    wire N__53000;
    wire N__52993;
    wire N__52988;
    wire N__52985;
    wire N__52982;
    wire N__52981;
    wire N__52978;
    wire N__52975;
    wire N__52974;
    wire N__52973;
    wire N__52972;
    wire N__52971;
    wire N__52970;
    wire N__52967;
    wire N__52964;
    wire N__52961;
    wire N__52958;
    wire N__52951;
    wire N__52948;
    wire N__52947;
    wire N__52942;
    wire N__52939;
    wire N__52934;
    wire N__52929;
    wire N__52924;
    wire N__52919;
    wire N__52914;
    wire N__52911;
    wire N__52902;
    wire N__52891;
    wire N__52890;
    wire N__52889;
    wire N__52888;
    wire N__52887;
    wire N__52886;
    wire N__52885;
    wire N__52884;
    wire N__52881;
    wire N__52878;
    wire N__52875;
    wire N__52874;
    wire N__52873;
    wire N__52872;
    wire N__52871;
    wire N__52870;
    wire N__52869;
    wire N__52868;
    wire N__52867;
    wire N__52864;
    wire N__52861;
    wire N__52860;
    wire N__52859;
    wire N__52858;
    wire N__52855;
    wire N__52852;
    wire N__52849;
    wire N__52848;
    wire N__52847;
    wire N__52846;
    wire N__52845;
    wire N__52844;
    wire N__52843;
    wire N__52840;
    wire N__52837;
    wire N__52834;
    wire N__52831;
    wire N__52828;
    wire N__52825;
    wire N__52822;
    wire N__52819;
    wire N__52816;
    wire N__52815;
    wire N__52812;
    wire N__52809;
    wire N__52804;
    wire N__52801;
    wire N__52798;
    wire N__52795;
    wire N__52792;
    wire N__52787;
    wire N__52784;
    wire N__52781;
    wire N__52778;
    wire N__52775;
    wire N__52772;
    wire N__52769;
    wire N__52764;
    wire N__52749;
    wire N__52746;
    wire N__52745;
    wire N__52744;
    wire N__52741;
    wire N__52738;
    wire N__52731;
    wire N__52728;
    wire N__52725;
    wire N__52710;
    wire N__52703;
    wire N__52700;
    wire N__52697;
    wire N__52694;
    wire N__52691;
    wire N__52686;
    wire N__52679;
    wire N__52674;
    wire N__52663;
    wire N__52660;
    wire N__52659;
    wire N__52654;
    wire N__52651;
    wire N__52650;
    wire N__52649;
    wire N__52646;
    wire N__52641;
    wire N__52638;
    wire N__52633;
    wire N__52630;
    wire N__52629;
    wire N__52626;
    wire N__52623;
    wire N__52618;
    wire N__52615;
    wire N__52612;
    wire N__52609;
    wire N__52608;
    wire N__52605;
    wire N__52602;
    wire N__52597;
    wire N__52596;
    wire N__52593;
    wire N__52590;
    wire N__52585;
    wire N__52582;
    wire N__52579;
    wire N__52576;
    wire N__52573;
    wire N__52570;
    wire N__52567;
    wire N__52564;
    wire N__52561;
    wire N__52558;
    wire N__52555;
    wire N__52552;
    wire N__52549;
    wire N__52546;
    wire N__52543;
    wire N__52540;
    wire N__52539;
    wire N__52536;
    wire N__52535;
    wire N__52534;
    wire N__52531;
    wire N__52528;
    wire N__52525;
    wire N__52522;
    wire N__52513;
    wire N__52510;
    wire N__52509;
    wire N__52506;
    wire N__52505;
    wire N__52502;
    wire N__52499;
    wire N__52496;
    wire N__52493;
    wire N__52490;
    wire N__52487;
    wire N__52480;
    wire N__52477;
    wire N__52476;
    wire N__52475;
    wire N__52470;
    wire N__52467;
    wire N__52462;
    wire N__52461;
    wire N__52456;
    wire N__52453;
    wire N__52450;
    wire N__52447;
    wire N__52444;
    wire N__52443;
    wire N__52440;
    wire N__52437;
    wire N__52432;
    wire N__52429;
    wire N__52426;
    wire N__52423;
    wire N__52420;
    wire N__52417;
    wire N__52414;
    wire N__52411;
    wire N__52408;
    wire N__52407;
    wire N__52404;
    wire N__52401;
    wire N__52398;
    wire N__52395;
    wire N__52392;
    wire N__52391;
    wire N__52386;
    wire N__52383;
    wire N__52378;
    wire N__52377;
    wire N__52376;
    wire N__52375;
    wire N__52372;
    wire N__52367;
    wire N__52364;
    wire N__52361;
    wire N__52358;
    wire N__52351;
    wire N__52348;
    wire N__52345;
    wire N__52344;
    wire N__52343;
    wire N__52340;
    wire N__52335;
    wire N__52330;
    wire N__52329;
    wire N__52326;
    wire N__52323;
    wire N__52320;
    wire N__52317;
    wire N__52314;
    wire N__52309;
    wire N__52306;
    wire N__52303;
    wire N__52300;
    wire N__52297;
    wire N__52294;
    wire N__52291;
    wire N__52288;
    wire N__52285;
    wire N__52282;
    wire N__52279;
    wire N__52276;
    wire N__52275;
    wire N__52274;
    wire N__52271;
    wire N__52268;
    wire N__52265;
    wire N__52262;
    wire N__52259;
    wire N__52256;
    wire N__52253;
    wire N__52246;
    wire N__52243;
    wire N__52240;
    wire N__52237;
    wire N__52234;
    wire N__52233;
    wire N__52230;
    wire N__52229;
    wire N__52226;
    wire N__52223;
    wire N__52220;
    wire N__52217;
    wire N__52210;
    wire N__52207;
    wire N__52206;
    wire N__52203;
    wire N__52202;
    wire N__52199;
    wire N__52196;
    wire N__52193;
    wire N__52190;
    wire N__52183;
    wire N__52180;
    wire N__52179;
    wire N__52178;
    wire N__52175;
    wire N__52172;
    wire N__52171;
    wire N__52168;
    wire N__52165;
    wire N__52162;
    wire N__52159;
    wire N__52156;
    wire N__52149;
    wire N__52144;
    wire N__52143;
    wire N__52138;
    wire N__52135;
    wire N__52134;
    wire N__52133;
    wire N__52132;
    wire N__52129;
    wire N__52122;
    wire N__52119;
    wire N__52116;
    wire N__52111;
    wire N__52108;
    wire N__52107;
    wire N__52106;
    wire N__52105;
    wire N__52102;
    wire N__52099;
    wire N__52098;
    wire N__52095;
    wire N__52092;
    wire N__52089;
    wire N__52086;
    wire N__52083;
    wire N__52072;
    wire N__52069;
    wire N__52068;
    wire N__52065;
    wire N__52062;
    wire N__52059;
    wire N__52058;
    wire N__52055;
    wire N__52054;
    wire N__52051;
    wire N__52050;
    wire N__52047;
    wire N__52044;
    wire N__52041;
    wire N__52038;
    wire N__52035;
    wire N__52034;
    wire N__52031;
    wire N__52028;
    wire N__52025;
    wire N__52020;
    wire N__52017;
    wire N__52006;
    wire N__52003;
    wire N__52000;
    wire N__51997;
    wire N__51996;
    wire N__51991;
    wire N__51990;
    wire N__51987;
    wire N__51984;
    wire N__51979;
    wire N__51978;
    wire N__51975;
    wire N__51974;
    wire N__51971;
    wire N__51970;
    wire N__51967;
    wire N__51964;
    wire N__51961;
    wire N__51958;
    wire N__51953;
    wire N__51950;
    wire N__51943;
    wire N__51942;
    wire N__51939;
    wire N__51938;
    wire N__51935;
    wire N__51932;
    wire N__51927;
    wire N__51924;
    wire N__51919;
    wire N__51918;
    wire N__51915;
    wire N__51914;
    wire N__51911;
    wire N__51910;
    wire N__51907;
    wire N__51904;
    wire N__51899;
    wire N__51892;
    wire N__51889;
    wire N__51886;
    wire N__51883;
    wire N__51880;
    wire N__51877;
    wire N__51874;
    wire N__51871;
    wire N__51868;
    wire N__51865;
    wire N__51862;
    wire N__51859;
    wire N__51856;
    wire N__51855;
    wire N__51854;
    wire N__51851;
    wire N__51846;
    wire N__51841;
    wire N__51838;
    wire N__51837;
    wire N__51836;
    wire N__51833;
    wire N__51830;
    wire N__51827;
    wire N__51820;
    wire N__51819;
    wire N__51816;
    wire N__51813;
    wire N__51810;
    wire N__51805;
    wire N__51802;
    wire N__51801;
    wire N__51800;
    wire N__51797;
    wire N__51794;
    wire N__51791;
    wire N__51788;
    wire N__51785;
    wire N__51778;
    wire N__51777;
    wire N__51776;
    wire N__51775;
    wire N__51774;
    wire N__51773;
    wire N__51768;
    wire N__51765;
    wire N__51762;
    wire N__51759;
    wire N__51756;
    wire N__51755;
    wire N__51754;
    wire N__51753;
    wire N__51750;
    wire N__51747;
    wire N__51744;
    wire N__51741;
    wire N__51738;
    wire N__51733;
    wire N__51730;
    wire N__51721;
    wire N__51712;
    wire N__51711;
    wire N__51710;
    wire N__51707;
    wire N__51704;
    wire N__51701;
    wire N__51700;
    wire N__51697;
    wire N__51694;
    wire N__51691;
    wire N__51688;
    wire N__51687;
    wire N__51686;
    wire N__51685;
    wire N__51684;
    wire N__51683;
    wire N__51680;
    wire N__51673;
    wire N__51670;
    wire N__51665;
    wire N__51660;
    wire N__51649;
    wire N__51646;
    wire N__51643;
    wire N__51640;
    wire N__51637;
    wire N__51634;
    wire N__51631;
    wire N__51630;
    wire N__51627;
    wire N__51624;
    wire N__51623;
    wire N__51622;
    wire N__51619;
    wire N__51616;
    wire N__51613;
    wire N__51610;
    wire N__51607;
    wire N__51598;
    wire N__51597;
    wire N__51596;
    wire N__51593;
    wire N__51592;
    wire N__51589;
    wire N__51586;
    wire N__51581;
    wire N__51578;
    wire N__51571;
    wire N__51568;
    wire N__51567;
    wire N__51566;
    wire N__51563;
    wire N__51560;
    wire N__51557;
    wire N__51550;
    wire N__51547;
    wire N__51544;
    wire N__51543;
    wire N__51540;
    wire N__51537;
    wire N__51534;
    wire N__51531;
    wire N__51526;
    wire N__51523;
    wire N__51520;
    wire N__51517;
    wire N__51514;
    wire N__51511;
    wire N__51508;
    wire N__51505;
    wire N__51502;
    wire N__51499;
    wire N__51496;
    wire N__51493;
    wire N__51490;
    wire N__51487;
    wire N__51484;
    wire N__51481;
    wire N__51478;
    wire N__51475;
    wire N__51474;
    wire N__51473;
    wire N__51472;
    wire N__51471;
    wire N__51470;
    wire N__51467;
    wire N__51466;
    wire N__51465;
    wire N__51464;
    wire N__51463;
    wire N__51458;
    wire N__51455;
    wire N__51452;
    wire N__51451;
    wire N__51450;
    wire N__51449;
    wire N__51448;
    wire N__51445;
    wire N__51444;
    wire N__51443;
    wire N__51440;
    wire N__51437;
    wire N__51436;
    wire N__51435;
    wire N__51434;
    wire N__51433;
    wire N__51426;
    wire N__51423;
    wire N__51420;
    wire N__51417;
    wire N__51414;
    wire N__51413;
    wire N__51412;
    wire N__51411;
    wire N__51410;
    wire N__51409;
    wire N__51404;
    wire N__51403;
    wire N__51402;
    wire N__51399;
    wire N__51398;
    wire N__51395;
    wire N__51390;
    wire N__51389;
    wire N__51388;
    wire N__51383;
    wire N__51380;
    wire N__51373;
    wire N__51372;
    wire N__51371;
    wire N__51368;
    wire N__51367;
    wire N__51366;
    wire N__51363;
    wire N__51356;
    wire N__51351;
    wire N__51348;
    wire N__51343;
    wire N__51340;
    wire N__51335;
    wire N__51332;
    wire N__51329;
    wire N__51326;
    wire N__51323;
    wire N__51322;
    wire N__51317;
    wire N__51312;
    wire N__51309;
    wire N__51304;
    wire N__51301;
    wire N__51296;
    wire N__51293;
    wire N__51290;
    wire N__51287;
    wire N__51282;
    wire N__51277;
    wire N__51272;
    wire N__51267;
    wire N__51264;
    wire N__51257;
    wire N__51250;
    wire N__51247;
    wire N__51244;
    wire N__51239;
    wire N__51236;
    wire N__51231;
    wire N__51224;
    wire N__51221;
    wire N__51218;
    wire N__51205;
    wire N__51204;
    wire N__51203;
    wire N__51200;
    wire N__51197;
    wire N__51194;
    wire N__51193;
    wire N__51192;
    wire N__51191;
    wire N__51190;
    wire N__51189;
    wire N__51182;
    wire N__51179;
    wire N__51176;
    wire N__51175;
    wire N__51174;
    wire N__51173;
    wire N__51172;
    wire N__51169;
    wire N__51166;
    wire N__51163;
    wire N__51162;
    wire N__51161;
    wire N__51160;
    wire N__51159;
    wire N__51158;
    wire N__51151;
    wire N__51148;
    wire N__51145;
    wire N__51142;
    wire N__51139;
    wire N__51132;
    wire N__51131;
    wire N__51130;
    wire N__51127;
    wire N__51124;
    wire N__51123;
    wire N__51122;
    wire N__51119;
    wire N__51114;
    wire N__51113;
    wire N__51112;
    wire N__51111;
    wire N__51104;
    wire N__51101;
    wire N__51100;
    wire N__51099;
    wire N__51098;
    wire N__51097;
    wire N__51096;
    wire N__51093;
    wire N__51090;
    wire N__51089;
    wire N__51088;
    wire N__51087;
    wire N__51086;
    wire N__51085;
    wire N__51082;
    wire N__51079;
    wire N__51074;
    wire N__51071;
    wire N__51070;
    wire N__51069;
    wire N__51068;
    wire N__51067;
    wire N__51066;
    wire N__51065;
    wire N__51064;
    wire N__51061;
    wire N__51056;
    wire N__51055;
    wire N__51054;
    wire N__51053;
    wire N__51052;
    wire N__51049;
    wire N__51046;
    wire N__51043;
    wire N__51042;
    wire N__51041;
    wire N__51036;
    wire N__51033;
    wire N__51030;
    wire N__51027;
    wire N__51024;
    wire N__51021;
    wire N__51016;
    wire N__51013;
    wire N__51012;
    wire N__51011;
    wire N__51010;
    wire N__51007;
    wire N__51004;
    wire N__51001;
    wire N__50998;
    wire N__50995;
    wire N__50988;
    wire N__50987;
    wire N__50984;
    wire N__50981;
    wire N__50980;
    wire N__50975;
    wire N__50974;
    wire N__50973;
    wire N__50970;
    wire N__50969;
    wire N__50966;
    wire N__50963;
    wire N__50962;
    wire N__50961;
    wire N__50956;
    wire N__50955;
    wire N__50954;
    wire N__50951;
    wire N__50948;
    wire N__50945;
    wire N__50942;
    wire N__50937;
    wire N__50930;
    wire N__50929;
    wire N__50924;
    wire N__50919;
    wire N__50914;
    wire N__50911;
    wire N__50904;
    wire N__50901;
    wire N__50888;
    wire N__50883;
    wire N__50880;
    wire N__50877;
    wire N__50874;
    wire N__50871;
    wire N__50866;
    wire N__50861;
    wire N__50858;
    wire N__50853;
    wire N__50850;
    wire N__50849;
    wire N__50846;
    wire N__50843;
    wire N__50830;
    wire N__50827;
    wire N__50826;
    wire N__50823;
    wire N__50820;
    wire N__50813;
    wire N__50810;
    wire N__50803;
    wire N__50802;
    wire N__50791;
    wire N__50784;
    wire N__50781;
    wire N__50780;
    wire N__50779;
    wire N__50778;
    wire N__50777;
    wire N__50768;
    wire N__50765;
    wire N__50762;
    wire N__50757;
    wire N__50752;
    wire N__50749;
    wire N__50744;
    wire N__50739;
    wire N__50732;
    wire N__50729;
    wire N__50710;
    wire N__50709;
    wire N__50706;
    wire N__50703;
    wire N__50700;
    wire N__50699;
    wire N__50696;
    wire N__50693;
    wire N__50690;
    wire N__50685;
    wire N__50680;
    wire N__50679;
    wire N__50678;
    wire N__50675;
    wire N__50674;
    wire N__50673;
    wire N__50670;
    wire N__50669;
    wire N__50668;
    wire N__50667;
    wire N__50666;
    wire N__50665;
    wire N__50664;
    wire N__50663;
    wire N__50662;
    wire N__50661;
    wire N__50660;
    wire N__50659;
    wire N__50658;
    wire N__50655;
    wire N__50652;
    wire N__50651;
    wire N__50650;
    wire N__50649;
    wire N__50648;
    wire N__50647;
    wire N__50646;
    wire N__50643;
    wire N__50640;
    wire N__50637;
    wire N__50632;
    wire N__50629;
    wire N__50622;
    wire N__50621;
    wire N__50620;
    wire N__50617;
    wire N__50612;
    wire N__50611;
    wire N__50610;
    wire N__50609;
    wire N__50606;
    wire N__50601;
    wire N__50596;
    wire N__50595;
    wire N__50594;
    wire N__50591;
    wire N__50588;
    wire N__50583;
    wire N__50578;
    wire N__50567;
    wire N__50564;
    wire N__50561;
    wire N__50558;
    wire N__50553;
    wire N__50546;
    wire N__50541;
    wire N__50538;
    wire N__50537;
    wire N__50532;
    wire N__50527;
    wire N__50520;
    wire N__50517;
    wire N__50512;
    wire N__50507;
    wire N__50504;
    wire N__50501;
    wire N__50500;
    wire N__50499;
    wire N__50498;
    wire N__50495;
    wire N__50486;
    wire N__50481;
    wire N__50478;
    wire N__50475;
    wire N__50468;
    wire N__50455;
    wire N__50452;
    wire N__50449;
    wire N__50446;
    wire N__50443;
    wire N__50440;
    wire N__50439;
    wire N__50438;
    wire N__50435;
    wire N__50432;
    wire N__50429;
    wire N__50426;
    wire N__50423;
    wire N__50416;
    wire N__50413;
    wire N__50410;
    wire N__50407;
    wire N__50404;
    wire N__50403;
    wire N__50400;
    wire N__50397;
    wire N__50392;
    wire N__50389;
    wire N__50388;
    wire N__50385;
    wire N__50382;
    wire N__50381;
    wire N__50378;
    wire N__50375;
    wire N__50372;
    wire N__50369;
    wire N__50368;
    wire N__50365;
    wire N__50360;
    wire N__50357;
    wire N__50350;
    wire N__50349;
    wire N__50346;
    wire N__50345;
    wire N__50342;
    wire N__50341;
    wire N__50340;
    wire N__50339;
    wire N__50336;
    wire N__50333;
    wire N__50330;
    wire N__50325;
    wire N__50322;
    wire N__50321;
    wire N__50318;
    wire N__50315;
    wire N__50308;
    wire N__50307;
    wire N__50306;
    wire N__50303;
    wire N__50300;
    wire N__50295;
    wire N__50290;
    wire N__50281;
    wire N__50278;
    wire N__50275;
    wire N__50272;
    wire N__50269;
    wire N__50266;
    wire N__50263;
    wire N__50260;
    wire N__50259;
    wire N__50256;
    wire N__50253;
    wire N__50248;
    wire N__50245;
    wire N__50244;
    wire N__50241;
    wire N__50238;
    wire N__50233;
    wire N__50230;
    wire N__50229;
    wire N__50226;
    wire N__50223;
    wire N__50218;
    wire N__50215;
    wire N__50212;
    wire N__50209;
    wire N__50206;
    wire N__50205;
    wire N__50204;
    wire N__50201;
    wire N__50198;
    wire N__50195;
    wire N__50192;
    wire N__50191;
    wire N__50186;
    wire N__50183;
    wire N__50180;
    wire N__50177;
    wire N__50174;
    wire N__50167;
    wire N__50164;
    wire N__50161;
    wire N__50158;
    wire N__50157;
    wire N__50154;
    wire N__50151;
    wire N__50148;
    wire N__50145;
    wire N__50142;
    wire N__50139;
    wire N__50138;
    wire N__50135;
    wire N__50132;
    wire N__50129;
    wire N__50122;
    wire N__50119;
    wire N__50116;
    wire N__50113;
    wire N__50110;
    wire N__50107;
    wire N__50106;
    wire N__50103;
    wire N__50100;
    wire N__50097;
    wire N__50094;
    wire N__50091;
    wire N__50088;
    wire N__50085;
    wire N__50080;
    wire N__50077;
    wire N__50074;
    wire N__50073;
    wire N__50072;
    wire N__50065;
    wire N__50062;
    wire N__50059;
    wire N__50056;
    wire N__50053;
    wire N__50050;
    wire N__50047;
    wire N__50044;
    wire N__50041;
    wire N__50038;
    wire N__50035;
    wire N__50034;
    wire N__50031;
    wire N__50028;
    wire N__50025;
    wire N__50020;
    wire N__50017;
    wire N__50014;
    wire N__50011;
    wire N__50010;
    wire N__50007;
    wire N__50004;
    wire N__50001;
    wire N__49998;
    wire N__49993;
    wire N__49992;
    wire N__49989;
    wire N__49986;
    wire N__49981;
    wire N__49978;
    wire N__49975;
    wire N__49972;
    wire N__49969;
    wire N__49966;
    wire N__49963;
    wire N__49962;
    wire N__49959;
    wire N__49956;
    wire N__49953;
    wire N__49950;
    wire N__49947;
    wire N__49942;
    wire N__49939;
    wire N__49936;
    wire N__49935;
    wire N__49934;
    wire N__49931;
    wire N__49926;
    wire N__49921;
    wire N__49920;
    wire N__49919;
    wire N__49916;
    wire N__49913;
    wire N__49910;
    wire N__49905;
    wire N__49900;
    wire N__49897;
    wire N__49894;
    wire N__49891;
    wire N__49890;
    wire N__49889;
    wire N__49886;
    wire N__49883;
    wire N__49880;
    wire N__49873;
    wire N__49870;
    wire N__49867;
    wire N__49864;
    wire N__49861;
    wire N__49858;
    wire N__49857;
    wire N__49852;
    wire N__49851;
    wire N__49848;
    wire N__49845;
    wire N__49842;
    wire N__49837;
    wire N__49834;
    wire N__49831;
    wire N__49828;
    wire N__49825;
    wire N__49822;
    wire N__49821;
    wire N__49818;
    wire N__49815;
    wire N__49814;
    wire N__49811;
    wire N__49808;
    wire N__49805;
    wire N__49802;
    wire N__49795;
    wire N__49792;
    wire N__49789;
    wire N__49786;
    wire N__49783;
    wire N__49780;
    wire N__49779;
    wire N__49776;
    wire N__49773;
    wire N__49768;
    wire N__49765;
    wire N__49762;
    wire N__49759;
    wire N__49756;
    wire N__49755;
    wire N__49754;
    wire N__49753;
    wire N__49750;
    wire N__49745;
    wire N__49742;
    wire N__49737;
    wire N__49736;
    wire N__49733;
    wire N__49730;
    wire N__49727;
    wire N__49720;
    wire N__49717;
    wire N__49714;
    wire N__49711;
    wire N__49708;
    wire N__49707;
    wire N__49704;
    wire N__49703;
    wire N__49700;
    wire N__49697;
    wire N__49694;
    wire N__49693;
    wire N__49692;
    wire N__49691;
    wire N__49688;
    wire N__49683;
    wire N__49680;
    wire N__49675;
    wire N__49674;
    wire N__49669;
    wire N__49664;
    wire N__49661;
    wire N__49654;
    wire N__49651;
    wire N__49648;
    wire N__49645;
    wire N__49642;
    wire N__49641;
    wire N__49638;
    wire N__49635;
    wire N__49634;
    wire N__49631;
    wire N__49628;
    wire N__49625;
    wire N__49622;
    wire N__49619;
    wire N__49616;
    wire N__49609;
    wire N__49608;
    wire N__49605;
    wire N__49600;
    wire N__49597;
    wire N__49596;
    wire N__49593;
    wire N__49590;
    wire N__49589;
    wire N__49586;
    wire N__49581;
    wire N__49578;
    wire N__49573;
    wire N__49570;
    wire N__49569;
    wire N__49566;
    wire N__49565;
    wire N__49562;
    wire N__49561;
    wire N__49558;
    wire N__49555;
    wire N__49554;
    wire N__49553;
    wire N__49552;
    wire N__49551;
    wire N__49550;
    wire N__49549;
    wire N__49548;
    wire N__49545;
    wire N__49542;
    wire N__49539;
    wire N__49536;
    wire N__49531;
    wire N__49528;
    wire N__49525;
    wire N__49520;
    wire N__49519;
    wire N__49518;
    wire N__49517;
    wire N__49514;
    wire N__49513;
    wire N__49512;
    wire N__49501;
    wire N__49496;
    wire N__49493;
    wire N__49488;
    wire N__49485;
    wire N__49482;
    wire N__49477;
    wire N__49476;
    wire N__49475;
    wire N__49474;
    wire N__49473;
    wire N__49472;
    wire N__49457;
    wire N__49456;
    wire N__49455;
    wire N__49454;
    wire N__49453;
    wire N__49452;
    wire N__49451;
    wire N__49450;
    wire N__49449;
    wire N__49448;
    wire N__49447;
    wire N__49446;
    wire N__49445;
    wire N__49444;
    wire N__49443;
    wire N__49438;
    wire N__49431;
    wire N__49428;
    wire N__49427;
    wire N__49426;
    wire N__49425;
    wire N__49416;
    wire N__49415;
    wire N__49414;
    wire N__49413;
    wire N__49412;
    wire N__49411;
    wire N__49410;
    wire N__49407;
    wire N__49404;
    wire N__49403;
    wire N__49402;
    wire N__49397;
    wire N__49394;
    wire N__49393;
    wire N__49392;
    wire N__49391;
    wire N__49386;
    wire N__49383;
    wire N__49382;
    wire N__49381;
    wire N__49380;
    wire N__49379;
    wire N__49374;
    wire N__49371;
    wire N__49366;
    wire N__49359;
    wire N__49358;
    wire N__49357;
    wire N__49356;
    wire N__49353;
    wire N__49348;
    wire N__49345;
    wire N__49340;
    wire N__49337;
    wire N__49336;
    wire N__49335;
    wire N__49334;
    wire N__49333;
    wire N__49332;
    wire N__49331;
    wire N__49326;
    wire N__49323;
    wire N__49322;
    wire N__49321;
    wire N__49320;
    wire N__49317;
    wire N__49314;
    wire N__49311;
    wire N__49304;
    wire N__49299;
    wire N__49292;
    wire N__49289;
    wire N__49280;
    wire N__49275;
    wire N__49274;
    wire N__49273;
    wire N__49272;
    wire N__49271;
    wire N__49270;
    wire N__49269;
    wire N__49266;
    wire N__49261;
    wire N__49256;
    wire N__49255;
    wire N__49254;
    wire N__49253;
    wire N__49250;
    wire N__49243;
    wire N__49236;
    wire N__49231;
    wire N__49228;
    wire N__49223;
    wire N__49212;
    wire N__49207;
    wire N__49204;
    wire N__49203;
    wire N__49202;
    wire N__49201;
    wire N__49198;
    wire N__49193;
    wire N__49190;
    wire N__49183;
    wire N__49180;
    wire N__49179;
    wire N__49176;
    wire N__49173;
    wire N__49166;
    wire N__49161;
    wire N__49156;
    wire N__49153;
    wire N__49150;
    wire N__49145;
    wire N__49144;
    wire N__49141;
    wire N__49136;
    wire N__49133;
    wire N__49130;
    wire N__49125;
    wire N__49122;
    wire N__49119;
    wire N__49116;
    wire N__49111;
    wire N__49104;
    wire N__49097;
    wire N__49094;
    wire N__49087;
    wire N__49084;
    wire N__49081;
    wire N__49076;
    wire N__49071;
    wire N__49066;
    wire N__49061;
    wire N__49048;
    wire N__49047;
    wire N__49046;
    wire N__49045;
    wire N__49044;
    wire N__49041;
    wire N__49040;
    wire N__49037;
    wire N__49030;
    wire N__49027;
    wire N__49026;
    wire N__49025;
    wire N__49024;
    wire N__49023;
    wire N__49022;
    wire N__49021;
    wire N__49020;
    wire N__49019;
    wire N__49018;
    wire N__49017;
    wire N__49014;
    wire N__49013;
    wire N__49012;
    wire N__49009;
    wire N__49008;
    wire N__49007;
    wire N__49006;
    wire N__49005;
    wire N__49004;
    wire N__49003;
    wire N__49002;
    wire N__49001;
    wire N__49000;
    wire N__48999;
    wire N__48994;
    wire N__48987;
    wire N__48982;
    wire N__48981;
    wire N__48980;
    wire N__48979;
    wire N__48978;
    wire N__48977;
    wire N__48976;
    wire N__48975;
    wire N__48974;
    wire N__48971;
    wire N__48970;
    wire N__48969;
    wire N__48968;
    wire N__48965;
    wire N__48962;
    wire N__48957;
    wire N__48954;
    wire N__48953;
    wire N__48950;
    wire N__48949;
    wire N__48948;
    wire N__48947;
    wire N__48946;
    wire N__48945;
    wire N__48944;
    wire N__48943;
    wire N__48940;
    wire N__48939;
    wire N__48938;
    wire N__48935;
    wire N__48934;
    wire N__48933;
    wire N__48928;
    wire N__48923;
    wire N__48916;
    wire N__48909;
    wire N__48904;
    wire N__48901;
    wire N__48898;
    wire N__48897;
    wire N__48896;
    wire N__48895;
    wire N__48892;
    wire N__48891;
    wire N__48890;
    wire N__48889;
    wire N__48888;
    wire N__48887;
    wire N__48886;
    wire N__48877;
    wire N__48872;
    wire N__48869;
    wire N__48864;
    wire N__48861;
    wire N__48858;
    wire N__48851;
    wire N__48848;
    wire N__48847;
    wire N__48846;
    wire N__48845;
    wire N__48844;
    wire N__48841;
    wire N__48834;
    wire N__48833;
    wire N__48830;
    wire N__48827;
    wire N__48822;
    wire N__48819;
    wire N__48814;
    wire N__48811;
    wire N__48806;
    wire N__48801;
    wire N__48792;
    wire N__48789;
    wire N__48788;
    wire N__48783;
    wire N__48780;
    wire N__48777;
    wire N__48770;
    wire N__48763;
    wire N__48754;
    wire N__48747;
    wire N__48744;
    wire N__48743;
    wire N__48742;
    wire N__48741;
    wire N__48740;
    wire N__48739;
    wire N__48738;
    wire N__48737;
    wire N__48736;
    wire N__48735;
    wire N__48734;
    wire N__48733;
    wire N__48728;
    wire N__48723;
    wire N__48720;
    wire N__48717;
    wire N__48714;
    wire N__48709;
    wire N__48706;
    wire N__48703;
    wire N__48698;
    wire N__48697;
    wire N__48690;
    wire N__48687;
    wire N__48684;
    wire N__48681;
    wire N__48676;
    wire N__48667;
    wire N__48664;
    wire N__48659;
    wire N__48656;
    wire N__48647;
    wire N__48642;
    wire N__48637;
    wire N__48632;
    wire N__48629;
    wire N__48626;
    wire N__48615;
    wire N__48612;
    wire N__48605;
    wire N__48596;
    wire N__48571;
    wire N__48570;
    wire N__48567;
    wire N__48566;
    wire N__48563;
    wire N__48562;
    wire N__48559;
    wire N__48558;
    wire N__48557;
    wire N__48554;
    wire N__48553;
    wire N__48552;
    wire N__48551;
    wire N__48548;
    wire N__48545;
    wire N__48542;
    wire N__48537;
    wire N__48534;
    wire N__48533;
    wire N__48530;
    wire N__48527;
    wire N__48524;
    wire N__48519;
    wire N__48516;
    wire N__48511;
    wire N__48508;
    wire N__48503;
    wire N__48498;
    wire N__48493;
    wire N__48484;
    wire N__48481;
    wire N__48480;
    wire N__48477;
    wire N__48474;
    wire N__48471;
    wire N__48466;
    wire N__48463;
    wire N__48460;
    wire N__48457;
    wire N__48454;
    wire N__48451;
    wire N__48450;
    wire N__48449;
    wire N__48448;
    wire N__48445;
    wire N__48442;
    wire N__48437;
    wire N__48434;
    wire N__48431;
    wire N__48428;
    wire N__48425;
    wire N__48420;
    wire N__48415;
    wire N__48414;
    wire N__48411;
    wire N__48410;
    wire N__48405;
    wire N__48402;
    wire N__48401;
    wire N__48398;
    wire N__48393;
    wire N__48388;
    wire N__48385;
    wire N__48384;
    wire N__48383;
    wire N__48380;
    wire N__48375;
    wire N__48372;
    wire N__48369;
    wire N__48364;
    wire N__48361;
    wire N__48358;
    wire N__48355;
    wire N__48352;
    wire N__48351;
    wire N__48346;
    wire N__48343;
    wire N__48340;
    wire N__48337;
    wire N__48334;
    wire N__48331;
    wire N__48328;
    wire N__48325;
    wire N__48322;
    wire N__48321;
    wire N__48318;
    wire N__48317;
    wire N__48314;
    wire N__48311;
    wire N__48308;
    wire N__48305;
    wire N__48302;
    wire N__48299;
    wire N__48292;
    wire N__48289;
    wire N__48286;
    wire N__48283;
    wire N__48280;
    wire N__48279;
    wire N__48274;
    wire N__48271;
    wire N__48268;
    wire N__48265;
    wire N__48262;
    wire N__48259;
    wire N__48256;
    wire N__48255;
    wire N__48252;
    wire N__48249;
    wire N__48244;
    wire N__48241;
    wire N__48240;
    wire N__48237;
    wire N__48234;
    wire N__48233;
    wire N__48232;
    wire N__48229;
    wire N__48226;
    wire N__48221;
    wire N__48216;
    wire N__48213;
    wire N__48208;
    wire N__48205;
    wire N__48204;
    wire N__48201;
    wire N__48198;
    wire N__48197;
    wire N__48196;
    wire N__48193;
    wire N__48190;
    wire N__48185;
    wire N__48182;
    wire N__48177;
    wire N__48172;
    wire N__48171;
    wire N__48170;
    wire N__48169;
    wire N__48168;
    wire N__48165;
    wire N__48162;
    wire N__48159;
    wire N__48158;
    wire N__48155;
    wire N__48154;
    wire N__48153;
    wire N__48150;
    wire N__48145;
    wire N__48140;
    wire N__48139;
    wire N__48134;
    wire N__48131;
    wire N__48128;
    wire N__48125;
    wire N__48122;
    wire N__48119;
    wire N__48116;
    wire N__48113;
    wire N__48108;
    wire N__48101;
    wire N__48094;
    wire N__48091;
    wire N__48090;
    wire N__48089;
    wire N__48088;
    wire N__48081;
    wire N__48078;
    wire N__48075;
    wire N__48072;
    wire N__48069;
    wire N__48066;
    wire N__48063;
    wire N__48058;
    wire N__48055;
    wire N__48052;
    wire N__48049;
    wire N__48048;
    wire N__48047;
    wire N__48046;
    wire N__48043;
    wire N__48040;
    wire N__48037;
    wire N__48034;
    wire N__48029;
    wire N__48028;
    wire N__48027;
    wire N__48026;
    wire N__48023;
    wire N__48018;
    wire N__48015;
    wire N__48010;
    wire N__48001;
    wire N__47998;
    wire N__47997;
    wire N__47994;
    wire N__47993;
    wire N__47992;
    wire N__47989;
    wire N__47986;
    wire N__47983;
    wire N__47980;
    wire N__47971;
    wire N__47968;
    wire N__47967;
    wire N__47962;
    wire N__47959;
    wire N__47956;
    wire N__47953;
    wire N__47950;
    wire N__47949;
    wire N__47946;
    wire N__47943;
    wire N__47938;
    wire N__47937;
    wire N__47934;
    wire N__47931;
    wire N__47930;
    wire N__47927;
    wire N__47924;
    wire N__47921;
    wire N__47918;
    wire N__47911;
    wire N__47908;
    wire N__47907;
    wire N__47906;
    wire N__47903;
    wire N__47902;
    wire N__47901;
    wire N__47898;
    wire N__47895;
    wire N__47892;
    wire N__47889;
    wire N__47884;
    wire N__47883;
    wire N__47880;
    wire N__47877;
    wire N__47874;
    wire N__47871;
    wire N__47868;
    wire N__47865;
    wire N__47860;
    wire N__47857;
    wire N__47848;
    wire N__47845;
    wire N__47844;
    wire N__47841;
    wire N__47838;
    wire N__47835;
    wire N__47830;
    wire N__47827;
    wire N__47824;
    wire N__47823;
    wire N__47820;
    wire N__47817;
    wire N__47814;
    wire N__47809;
    wire N__47806;
    wire N__47803;
    wire N__47802;
    wire N__47799;
    wire N__47796;
    wire N__47793;
    wire N__47788;
    wire N__47787;
    wire N__47784;
    wire N__47781;
    wire N__47778;
    wire N__47775;
    wire N__47772;
    wire N__47767;
    wire N__47766;
    wire N__47763;
    wire N__47762;
    wire N__47759;
    wire N__47758;
    wire N__47755;
    wire N__47752;
    wire N__47749;
    wire N__47746;
    wire N__47737;
    wire N__47736;
    wire N__47733;
    wire N__47730;
    wire N__47727;
    wire N__47726;
    wire N__47725;
    wire N__47722;
    wire N__47719;
    wire N__47714;
    wire N__47707;
    wire N__47704;
    wire N__47701;
    wire N__47700;
    wire N__47697;
    wire N__47694;
    wire N__47693;
    wire N__47690;
    wire N__47689;
    wire N__47688;
    wire N__47685;
    wire N__47684;
    wire N__47681;
    wire N__47678;
    wire N__47675;
    wire N__47672;
    wire N__47669;
    wire N__47664;
    wire N__47661;
    wire N__47656;
    wire N__47651;
    wire N__47644;
    wire N__47641;
    wire N__47640;
    wire N__47637;
    wire N__47634;
    wire N__47633;
    wire N__47632;
    wire N__47631;
    wire N__47628;
    wire N__47625;
    wire N__47624;
    wire N__47623;
    wire N__47620;
    wire N__47617;
    wire N__47616;
    wire N__47615;
    wire N__47612;
    wire N__47607;
    wire N__47604;
    wire N__47601;
    wire N__47596;
    wire N__47591;
    wire N__47578;
    wire N__47575;
    wire N__47572;
    wire N__47569;
    wire N__47566;
    wire N__47563;
    wire N__47560;
    wire N__47557;
    wire N__47554;
    wire N__47551;
    wire N__47548;
    wire N__47547;
    wire N__47544;
    wire N__47541;
    wire N__47540;
    wire N__47539;
    wire N__47536;
    wire N__47529;
    wire N__47524;
    wire N__47523;
    wire N__47522;
    wire N__47519;
    wire N__47516;
    wire N__47513;
    wire N__47510;
    wire N__47509;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47501;
    wire N__47500;
    wire N__47497;
    wire N__47494;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47479;
    wire N__47476;
    wire N__47473;
    wire N__47468;
    wire N__47455;
    wire N__47454;
    wire N__47451;
    wire N__47450;
    wire N__47447;
    wire N__47446;
    wire N__47443;
    wire N__47440;
    wire N__47437;
    wire N__47434;
    wire N__47431;
    wire N__47422;
    wire N__47419;
    wire N__47416;
    wire N__47413;
    wire N__47410;
    wire N__47407;
    wire N__47404;
    wire N__47401;
    wire N__47398;
    wire N__47395;
    wire N__47392;
    wire N__47391;
    wire N__47388;
    wire N__47385;
    wire N__47384;
    wire N__47381;
    wire N__47380;
    wire N__47377;
    wire N__47374;
    wire N__47371;
    wire N__47368;
    wire N__47359;
    wire N__47356;
    wire N__47355;
    wire N__47352;
    wire N__47349;
    wire N__47348;
    wire N__47347;
    wire N__47342;
    wire N__47339;
    wire N__47336;
    wire N__47333;
    wire N__47326;
    wire N__47323;
    wire N__47322;
    wire N__47321;
    wire N__47320;
    wire N__47317;
    wire N__47314;
    wire N__47311;
    wire N__47308;
    wire N__47305;
    wire N__47300;
    wire N__47297;
    wire N__47294;
    wire N__47291;
    wire N__47288;
    wire N__47283;
    wire N__47280;
    wire N__47277;
    wire N__47274;
    wire N__47271;
    wire N__47266;
    wire N__47263;
    wire N__47260;
    wire N__47257;
    wire N__47254;
    wire N__47253;
    wire N__47250;
    wire N__47247;
    wire N__47246;
    wire N__47243;
    wire N__47240;
    wire N__47239;
    wire N__47236;
    wire N__47233;
    wire N__47230;
    wire N__47227;
    wire N__47218;
    wire N__47217;
    wire N__47216;
    wire N__47215;
    wire N__47214;
    wire N__47213;
    wire N__47212;
    wire N__47211;
    wire N__47210;
    wire N__47209;
    wire N__47208;
    wire N__47207;
    wire N__47206;
    wire N__47203;
    wire N__47202;
    wire N__47199;
    wire N__47198;
    wire N__47195;
    wire N__47194;
    wire N__47191;
    wire N__47190;
    wire N__47189;
    wire N__47186;
    wire N__47185;
    wire N__47182;
    wire N__47181;
    wire N__47178;
    wire N__47177;
    wire N__47176;
    wire N__47173;
    wire N__47172;
    wire N__47169;
    wire N__47168;
    wire N__47165;
    wire N__47164;
    wire N__47163;
    wire N__47160;
    wire N__47159;
    wire N__47156;
    wire N__47155;
    wire N__47152;
    wire N__47151;
    wire N__47150;
    wire N__47149;
    wire N__47148;
    wire N__47147;
    wire N__47146;
    wire N__47145;
    wire N__47144;
    wire N__47143;
    wire N__47142;
    wire N__47141;
    wire N__47140;
    wire N__47139;
    wire N__47136;
    wire N__47121;
    wire N__47106;
    wire N__47091;
    wire N__47076;
    wire N__47075;
    wire N__47072;
    wire N__47071;
    wire N__47068;
    wire N__47067;
    wire N__47064;
    wire N__47063;
    wire N__47062;
    wire N__47059;
    wire N__47058;
    wire N__47055;
    wire N__47054;
    wire N__47051;
    wire N__47050;
    wire N__47049;
    wire N__47046;
    wire N__47045;
    wire N__47042;
    wire N__47041;
    wire N__47038;
    wire N__47037;
    wire N__47036;
    wire N__47033;
    wire N__47032;
    wire N__47029;
    wire N__47028;
    wire N__47025;
    wire N__47024;
    wire N__47023;
    wire N__47022;
    wire N__47021;
    wire N__47020;
    wire N__47019;
    wire N__47018;
    wire N__47017;
    wire N__47016;
    wire N__47015;
    wire N__47014;
    wire N__47013;
    wire N__47012;
    wire N__47003;
    wire N__47000;
    wire N__46985;
    wire N__46970;
    wire N__46955;
    wire N__46940;
    wire N__46939;
    wire N__46936;
    wire N__46935;
    wire N__46932;
    wire N__46931;
    wire N__46928;
    wire N__46927;
    wire N__46926;
    wire N__46923;
    wire N__46922;
    wire N__46919;
    wire N__46918;
    wire N__46915;
    wire N__46914;
    wire N__46913;
    wire N__46910;
    wire N__46909;
    wire N__46906;
    wire N__46905;
    wire N__46902;
    wire N__46901;
    wire N__46900;
    wire N__46897;
    wire N__46896;
    wire N__46893;
    wire N__46892;
    wire N__46889;
    wire N__46888;
    wire N__46887;
    wire N__46886;
    wire N__46885;
    wire N__46884;
    wire N__46883;
    wire N__46882;
    wire N__46881;
    wire N__46880;
    wire N__46879;
    wire N__46878;
    wire N__46877;
    wire N__46876;
    wire N__46865;
    wire N__46862;
    wire N__46847;
    wire N__46832;
    wire N__46817;
    wire N__46802;
    wire N__46801;
    wire N__46798;
    wire N__46797;
    wire N__46794;
    wire N__46793;
    wire N__46790;
    wire N__46789;
    wire N__46788;
    wire N__46785;
    wire N__46784;
    wire N__46781;
    wire N__46780;
    wire N__46777;
    wire N__46776;
    wire N__46775;
    wire N__46772;
    wire N__46771;
    wire N__46768;
    wire N__46767;
    wire N__46764;
    wire N__46763;
    wire N__46762;
    wire N__46759;
    wire N__46758;
    wire N__46755;
    wire N__46754;
    wire N__46751;
    wire N__46750;
    wire N__46749;
    wire N__46748;
    wire N__46747;
    wire N__46746;
    wire N__46745;
    wire N__46744;
    wire N__46743;
    wire N__46742;
    wire N__46741;
    wire N__46730;
    wire N__46727;
    wire N__46712;
    wire N__46697;
    wire N__46682;
    wire N__46667;
    wire N__46666;
    wire N__46663;
    wire N__46662;
    wire N__46659;
    wire N__46658;
    wire N__46655;
    wire N__46654;
    wire N__46653;
    wire N__46650;
    wire N__46649;
    wire N__46646;
    wire N__46645;
    wire N__46642;
    wire N__46641;
    wire N__46640;
    wire N__46637;
    wire N__46636;
    wire N__46633;
    wire N__46632;
    wire N__46629;
    wire N__46628;
    wire N__46627;
    wire N__46626;
    wire N__46625;
    wire N__46624;
    wire N__46623;
    wire N__46622;
    wire N__46621;
    wire N__46620;
    wire N__46619;
    wire N__46618;
    wire N__46617;
    wire N__46616;
    wire N__46603;
    wire N__46588;
    wire N__46573;
    wire N__46558;
    wire N__46557;
    wire N__46554;
    wire N__46553;
    wire N__46550;
    wire N__46549;
    wire N__46546;
    wire N__46545;
    wire N__46544;
    wire N__46541;
    wire N__46540;
    wire N__46537;
    wire N__46536;
    wire N__46533;
    wire N__46532;
    wire N__46531;
    wire N__46530;
    wire N__46529;
    wire N__46528;
    wire N__46527;
    wire N__46526;
    wire N__46525;
    wire N__46524;
    wire N__46523;
    wire N__46522;
    wire N__46521;
    wire N__46520;
    wire N__46519;
    wire N__46518;
    wire N__46517;
    wire N__46516;
    wire N__46515;
    wire N__46514;
    wire N__46513;
    wire N__46512;
    wire N__46511;
    wire N__46510;
    wire N__46509;
    wire N__46508;
    wire N__46507;
    wire N__46504;
    wire N__46503;
    wire N__46500;
    wire N__46499;
    wire N__46496;
    wire N__46495;
    wire N__46494;
    wire N__46493;
    wire N__46492;
    wire N__46491;
    wire N__46488;
    wire N__46487;
    wire N__46484;
    wire N__46483;
    wire N__46480;
    wire N__46479;
    wire N__46470;
    wire N__46455;
    wire N__46440;
    wire N__46433;
    wire N__46424;
    wire N__46417;
    wire N__46408;
    wire N__46401;
    wire N__46392;
    wire N__46391;
    wire N__46388;
    wire N__46387;
    wire N__46384;
    wire N__46383;
    wire N__46380;
    wire N__46379;
    wire N__46364;
    wire N__46363;
    wire N__46360;
    wire N__46359;
    wire N__46356;
    wire N__46355;
    wire N__46352;
    wire N__46351;
    wire N__46336;
    wire N__46329;
    wire N__46316;
    wire N__46301;
    wire N__46298;
    wire N__46283;
    wire N__46282;
    wire N__46281;
    wire N__46280;
    wire N__46279;
    wire N__46278;
    wire N__46277;
    wire N__46276;
    wire N__46275;
    wire N__46274;
    wire N__46273;
    wire N__46272;
    wire N__46271;
    wire N__46270;
    wire N__46269;
    wire N__46268;
    wire N__46267;
    wire N__46266;
    wire N__46265;
    wire N__46264;
    wire N__46263;
    wire N__46262;
    wire N__46259;
    wire N__46252;
    wire N__46247;
    wire N__46240;
    wire N__46231;
    wire N__46224;
    wire N__46215;
    wire N__46208;
    wire N__46199;
    wire N__46180;
    wire N__46177;
    wire N__46176;
    wire N__46175;
    wire N__46174;
    wire N__46171;
    wire N__46168;
    wire N__46165;
    wire N__46162;
    wire N__46159;
    wire N__46158;
    wire N__46155;
    wire N__46152;
    wire N__46149;
    wire N__46148;
    wire N__46147;
    wire N__46144;
    wire N__46141;
    wire N__46138;
    wire N__46135;
    wire N__46132;
    wire N__46129;
    wire N__46126;
    wire N__46121;
    wire N__46116;
    wire N__46113;
    wire N__46110;
    wire N__46109;
    wire N__46104;
    wire N__46099;
    wire N__46096;
    wire N__46093;
    wire N__46090;
    wire N__46087;
    wire N__46084;
    wire N__46075;
    wire N__46072;
    wire N__46069;
    wire N__46066;
    wire N__46063;
    wire N__46060;
    wire N__46057;
    wire N__46054;
    wire N__46051;
    wire N__46050;
    wire N__46049;
    wire N__46048;
    wire N__46045;
    wire N__46040;
    wire N__46039;
    wire N__46036;
    wire N__46031;
    wire N__46030;
    wire N__46027;
    wire N__46024;
    wire N__46021;
    wire N__46018;
    wire N__46015;
    wire N__46014;
    wire N__46011;
    wire N__46006;
    wire N__46003;
    wire N__46000;
    wire N__45999;
    wire N__45996;
    wire N__45993;
    wire N__45990;
    wire N__45987;
    wire N__45984;
    wire N__45981;
    wire N__45978;
    wire N__45975;
    wire N__45964;
    wire N__45961;
    wire N__45958;
    wire N__45955;
    wire N__45952;
    wire N__45949;
    wire N__45946;
    wire N__45943;
    wire N__45942;
    wire N__45937;
    wire N__45936;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45922;
    wire N__45919;
    wire N__45916;
    wire N__45913;
    wire N__45910;
    wire N__45907;
    wire N__45904;
    wire N__45903;
    wire N__45900;
    wire N__45897;
    wire N__45896;
    wire N__45891;
    wire N__45888;
    wire N__45885;
    wire N__45880;
    wire N__45877;
    wire N__45876;
    wire N__45873;
    wire N__45870;
    wire N__45869;
    wire N__45866;
    wire N__45863;
    wire N__45860;
    wire N__45857;
    wire N__45850;
    wire N__45847;
    wire N__45844;
    wire N__45841;
    wire N__45838;
    wire N__45837;
    wire N__45834;
    wire N__45831;
    wire N__45830;
    wire N__45827;
    wire N__45824;
    wire N__45821;
    wire N__45818;
    wire N__45811;
    wire N__45808;
    wire N__45805;
    wire N__45802;
    wire N__45799;
    wire N__45798;
    wire N__45795;
    wire N__45792;
    wire N__45791;
    wire N__45788;
    wire N__45785;
    wire N__45782;
    wire N__45779;
    wire N__45772;
    wire N__45769;
    wire N__45766;
    wire N__45763;
    wire N__45760;
    wire N__45759;
    wire N__45756;
    wire N__45753;
    wire N__45750;
    wire N__45749;
    wire N__45746;
    wire N__45743;
    wire N__45740;
    wire N__45737;
    wire N__45730;
    wire N__45727;
    wire N__45724;
    wire N__45721;
    wire N__45718;
    wire N__45715;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45707;
    wire N__45704;
    wire N__45701;
    wire N__45698;
    wire N__45695;
    wire N__45688;
    wire N__45685;
    wire N__45682;
    wire N__45679;
    wire N__45676;
    wire N__45675;
    wire N__45674;
    wire N__45671;
    wire N__45668;
    wire N__45665;
    wire N__45662;
    wire N__45655;
    wire N__45652;
    wire N__45649;
    wire N__45646;
    wire N__45643;
    wire N__45640;
    wire N__45637;
    wire N__45634;
    wire N__45631;
    wire N__45630;
    wire N__45629;
    wire N__45626;
    wire N__45623;
    wire N__45620;
    wire N__45613;
    wire N__45610;
    wire N__45607;
    wire N__45604;
    wire N__45601;
    wire N__45598;
    wire N__45595;
    wire N__45592;
    wire N__45589;
    wire N__45586;
    wire N__45583;
    wire N__45580;
    wire N__45579;
    wire N__45576;
    wire N__45573;
    wire N__45570;
    wire N__45569;
    wire N__45566;
    wire N__45563;
    wire N__45560;
    wire N__45557;
    wire N__45550;
    wire N__45547;
    wire N__45544;
    wire N__45541;
    wire N__45538;
    wire N__45535;
    wire N__45534;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45524;
    wire N__45521;
    wire N__45518;
    wire N__45515;
    wire N__45512;
    wire N__45505;
    wire N__45502;
    wire N__45499;
    wire N__45498;
    wire N__45495;
    wire N__45492;
    wire N__45491;
    wire N__45488;
    wire N__45485;
    wire N__45482;
    wire N__45477;
    wire N__45472;
    wire N__45469;
    wire N__45466;
    wire N__45463;
    wire N__45460;
    wire N__45457;
    wire N__45454;
    wire N__45451;
    wire N__45448;
    wire N__45445;
    wire N__45442;
    wire N__45439;
    wire N__45436;
    wire N__45435;
    wire N__45432;
    wire N__45429;
    wire N__45426;
    wire N__45425;
    wire N__45422;
    wire N__45419;
    wire N__45416;
    wire N__45413;
    wire N__45406;
    wire N__45403;
    wire N__45400;
    wire N__45397;
    wire N__45394;
    wire N__45391;
    wire N__45388;
    wire N__45385;
    wire N__45384;
    wire N__45381;
    wire N__45378;
    wire N__45375;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45363;
    wire N__45362;
    wire N__45359;
    wire N__45356;
    wire N__45353;
    wire N__45346;
    wire N__45343;
    wire N__45340;
    wire N__45337;
    wire N__45334;
    wire N__45331;
    wire N__45328;
    wire N__45327;
    wire N__45324;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45314;
    wire N__45309;
    wire N__45306;
    wire N__45301;
    wire N__45298;
    wire N__45295;
    wire N__45292;
    wire N__45289;
    wire N__45286;
    wire N__45283;
    wire N__45280;
    wire N__45279;
    wire N__45276;
    wire N__45273;
    wire N__45270;
    wire N__45267;
    wire N__45266;
    wire N__45261;
    wire N__45258;
    wire N__45255;
    wire N__45250;
    wire N__45247;
    wire N__45244;
    wire N__45241;
    wire N__45238;
    wire N__45235;
    wire N__45232;
    wire N__45229;
    wire N__45226;
    wire N__45225;
    wire N__45222;
    wire N__45219;
    wire N__45216;
    wire N__45215;
    wire N__45212;
    wire N__45209;
    wire N__45206;
    wire N__45203;
    wire N__45196;
    wire N__45193;
    wire N__45190;
    wire N__45187;
    wire N__45184;
    wire N__45181;
    wire N__45178;
    wire N__45175;
    wire N__45174;
    wire N__45171;
    wire N__45168;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45156;
    wire N__45155;
    wire N__45152;
    wire N__45149;
    wire N__45146;
    wire N__45139;
    wire N__45136;
    wire N__45133;
    wire N__45130;
    wire N__45127;
    wire N__45124;
    wire N__45121;
    wire N__45118;
    wire N__45115;
    wire N__45112;
    wire N__45109;
    wire N__45106;
    wire N__45103;
    wire N__45100;
    wire N__45097;
    wire N__45094;
    wire N__45091;
    wire N__45088;
    wire N__45085;
    wire N__45082;
    wire N__45081;
    wire N__45078;
    wire N__45077;
    wire N__45074;
    wire N__45073;
    wire N__45070;
    wire N__45069;
    wire N__45066;
    wire N__45065;
    wire N__45064;
    wire N__45061;
    wire N__45058;
    wire N__45055;
    wire N__45052;
    wire N__45049;
    wire N__45044;
    wire N__45039;
    wire N__45034;
    wire N__45027;
    wire N__45022;
    wire N__45019;
    wire N__45018;
    wire N__45015;
    wire N__45012;
    wire N__45007;
    wire N__45004;
    wire N__45001;
    wire N__44998;
    wire N__44995;
    wire N__44992;
    wire N__44989;
    wire N__44986;
    wire N__44983;
    wire N__44980;
    wire N__44977;
    wire N__44974;
    wire N__44971;
    wire N__44968;
    wire N__44965;
    wire N__44962;
    wire N__44959;
    wire N__44956;
    wire N__44953;
    wire N__44950;
    wire N__44947;
    wire N__44944;
    wire N__44941;
    wire N__44938;
    wire N__44935;
    wire N__44932;
    wire N__44929;
    wire N__44926;
    wire N__44925;
    wire N__44922;
    wire N__44921;
    wire N__44918;
    wire N__44915;
    wire N__44912;
    wire N__44905;
    wire N__44902;
    wire N__44899;
    wire N__44898;
    wire N__44895;
    wire N__44892;
    wire N__44889;
    wire N__44886;
    wire N__44881;
    wire N__44880;
    wire N__44877;
    wire N__44874;
    wire N__44871;
    wire N__44866;
    wire N__44863;
    wire N__44860;
    wire N__44857;
    wire N__44854;
    wire N__44851;
    wire N__44848;
    wire N__44845;
    wire N__44842;
    wire N__44839;
    wire N__44836;
    wire N__44833;
    wire N__44830;
    wire N__44827;
    wire N__44824;
    wire N__44821;
    wire N__44818;
    wire N__44817;
    wire N__44814;
    wire N__44811;
    wire N__44806;
    wire N__44803;
    wire N__44802;
    wire N__44799;
    wire N__44794;
    wire N__44791;
    wire N__44790;
    wire N__44787;
    wire N__44784;
    wire N__44781;
    wire N__44778;
    wire N__44773;
    wire N__44770;
    wire N__44767;
    wire N__44764;
    wire N__44761;
    wire N__44758;
    wire N__44755;
    wire N__44752;
    wire N__44749;
    wire N__44746;
    wire N__44743;
    wire N__44740;
    wire N__44737;
    wire N__44734;
    wire N__44731;
    wire N__44728;
    wire N__44725;
    wire N__44724;
    wire N__44723;
    wire N__44720;
    wire N__44715;
    wire N__44710;
    wire N__44707;
    wire N__44704;
    wire N__44703;
    wire N__44702;
    wire N__44699;
    wire N__44698;
    wire N__44697;
    wire N__44696;
    wire N__44695;
    wire N__44692;
    wire N__44689;
    wire N__44686;
    wire N__44683;
    wire N__44678;
    wire N__44673;
    wire N__44662;
    wire N__44661;
    wire N__44660;
    wire N__44659;
    wire N__44656;
    wire N__44655;
    wire N__44654;
    wire N__44653;
    wire N__44650;
    wire N__44647;
    wire N__44644;
    wire N__44637;
    wire N__44634;
    wire N__44623;
    wire N__44620;
    wire N__44619;
    wire N__44618;
    wire N__44615;
    wire N__44612;
    wire N__44609;
    wire N__44608;
    wire N__44607;
    wire N__44606;
    wire N__44603;
    wire N__44600;
    wire N__44597;
    wire N__44592;
    wire N__44591;
    wire N__44588;
    wire N__44583;
    wire N__44578;
    wire N__44575;
    wire N__44572;
    wire N__44567;
    wire N__44560;
    wire N__44559;
    wire N__44556;
    wire N__44553;
    wire N__44550;
    wire N__44545;
    wire N__44542;
    wire N__44541;
    wire N__44538;
    wire N__44535;
    wire N__44534;
    wire N__44529;
    wire N__44526;
    wire N__44523;
    wire N__44518;
    wire N__44515;
    wire N__44512;
    wire N__44509;
    wire N__44506;
    wire N__44505;
    wire N__44502;
    wire N__44499;
    wire N__44496;
    wire N__44493;
    wire N__44492;
    wire N__44491;
    wire N__44488;
    wire N__44485;
    wire N__44480;
    wire N__44473;
    wire N__44470;
    wire N__44469;
    wire N__44468;
    wire N__44465;
    wire N__44462;
    wire N__44459;
    wire N__44454;
    wire N__44449;
    wire N__44448;
    wire N__44445;
    wire N__44444;
    wire N__44443;
    wire N__44440;
    wire N__44437;
    wire N__44432;
    wire N__44429;
    wire N__44424;
    wire N__44419;
    wire N__44416;
    wire N__44415;
    wire N__44412;
    wire N__44409;
    wire N__44406;
    wire N__44401;
    wire N__44400;
    wire N__44399;
    wire N__44398;
    wire N__44395;
    wire N__44388;
    wire N__44383;
    wire N__44380;
    wire N__44379;
    wire N__44378;
    wire N__44375;
    wire N__44372;
    wire N__44369;
    wire N__44362;
    wire N__44361;
    wire N__44356;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44344;
    wire N__44343;
    wire N__44340;
    wire N__44337;
    wire N__44336;
    wire N__44333;
    wire N__44330;
    wire N__44327;
    wire N__44320;
    wire N__44317;
    wire N__44314;
    wire N__44311;
    wire N__44310;
    wire N__44309;
    wire N__44308;
    wire N__44305;
    wire N__44302;
    wire N__44299;
    wire N__44298;
    wire N__44297;
    wire N__44294;
    wire N__44293;
    wire N__44292;
    wire N__44287;
    wire N__44282;
    wire N__44279;
    wire N__44272;
    wire N__44263;
    wire N__44260;
    wire N__44257;
    wire N__44256;
    wire N__44255;
    wire N__44252;
    wire N__44251;
    wire N__44248;
    wire N__44245;
    wire N__44242;
    wire N__44239;
    wire N__44236;
    wire N__44227;
    wire N__44224;
    wire N__44221;
    wire N__44220;
    wire N__44217;
    wire N__44214;
    wire N__44211;
    wire N__44206;
    wire N__44203;
    wire N__44200;
    wire N__44197;
    wire N__44194;
    wire N__44191;
    wire N__44188;
    wire N__44185;
    wire N__44182;
    wire N__44181;
    wire N__44178;
    wire N__44175;
    wire N__44172;
    wire N__44167;
    wire N__44166;
    wire N__44165;
    wire N__44162;
    wire N__44159;
    wire N__44156;
    wire N__44153;
    wire N__44150;
    wire N__44147;
    wire N__44146;
    wire N__44145;
    wire N__44142;
    wire N__44137;
    wire N__44136;
    wire N__44135;
    wire N__44132;
    wire N__44129;
    wire N__44126;
    wire N__44123;
    wire N__44120;
    wire N__44115;
    wire N__44104;
    wire N__44103;
    wire N__44100;
    wire N__44099;
    wire N__44096;
    wire N__44093;
    wire N__44090;
    wire N__44087;
    wire N__44080;
    wire N__44079;
    wire N__44078;
    wire N__44073;
    wire N__44070;
    wire N__44065;
    wire N__44064;
    wire N__44061;
    wire N__44058;
    wire N__44053;
    wire N__44050;
    wire N__44049;
    wire N__44048;
    wire N__44045;
    wire N__44042;
    wire N__44039;
    wire N__44038;
    wire N__44035;
    wire N__44032;
    wire N__44029;
    wire N__44026;
    wire N__44021;
    wire N__44014;
    wire N__44013;
    wire N__44012;
    wire N__44009;
    wire N__44006;
    wire N__44003;
    wire N__44000;
    wire N__43993;
    wire N__43990;
    wire N__43987;
    wire N__43984;
    wire N__43981;
    wire N__43978;
    wire N__43975;
    wire N__43972;
    wire N__43971;
    wire N__43970;
    wire N__43967;
    wire N__43962;
    wire N__43959;
    wire N__43956;
    wire N__43951;
    wire N__43948;
    wire N__43945;
    wire N__43942;
    wire N__43939;
    wire N__43936;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43921;
    wire N__43920;
    wire N__43919;
    wire N__43918;
    wire N__43915;
    wire N__43910;
    wire N__43907;
    wire N__43904;
    wire N__43901;
    wire N__43900;
    wire N__43899;
    wire N__43892;
    wire N__43889;
    wire N__43886;
    wire N__43879;
    wire N__43878;
    wire N__43875;
    wire N__43872;
    wire N__43871;
    wire N__43870;
    wire N__43869;
    wire N__43868;
    wire N__43865;
    wire N__43862;
    wire N__43859;
    wire N__43856;
    wire N__43851;
    wire N__43848;
    wire N__43837;
    wire N__43834;
    wire N__43833;
    wire N__43830;
    wire N__43827;
    wire N__43822;
    wire N__43819;
    wire N__43818;
    wire N__43817;
    wire N__43814;
    wire N__43811;
    wire N__43810;
    wire N__43809;
    wire N__43808;
    wire N__43807;
    wire N__43806;
    wire N__43803;
    wire N__43800;
    wire N__43797;
    wire N__43794;
    wire N__43791;
    wire N__43784;
    wire N__43771;
    wire N__43770;
    wire N__43767;
    wire N__43764;
    wire N__43759;
    wire N__43756;
    wire N__43753;
    wire N__43752;
    wire N__43751;
    wire N__43748;
    wire N__43745;
    wire N__43742;
    wire N__43735;
    wire N__43732;
    wire N__43729;
    wire N__43728;
    wire N__43725;
    wire N__43724;
    wire N__43723;
    wire N__43720;
    wire N__43715;
    wire N__43712;
    wire N__43705;
    wire N__43702;
    wire N__43699;
    wire N__43696;
    wire N__43693;
    wire N__43690;
    wire N__43687;
    wire N__43684;
    wire N__43681;
    wire N__43678;
    wire N__43675;
    wire N__43672;
    wire N__43669;
    wire N__43666;
    wire N__43663;
    wire N__43660;
    wire N__43657;
    wire N__43654;
    wire N__43651;
    wire N__43648;
    wire N__43645;
    wire N__43644;
    wire N__43639;
    wire N__43636;
    wire N__43633;
    wire N__43630;
    wire N__43629;
    wire N__43626;
    wire N__43623;
    wire N__43620;
    wire N__43617;
    wire N__43612;
    wire N__43609;
    wire N__43606;
    wire N__43605;
    wire N__43604;
    wire N__43599;
    wire N__43596;
    wire N__43591;
    wire N__43588;
    wire N__43585;
    wire N__43582;
    wire N__43579;
    wire N__43576;
    wire N__43573;
    wire N__43572;
    wire N__43571;
    wire N__43564;
    wire N__43561;
    wire N__43558;
    wire N__43557;
    wire N__43552;
    wire N__43549;
    wire N__43546;
    wire N__43543;
    wire N__43540;
    wire N__43539;
    wire N__43536;
    wire N__43533;
    wire N__43532;
    wire N__43531;
    wire N__43526;
    wire N__43523;
    wire N__43520;
    wire N__43517;
    wire N__43510;
    wire N__43507;
    wire N__43504;
    wire N__43503;
    wire N__43502;
    wire N__43499;
    wire N__43496;
    wire N__43493;
    wire N__43488;
    wire N__43487;
    wire N__43484;
    wire N__43481;
    wire N__43478;
    wire N__43475;
    wire N__43472;
    wire N__43465;
    wire N__43462;
    wire N__43459;
    wire N__43456;
    wire N__43455;
    wire N__43452;
    wire N__43451;
    wire N__43448;
    wire N__43445;
    wire N__43444;
    wire N__43441;
    wire N__43436;
    wire N__43433;
    wire N__43430;
    wire N__43427;
    wire N__43420;
    wire N__43417;
    wire N__43414;
    wire N__43411;
    wire N__43410;
    wire N__43407;
    wire N__43404;
    wire N__43401;
    wire N__43398;
    wire N__43395;
    wire N__43394;
    wire N__43393;
    wire N__43388;
    wire N__43385;
    wire N__43382;
    wire N__43379;
    wire N__43372;
    wire N__43369;
    wire N__43366;
    wire N__43363;
    wire N__43362;
    wire N__43361;
    wire N__43358;
    wire N__43353;
    wire N__43350;
    wire N__43345;
    wire N__43344;
    wire N__43343;
    wire N__43342;
    wire N__43341;
    wire N__43340;
    wire N__43333;
    wire N__43330;
    wire N__43325;
    wire N__43322;
    wire N__43319;
    wire N__43314;
    wire N__43311;
    wire N__43306;
    wire N__43303;
    wire N__43300;
    wire N__43297;
    wire N__43294;
    wire N__43291;
    wire N__43290;
    wire N__43287;
    wire N__43284;
    wire N__43279;
    wire N__43276;
    wire N__43273;
    wire N__43270;
    wire N__43269;
    wire N__43268;
    wire N__43267;
    wire N__43266;
    wire N__43265;
    wire N__43264;
    wire N__43263;
    wire N__43262;
    wire N__43261;
    wire N__43260;
    wire N__43259;
    wire N__43258;
    wire N__43251;
    wire N__43246;
    wire N__43245;
    wire N__43244;
    wire N__43243;
    wire N__43240;
    wire N__43239;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43227;
    wire N__43220;
    wire N__43219;
    wire N__43218;
    wire N__43217;
    wire N__43216;
    wire N__43215;
    wire N__43210;
    wire N__43199;
    wire N__43194;
    wire N__43193;
    wire N__43192;
    wire N__43185;
    wire N__43182;
    wire N__43179;
    wire N__43176;
    wire N__43175;
    wire N__43172;
    wire N__43171;
    wire N__43170;
    wire N__43169;
    wire N__43166;
    wire N__43161;
    wire N__43158;
    wire N__43157;
    wire N__43156;
    wire N__43155;
    wire N__43154;
    wire N__43151;
    wire N__43148;
    wire N__43139;
    wire N__43136;
    wire N__43133;
    wire N__43130;
    wire N__43125;
    wire N__43120;
    wire N__43117;
    wire N__43112;
    wire N__43111;
    wire N__43110;
    wire N__43109;
    wire N__43106;
    wire N__43103;
    wire N__43096;
    wire N__43091;
    wire N__43080;
    wire N__43079;
    wire N__43072;
    wire N__43067;
    wire N__43064;
    wire N__43059;
    wire N__43056;
    wire N__43045;
    wire N__43044;
    wire N__43043;
    wire N__43038;
    wire N__43035;
    wire N__43032;
    wire N__43031;
    wire N__43028;
    wire N__43025;
    wire N__43022;
    wire N__43019;
    wire N__43016;
    wire N__43009;
    wire N__43008;
    wire N__43007;
    wire N__43004;
    wire N__43001;
    wire N__42998;
    wire N__42995;
    wire N__42990;
    wire N__42985;
    wire N__42982;
    wire N__42979;
    wire N__42978;
    wire N__42975;
    wire N__42972;
    wire N__42971;
    wire N__42966;
    wire N__42963;
    wire N__42958;
    wire N__42955;
    wire N__42954;
    wire N__42951;
    wire N__42948;
    wire N__42943;
    wire N__42940;
    wire N__42937;
    wire N__42936;
    wire N__42935;
    wire N__42932;
    wire N__42929;
    wire N__42928;
    wire N__42925;
    wire N__42922;
    wire N__42919;
    wire N__42916;
    wire N__42913;
    wire N__42910;
    wire N__42907;
    wire N__42898;
    wire N__42895;
    wire N__42892;
    wire N__42889;
    wire N__42886;
    wire N__42885;
    wire N__42884;
    wire N__42881;
    wire N__42880;
    wire N__42877;
    wire N__42874;
    wire N__42871;
    wire N__42870;
    wire N__42867;
    wire N__42864;
    wire N__42859;
    wire N__42856;
    wire N__42853;
    wire N__42850;
    wire N__42847;
    wire N__42844;
    wire N__42835;
    wire N__42834;
    wire N__42833;
    wire N__42830;
    wire N__42827;
    wire N__42826;
    wire N__42825;
    wire N__42822;
    wire N__42819;
    wire N__42816;
    wire N__42813;
    wire N__42810;
    wire N__42799;
    wire N__42798;
    wire N__42797;
    wire N__42796;
    wire N__42795;
    wire N__42794;
    wire N__42793;
    wire N__42792;
    wire N__42791;
    wire N__42790;
    wire N__42789;
    wire N__42788;
    wire N__42787;
    wire N__42786;
    wire N__42785;
    wire N__42782;
    wire N__42779;
    wire N__42770;
    wire N__42769;
    wire N__42768;
    wire N__42767;
    wire N__42766;
    wire N__42755;
    wire N__42752;
    wire N__42745;
    wire N__42744;
    wire N__42743;
    wire N__42740;
    wire N__42737;
    wire N__42734;
    wire N__42729;
    wire N__42724;
    wire N__42721;
    wire N__42716;
    wire N__42711;
    wire N__42710;
    wire N__42709;
    wire N__42708;
    wire N__42707;
    wire N__42706;
    wire N__42705;
    wire N__42704;
    wire N__42703;
    wire N__42700;
    wire N__42693;
    wire N__42690;
    wire N__42687;
    wire N__42682;
    wire N__42675;
    wire N__42664;
    wire N__42649;
    wire N__42646;
    wire N__42643;
    wire N__42640;
    wire N__42639;
    wire N__42638;
    wire N__42635;
    wire N__42632;
    wire N__42629;
    wire N__42624;
    wire N__42621;
    wire N__42616;
    wire N__42615;
    wire N__42612;
    wire N__42611;
    wire N__42610;
    wire N__42605;
    wire N__42602;
    wire N__42599;
    wire N__42594;
    wire N__42589;
    wire N__42586;
    wire N__42585;
    wire N__42584;
    wire N__42581;
    wire N__42578;
    wire N__42575;
    wire N__42568;
    wire N__42567;
    wire N__42564;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42550;
    wire N__42547;
    wire N__42546;
    wire N__42545;
    wire N__42542;
    wire N__42539;
    wire N__42538;
    wire N__42535;
    wire N__42532;
    wire N__42529;
    wire N__42524;
    wire N__42521;
    wire N__42518;
    wire N__42515;
    wire N__42508;
    wire N__42507;
    wire N__42506;
    wire N__42503;
    wire N__42502;
    wire N__42499;
    wire N__42498;
    wire N__42495;
    wire N__42494;
    wire N__42493;
    wire N__42490;
    wire N__42487;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42473;
    wire N__42470;
    wire N__42463;
    wire N__42460;
    wire N__42453;
    wire N__42448;
    wire N__42445;
    wire N__42442;
    wire N__42439;
    wire N__42436;
    wire N__42433;
    wire N__42430;
    wire N__42429;
    wire N__42426;
    wire N__42423;
    wire N__42420;
    wire N__42417;
    wire N__42412;
    wire N__42409;
    wire N__42406;
    wire N__42403;
    wire N__42400;
    wire N__42397;
    wire N__42396;
    wire N__42395;
    wire N__42392;
    wire N__42389;
    wire N__42386;
    wire N__42385;
    wire N__42382;
    wire N__42379;
    wire N__42376;
    wire N__42375;
    wire N__42372;
    wire N__42367;
    wire N__42364;
    wire N__42361;
    wire N__42352;
    wire N__42351;
    wire N__42348;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42338;
    wire N__42337;
    wire N__42336;
    wire N__42333;
    wire N__42330;
    wire N__42325;
    wire N__42322;
    wire N__42315;
    wire N__42310;
    wire N__42307;
    wire N__42306;
    wire N__42303;
    wire N__42300;
    wire N__42297;
    wire N__42294;
    wire N__42293;
    wire N__42290;
    wire N__42287;
    wire N__42286;
    wire N__42283;
    wire N__42280;
    wire N__42277;
    wire N__42274;
    wire N__42265;
    wire N__42262;
    wire N__42259;
    wire N__42256;
    wire N__42253;
    wire N__42252;
    wire N__42251;
    wire N__42250;
    wire N__42249;
    wire N__42248;
    wire N__42245;
    wire N__42242;
    wire N__42241;
    wire N__42240;
    wire N__42239;
    wire N__42238;
    wire N__42237;
    wire N__42236;
    wire N__42235;
    wire N__42234;
    wire N__42233;
    wire N__42232;
    wire N__42231;
    wire N__42224;
    wire N__42223;
    wire N__42222;
    wire N__42221;
    wire N__42210;
    wire N__42209;
    wire N__42208;
    wire N__42205;
    wire N__42204;
    wire N__42203;
    wire N__42202;
    wire N__42199;
    wire N__42190;
    wire N__42187;
    wire N__42184;
    wire N__42181;
    wire N__42180;
    wire N__42177;
    wire N__42172;
    wire N__42169;
    wire N__42168;
    wire N__42167;
    wire N__42164;
    wire N__42155;
    wire N__42152;
    wire N__42151;
    wire N__42150;
    wire N__42147;
    wire N__42138;
    wire N__42133;
    wire N__42128;
    wire N__42123;
    wire N__42120;
    wire N__42115;
    wire N__42108;
    wire N__42107;
    wire N__42106;
    wire N__42103;
    wire N__42100;
    wire N__42097;
    wire N__42090;
    wire N__42085;
    wire N__42082;
    wire N__42079;
    wire N__42076;
    wire N__42071;
    wire N__42062;
    wire N__42059;
    wire N__42056;
    wire N__42053;
    wire N__42046;
    wire N__42045;
    wire N__42042;
    wire N__42041;
    wire N__42038;
    wire N__42035;
    wire N__42034;
    wire N__42031;
    wire N__42030;
    wire N__42027;
    wire N__42024;
    wire N__42021;
    wire N__42018;
    wire N__42015;
    wire N__42010;
    wire N__42007;
    wire N__41998;
    wire N__41995;
    wire N__41994;
    wire N__41993;
    wire N__41992;
    wire N__41989;
    wire N__41986;
    wire N__41981;
    wire N__41976;
    wire N__41971;
    wire N__41968;
    wire N__41967;
    wire N__41964;
    wire N__41961;
    wire N__41960;
    wire N__41957;
    wire N__41954;
    wire N__41951;
    wire N__41950;
    wire N__41947;
    wire N__41944;
    wire N__41941;
    wire N__41938;
    wire N__41935;
    wire N__41930;
    wire N__41923;
    wire N__41920;
    wire N__41917;
    wire N__41914;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41904;
    wire N__41899;
    wire N__41896;
    wire N__41893;
    wire N__41890;
    wire N__41889;
    wire N__41888;
    wire N__41885;
    wire N__41880;
    wire N__41877;
    wire N__41872;
    wire N__41871;
    wire N__41870;
    wire N__41869;
    wire N__41866;
    wire N__41863;
    wire N__41862;
    wire N__41859;
    wire N__41856;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41844;
    wire N__41843;
    wire N__41840;
    wire N__41833;
    wire N__41830;
    wire N__41827;
    wire N__41822;
    wire N__41815;
    wire N__41812;
    wire N__41811;
    wire N__41810;
    wire N__41807;
    wire N__41804;
    wire N__41801;
    wire N__41800;
    wire N__41799;
    wire N__41796;
    wire N__41791;
    wire N__41788;
    wire N__41785;
    wire N__41784;
    wire N__41781;
    wire N__41774;
    wire N__41771;
    wire N__41768;
    wire N__41765;
    wire N__41758;
    wire N__41755;
    wire N__41754;
    wire N__41751;
    wire N__41750;
    wire N__41747;
    wire N__41746;
    wire N__41745;
    wire N__41744;
    wire N__41741;
    wire N__41738;
    wire N__41735;
    wire N__41728;
    wire N__41723;
    wire N__41722;
    wire N__41719;
    wire N__41714;
    wire N__41711;
    wire N__41704;
    wire N__41701;
    wire N__41700;
    wire N__41697;
    wire N__41696;
    wire N__41693;
    wire N__41690;
    wire N__41687;
    wire N__41684;
    wire N__41683;
    wire N__41682;
    wire N__41679;
    wire N__41674;
    wire N__41673;
    wire N__41670;
    wire N__41667;
    wire N__41662;
    wire N__41657;
    wire N__41650;
    wire N__41649;
    wire N__41648;
    wire N__41647;
    wire N__41646;
    wire N__41645;
    wire N__41642;
    wire N__41635;
    wire N__41632;
    wire N__41629;
    wire N__41628;
    wire N__41623;
    wire N__41620;
    wire N__41615;
    wire N__41612;
    wire N__41605;
    wire N__41602;
    wire N__41601;
    wire N__41598;
    wire N__41595;
    wire N__41592;
    wire N__41587;
    wire N__41584;
    wire N__41581;
    wire N__41578;
    wire N__41577;
    wire N__41574;
    wire N__41571;
    wire N__41568;
    wire N__41563;
    wire N__41560;
    wire N__41557;
    wire N__41554;
    wire N__41551;
    wire N__41548;
    wire N__41547;
    wire N__41546;
    wire N__41541;
    wire N__41538;
    wire N__41535;
    wire N__41534;
    wire N__41531;
    wire N__41528;
    wire N__41525;
    wire N__41522;
    wire N__41519;
    wire N__41512;
    wire N__41509;
    wire N__41506;
    wire N__41503;
    wire N__41500;
    wire N__41497;
    wire N__41496;
    wire N__41493;
    wire N__41492;
    wire N__41491;
    wire N__41490;
    wire N__41487;
    wire N__41486;
    wire N__41485;
    wire N__41484;
    wire N__41479;
    wire N__41476;
    wire N__41471;
    wire N__41468;
    wire N__41467;
    wire N__41462;
    wire N__41459;
    wire N__41458;
    wire N__41457;
    wire N__41456;
    wire N__41455;
    wire N__41454;
    wire N__41451;
    wire N__41446;
    wire N__41445;
    wire N__41444;
    wire N__41443;
    wire N__41440;
    wire N__41437;
    wire N__41434;
    wire N__41429;
    wire N__41422;
    wire N__41419;
    wire N__41416;
    wire N__41413;
    wire N__41406;
    wire N__41399;
    wire N__41386;
    wire N__41383;
    wire N__41382;
    wire N__41379;
    wire N__41378;
    wire N__41377;
    wire N__41376;
    wire N__41375;
    wire N__41374;
    wire N__41373;
    wire N__41370;
    wire N__41367;
    wire N__41362;
    wire N__41353;
    wire N__41344;
    wire N__41343;
    wire N__41342;
    wire N__41339;
    wire N__41334;
    wire N__41331;
    wire N__41328;
    wire N__41327;
    wire N__41324;
    wire N__41321;
    wire N__41318;
    wire N__41315;
    wire N__41312;
    wire N__41305;
    wire N__41302;
    wire N__41299;
    wire N__41296;
    wire N__41293;
    wire N__41290;
    wire N__41287;
    wire N__41284;
    wire N__41281;
    wire N__41278;
    wire N__41277;
    wire N__41274;
    wire N__41271;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41257;
    wire N__41254;
    wire N__41253;
    wire N__41250;
    wire N__41247;
    wire N__41244;
    wire N__41239;
    wire N__41236;
    wire N__41233;
    wire N__41230;
    wire N__41227;
    wire N__41224;
    wire N__41221;
    wire N__41218;
    wire N__41215;
    wire N__41212;
    wire N__41209;
    wire N__41208;
    wire N__41205;
    wire N__41202;
    wire N__41197;
    wire N__41194;
    wire N__41191;
    wire N__41188;
    wire N__41185;
    wire N__41182;
    wire N__41179;
    wire N__41178;
    wire N__41173;
    wire N__41170;
    wire N__41167;
    wire N__41164;
    wire N__41161;
    wire N__41158;
    wire N__41155;
    wire N__41152;
    wire N__41151;
    wire N__41148;
    wire N__41147;
    wire N__41146;
    wire N__41143;
    wire N__41140;
    wire N__41135;
    wire N__41132;
    wire N__41129;
    wire N__41122;
    wire N__41119;
    wire N__41116;
    wire N__41113;
    wire N__41110;
    wire N__41107;
    wire N__41104;
    wire N__41101;
    wire N__41100;
    wire N__41099;
    wire N__41096;
    wire N__41093;
    wire N__41090;
    wire N__41087;
    wire N__41084;
    wire N__41083;
    wire N__41076;
    wire N__41073;
    wire N__41070;
    wire N__41065;
    wire N__41062;
    wire N__41059;
    wire N__41056;
    wire N__41053;
    wire N__41052;
    wire N__41049;
    wire N__41048;
    wire N__41045;
    wire N__41042;
    wire N__41041;
    wire N__41038;
    wire N__41035;
    wire N__41032;
    wire N__41029;
    wire N__41020;
    wire N__41017;
    wire N__41014;
    wire N__41011;
    wire N__41008;
    wire N__41007;
    wire N__41004;
    wire N__41003;
    wire N__41000;
    wire N__40997;
    wire N__40996;
    wire N__40993;
    wire N__40990;
    wire N__40987;
    wire N__40984;
    wire N__40981;
    wire N__40978;
    wire N__40975;
    wire N__40966;
    wire N__40963;
    wire N__40960;
    wire N__40957;
    wire N__40954;
    wire N__40953;
    wire N__40952;
    wire N__40951;
    wire N__40950;
    wire N__40947;
    wire N__40946;
    wire N__40945;
    wire N__40944;
    wire N__40941;
    wire N__40938;
    wire N__40935;
    wire N__40934;
    wire N__40931;
    wire N__40928;
    wire N__40927;
    wire N__40924;
    wire N__40921;
    wire N__40918;
    wire N__40915;
    wire N__40912;
    wire N__40909;
    wire N__40906;
    wire N__40903;
    wire N__40900;
    wire N__40897;
    wire N__40894;
    wire N__40891;
    wire N__40886;
    wire N__40883;
    wire N__40880;
    wire N__40877;
    wire N__40874;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40858;
    wire N__40855;
    wire N__40852;
    wire N__40849;
    wire N__40846;
    wire N__40843;
    wire N__40840;
    wire N__40837;
    wire N__40834;
    wire N__40829;
    wire N__40826;
    wire N__40821;
    wire N__40818;
    wire N__40807;
    wire N__40804;
    wire N__40801;
    wire N__40798;
    wire N__40795;
    wire N__40792;
    wire N__40789;
    wire N__40786;
    wire N__40783;
    wire N__40780;
    wire N__40777;
    wire N__40776;
    wire N__40775;
    wire N__40770;
    wire N__40767;
    wire N__40764;
    wire N__40761;
    wire N__40758;
    wire N__40755;
    wire N__40750;
    wire N__40749;
    wire N__40746;
    wire N__40745;
    wire N__40744;
    wire N__40741;
    wire N__40738;
    wire N__40735;
    wire N__40734;
    wire N__40731;
    wire N__40728;
    wire N__40725;
    wire N__40722;
    wire N__40717;
    wire N__40714;
    wire N__40705;
    wire N__40702;
    wire N__40701;
    wire N__40698;
    wire N__40695;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40678;
    wire N__40675;
    wire N__40672;
    wire N__40671;
    wire N__40670;
    wire N__40667;
    wire N__40662;
    wire N__40657;
    wire N__40654;
    wire N__40653;
    wire N__40652;
    wire N__40649;
    wire N__40644;
    wire N__40641;
    wire N__40638;
    wire N__40633;
    wire N__40630;
    wire N__40629;
    wire N__40628;
    wire N__40625;
    wire N__40624;
    wire N__40623;
    wire N__40618;
    wire N__40615;
    wire N__40610;
    wire N__40607;
    wire N__40600;
    wire N__40599;
    wire N__40598;
    wire N__40597;
    wire N__40596;
    wire N__40595;
    wire N__40592;
    wire N__40589;
    wire N__40586;
    wire N__40585;
    wire N__40582;
    wire N__40577;
    wire N__40576;
    wire N__40575;
    wire N__40572;
    wire N__40569;
    wire N__40562;
    wire N__40559;
    wire N__40556;
    wire N__40553;
    wire N__40540;
    wire N__40539;
    wire N__40536;
    wire N__40535;
    wire N__40528;
    wire N__40527;
    wire N__40524;
    wire N__40521;
    wire N__40516;
    wire N__40513;
    wire N__40512;
    wire N__40509;
    wire N__40506;
    wire N__40505;
    wire N__40502;
    wire N__40497;
    wire N__40492;
    wire N__40489;
    wire N__40486;
    wire N__40483;
    wire N__40480;
    wire N__40477;
    wire N__40474;
    wire N__40471;
    wire N__40468;
    wire N__40465;
    wire N__40462;
    wire N__40459;
    wire N__40456;
    wire N__40455;
    wire N__40454;
    wire N__40453;
    wire N__40448;
    wire N__40447;
    wire N__40446;
    wire N__40445;
    wire N__40440;
    wire N__40437;
    wire N__40430;
    wire N__40423;
    wire N__40420;
    wire N__40419;
    wire N__40418;
    wire N__40415;
    wire N__40412;
    wire N__40409;
    wire N__40402;
    wire N__40401;
    wire N__40396;
    wire N__40393;
    wire N__40390;
    wire N__40387;
    wire N__40384;
    wire N__40381;
    wire N__40378;
    wire N__40375;
    wire N__40372;
    wire N__40369;
    wire N__40368;
    wire N__40367;
    wire N__40366;
    wire N__40363;
    wire N__40360;
    wire N__40359;
    wire N__40356;
    wire N__40355;
    wire N__40352;
    wire N__40349;
    wire N__40346;
    wire N__40343;
    wire N__40340;
    wire N__40337;
    wire N__40334;
    wire N__40331;
    wire N__40328;
    wire N__40325;
    wire N__40312;
    wire N__40309;
    wire N__40306;
    wire N__40305;
    wire N__40304;
    wire N__40301;
    wire N__40298;
    wire N__40295;
    wire N__40294;
    wire N__40291;
    wire N__40288;
    wire N__40285;
    wire N__40284;
    wire N__40281;
    wire N__40276;
    wire N__40273;
    wire N__40268;
    wire N__40261;
    wire N__40258;
    wire N__40257;
    wire N__40254;
    wire N__40251;
    wire N__40246;
    wire N__40243;
    wire N__40242;
    wire N__40241;
    wire N__40238;
    wire N__40233;
    wire N__40232;
    wire N__40229;
    wire N__40226;
    wire N__40223;
    wire N__40218;
    wire N__40213;
    wire N__40210;
    wire N__40209;
    wire N__40208;
    wire N__40205;
    wire N__40202;
    wire N__40199;
    wire N__40198;
    wire N__40195;
    wire N__40192;
    wire N__40189;
    wire N__40186;
    wire N__40179;
    wire N__40174;
    wire N__40171;
    wire N__40170;
    wire N__40169;
    wire N__40166;
    wire N__40163;
    wire N__40160;
    wire N__40159;
    wire N__40158;
    wire N__40157;
    wire N__40154;
    wire N__40151;
    wire N__40150;
    wire N__40149;
    wire N__40146;
    wire N__40143;
    wire N__40138;
    wire N__40133;
    wire N__40128;
    wire N__40125;
    wire N__40120;
    wire N__40115;
    wire N__40114;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40104;
    wire N__40099;
    wire N__40090;
    wire N__40087;
    wire N__40084;
    wire N__40081;
    wire N__40078;
    wire N__40075;
    wire N__40072;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40060;
    wire N__40059;
    wire N__40058;
    wire N__40057;
    wire N__40056;
    wire N__40053;
    wire N__40050;
    wire N__40047;
    wire N__40044;
    wire N__40041;
    wire N__40040;
    wire N__40039;
    wire N__40036;
    wire N__40033;
    wire N__40028;
    wire N__40025;
    wire N__40022;
    wire N__40019;
    wire N__40014;
    wire N__40011;
    wire N__40008;
    wire N__40005;
    wire N__39994;
    wire N__39991;
    wire N__39988;
    wire N__39985;
    wire N__39982;
    wire N__39979;
    wire N__39976;
    wire N__39975;
    wire N__39974;
    wire N__39971;
    wire N__39968;
    wire N__39967;
    wire N__39966;
    wire N__39963;
    wire N__39960;
    wire N__39957;
    wire N__39952;
    wire N__39943;
    wire N__39940;
    wire N__39937;
    wire N__39934;
    wire N__39933;
    wire N__39930;
    wire N__39927;
    wire N__39924;
    wire N__39919;
    wire N__39916;
    wire N__39913;
    wire N__39910;
    wire N__39907;
    wire N__39904;
    wire N__39903;
    wire N__39902;
    wire N__39899;
    wire N__39898;
    wire N__39895;
    wire N__39894;
    wire N__39893;
    wire N__39890;
    wire N__39889;
    wire N__39886;
    wire N__39883;
    wire N__39880;
    wire N__39875;
    wire N__39872;
    wire N__39869;
    wire N__39866;
    wire N__39863;
    wire N__39858;
    wire N__39847;
    wire N__39846;
    wire N__39841;
    wire N__39838;
    wire N__39837;
    wire N__39836;
    wire N__39835;
    wire N__39834;
    wire N__39833;
    wire N__39832;
    wire N__39829;
    wire N__39826;
    wire N__39823;
    wire N__39822;
    wire N__39819;
    wire N__39818;
    wire N__39817;
    wire N__39816;
    wire N__39815;
    wire N__39814;
    wire N__39811;
    wire N__39808;
    wire N__39807;
    wire N__39806;
    wire N__39805;
    wire N__39804;
    wire N__39801;
    wire N__39800;
    wire N__39799;
    wire N__39796;
    wire N__39791;
    wire N__39788;
    wire N__39785;
    wire N__39782;
    wire N__39781;
    wire N__39780;
    wire N__39779;
    wire N__39778;
    wire N__39777;
    wire N__39776;
    wire N__39775;
    wire N__39774;
    wire N__39773;
    wire N__39772;
    wire N__39771;
    wire N__39768;
    wire N__39763;
    wire N__39760;
    wire N__39759;
    wire N__39758;
    wire N__39757;
    wire N__39756;
    wire N__39751;
    wire N__39750;
    wire N__39749;
    wire N__39744;
    wire N__39741;
    wire N__39738;
    wire N__39735;
    wire N__39734;
    wire N__39733;
    wire N__39732;
    wire N__39727;
    wire N__39726;
    wire N__39721;
    wire N__39720;
    wire N__39715;
    wire N__39712;
    wire N__39709;
    wire N__39702;
    wire N__39701;
    wire N__39700;
    wire N__39697;
    wire N__39690;
    wire N__39687;
    wire N__39682;
    wire N__39679;
    wire N__39676;
    wire N__39673;
    wire N__39668;
    wire N__39663;
    wire N__39660;
    wire N__39655;
    wire N__39650;
    wire N__39647;
    wire N__39644;
    wire N__39639;
    wire N__39636;
    wire N__39633;
    wire N__39630;
    wire N__39627;
    wire N__39626;
    wire N__39623;
    wire N__39616;
    wire N__39613;
    wire N__39608;
    wire N__39603;
    wire N__39598;
    wire N__39591;
    wire N__39586;
    wire N__39583;
    wire N__39574;
    wire N__39569;
    wire N__39564;
    wire N__39561;
    wire N__39558;
    wire N__39555;
    wire N__39552;
    wire N__39541;
    wire N__39534;
    wire N__39525;
    wire N__39514;
    wire N__39511;
    wire N__39508;
    wire N__39505;
    wire N__39502;
    wire N__39499;
    wire N__39496;
    wire N__39495;
    wire N__39492;
    wire N__39489;
    wire N__39488;
    wire N__39487;
    wire N__39486;
    wire N__39481;
    wire N__39478;
    wire N__39477;
    wire N__39476;
    wire N__39475;
    wire N__39472;
    wire N__39469;
    wire N__39466;
    wire N__39463;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39447;
    wire N__39440;
    wire N__39433;
    wire N__39430;
    wire N__39427;
    wire N__39426;
    wire N__39423;
    wire N__39420;
    wire N__39417;
    wire N__39414;
    wire N__39411;
    wire N__39408;
    wire N__39403;
    wire N__39400;
    wire N__39397;
    wire N__39394;
    wire N__39393;
    wire N__39392;
    wire N__39391;
    wire N__39390;
    wire N__39387;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39372;
    wire N__39367;
    wire N__39364;
    wire N__39361;
    wire N__39360;
    wire N__39355;
    wire N__39350;
    wire N__39347;
    wire N__39340;
    wire N__39337;
    wire N__39334;
    wire N__39331;
    wire N__39328;
    wire N__39325;
    wire N__39324;
    wire N__39321;
    wire N__39320;
    wire N__39319;
    wire N__39318;
    wire N__39317;
    wire N__39314;
    wire N__39311;
    wire N__39308;
    wire N__39301;
    wire N__39292;
    wire N__39289;
    wire N__39288;
    wire N__39285;
    wire N__39282;
    wire N__39279;
    wire N__39274;
    wire N__39273;
    wire N__39270;
    wire N__39269;
    wire N__39268;
    wire N__39265;
    wire N__39264;
    wire N__39261;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39249;
    wire N__39248;
    wire N__39243;
    wire N__39236;
    wire N__39233;
    wire N__39230;
    wire N__39225;
    wire N__39220;
    wire N__39217;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39205;
    wire N__39202;
    wire N__39199;
    wire N__39196;
    wire N__39193;
    wire N__39190;
    wire N__39189;
    wire N__39186;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39166;
    wire N__39163;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39148;
    wire N__39145;
    wire N__39142;
    wire N__39139;
    wire N__39138;
    wire N__39135;
    wire N__39132;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39115;
    wire N__39114;
    wire N__39111;
    wire N__39108;
    wire N__39105;
    wire N__39102;
    wire N__39101;
    wire N__39098;
    wire N__39095;
    wire N__39092;
    wire N__39091;
    wire N__39090;
    wire N__39089;
    wire N__39086;
    wire N__39081;
    wire N__39078;
    wire N__39073;
    wire N__39064;
    wire N__39061;
    wire N__39060;
    wire N__39057;
    wire N__39056;
    wire N__39053;
    wire N__39050;
    wire N__39047;
    wire N__39040;
    wire N__39037;
    wire N__39036;
    wire N__39035;
    wire N__39032;
    wire N__39029;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39016;
    wire N__39015;
    wire N__39014;
    wire N__39009;
    wire N__39006;
    wire N__39001;
    wire N__38998;
    wire N__38989;
    wire N__38986;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38976;
    wire N__38971;
    wire N__38968;
    wire N__38967;
    wire N__38966;
    wire N__38965;
    wire N__38958;
    wire N__38955;
    wire N__38950;
    wire N__38947;
    wire N__38944;
    wire N__38941;
    wire N__38938;
    wire N__38935;
    wire N__38934;
    wire N__38931;
    wire N__38928;
    wire N__38925;
    wire N__38922;
    wire N__38917;
    wire N__38916;
    wire N__38915;
    wire N__38914;
    wire N__38911;
    wire N__38906;
    wire N__38905;
    wire N__38902;
    wire N__38897;
    wire N__38894;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38878;
    wire N__38875;
    wire N__38874;
    wire N__38871;
    wire N__38870;
    wire N__38869;
    wire N__38866;
    wire N__38863;
    wire N__38860;
    wire N__38859;
    wire N__38856;
    wire N__38851;
    wire N__38848;
    wire N__38847;
    wire N__38844;
    wire N__38841;
    wire N__38838;
    wire N__38835;
    wire N__38832;
    wire N__38821;
    wire N__38818;
    wire N__38815;
    wire N__38812;
    wire N__38809;
    wire N__38806;
    wire N__38803;
    wire N__38800;
    wire N__38797;
    wire N__38794;
    wire N__38791;
    wire N__38788;
    wire N__38785;
    wire N__38784;
    wire N__38783;
    wire N__38780;
    wire N__38777;
    wire N__38774;
    wire N__38773;
    wire N__38772;
    wire N__38771;
    wire N__38768;
    wire N__38765;
    wire N__38762;
    wire N__38757;
    wire N__38756;
    wire N__38753;
    wire N__38750;
    wire N__38745;
    wire N__38742;
    wire N__38739;
    wire N__38728;
    wire N__38725;
    wire N__38724;
    wire N__38723;
    wire N__38722;
    wire N__38719;
    wire N__38716;
    wire N__38715;
    wire N__38714;
    wire N__38711;
    wire N__38708;
    wire N__38705;
    wire N__38702;
    wire N__38697;
    wire N__38694;
    wire N__38687;
    wire N__38684;
    wire N__38677;
    wire N__38676;
    wire N__38671;
    wire N__38668;
    wire N__38667;
    wire N__38666;
    wire N__38663;
    wire N__38662;
    wire N__38659;
    wire N__38656;
    wire N__38653;
    wire N__38652;
    wire N__38649;
    wire N__38648;
    wire N__38645;
    wire N__38642;
    wire N__38639;
    wire N__38636;
    wire N__38633;
    wire N__38630;
    wire N__38627;
    wire N__38622;
    wire N__38611;
    wire N__38610;
    wire N__38607;
    wire N__38602;
    wire N__38599;
    wire N__38596;
    wire N__38593;
    wire N__38590;
    wire N__38587;
    wire N__38586;
    wire N__38583;
    wire N__38580;
    wire N__38579;
    wire N__38576;
    wire N__38573;
    wire N__38570;
    wire N__38563;
    wire N__38560;
    wire N__38557;
    wire N__38556;
    wire N__38553;
    wire N__38550;
    wire N__38545;
    wire N__38542;
    wire N__38539;
    wire N__38536;
    wire N__38533;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38521;
    wire N__38518;
    wire N__38515;
    wire N__38512;
    wire N__38509;
    wire N__38506;
    wire N__38505;
    wire N__38504;
    wire N__38503;
    wire N__38502;
    wire N__38501;
    wire N__38500;
    wire N__38499;
    wire N__38498;
    wire N__38497;
    wire N__38496;
    wire N__38493;
    wire N__38492;
    wire N__38491;
    wire N__38488;
    wire N__38485;
    wire N__38482;
    wire N__38473;
    wire N__38470;
    wire N__38467;
    wire N__38466;
    wire N__38465;
    wire N__38462;
    wire N__38461;
    wire N__38460;
    wire N__38459;
    wire N__38458;
    wire N__38457;
    wire N__38454;
    wire N__38449;
    wire N__38446;
    wire N__38443;
    wire N__38434;
    wire N__38431;
    wire N__38424;
    wire N__38419;
    wire N__38416;
    wire N__38413;
    wire N__38412;
    wire N__38411;
    wire N__38410;
    wire N__38405;
    wire N__38402;
    wire N__38397;
    wire N__38396;
    wire N__38395;
    wire N__38388;
    wire N__38383;
    wire N__38378;
    wire N__38377;
    wire N__38374;
    wire N__38367;
    wire N__38364;
    wire N__38361;
    wire N__38360;
    wire N__38359;
    wire N__38358;
    wire N__38357;
    wire N__38356;
    wire N__38353;
    wire N__38348;
    wire N__38343;
    wire N__38336;
    wire N__38327;
    wire N__38324;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38302;
    wire N__38299;
    wire N__38296;
    wire N__38295;
    wire N__38294;
    wire N__38291;
    wire N__38288;
    wire N__38285;
    wire N__38282;
    wire N__38279;
    wire N__38276;
    wire N__38273;
    wire N__38270;
    wire N__38267;
    wire N__38264;
    wire N__38257;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38247;
    wire N__38246;
    wire N__38245;
    wire N__38244;
    wire N__38243;
    wire N__38242;
    wire N__38239;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38222;
    wire N__38221;
    wire N__38218;
    wire N__38215;
    wire N__38212;
    wire N__38209;
    wire N__38204;
    wire N__38201;
    wire N__38196;
    wire N__38193;
    wire N__38188;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38170;
    wire N__38167;
    wire N__38164;
    wire N__38163;
    wire N__38160;
    wire N__38157;
    wire N__38154;
    wire N__38149;
    wire N__38146;
    wire N__38143;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38131;
    wire N__38128;
    wire N__38127;
    wire N__38122;
    wire N__38119;
    wire N__38116;
    wire N__38113;
    wire N__38110;
    wire N__38109;
    wire N__38108;
    wire N__38107;
    wire N__38104;
    wire N__38101;
    wire N__38098;
    wire N__38095;
    wire N__38088;
    wire N__38083;
    wire N__38080;
    wire N__38077;
    wire N__38074;
    wire N__38071;
    wire N__38070;
    wire N__38067;
    wire N__38064;
    wire N__38063;
    wire N__38060;
    wire N__38059;
    wire N__38056;
    wire N__38053;
    wire N__38050;
    wire N__38047;
    wire N__38046;
    wire N__38043;
    wire N__38040;
    wire N__38035;
    wire N__38032;
    wire N__38025;
    wire N__38020;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38008;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__37998;
    wire N__37993;
    wire N__37990;
    wire N__37987;
    wire N__37984;
    wire N__37981;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37960;
    wire N__37957;
    wire N__37954;
    wire N__37951;
    wire N__37948;
    wire N__37945;
    wire N__37944;
    wire N__37941;
    wire N__37940;
    wire N__37937;
    wire N__37934;
    wire N__37931;
    wire N__37928;
    wire N__37921;
    wire N__37918;
    wire N__37915;
    wire N__37914;
    wire N__37913;
    wire N__37910;
    wire N__37907;
    wire N__37904;
    wire N__37903;
    wire N__37896;
    wire N__37893;
    wire N__37890;
    wire N__37885;
    wire N__37882;
    wire N__37881;
    wire N__37880;
    wire N__37877;
    wire N__37876;
    wire N__37873;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37857;
    wire N__37852;
    wire N__37849;
    wire N__37848;
    wire N__37847;
    wire N__37846;
    wire N__37843;
    wire N__37840;
    wire N__37837;
    wire N__37834;
    wire N__37831;
    wire N__37828;
    wire N__37819;
    wire N__37818;
    wire N__37815;
    wire N__37812;
    wire N__37807;
    wire N__37804;
    wire N__37803;
    wire N__37800;
    wire N__37799;
    wire N__37796;
    wire N__37793;
    wire N__37790;
    wire N__37789;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37774;
    wire N__37769;
    wire N__37762;
    wire N__37759;
    wire N__37756;
    wire N__37753;
    wire N__37752;
    wire N__37751;
    wire N__37750;
    wire N__37747;
    wire N__37744;
    wire N__37741;
    wire N__37738;
    wire N__37735;
    wire N__37726;
    wire N__37723;
    wire N__37720;
    wire N__37717;
    wire N__37716;
    wire N__37715;
    wire N__37714;
    wire N__37711;
    wire N__37708;
    wire N__37703;
    wire N__37698;
    wire N__37693;
    wire N__37690;
    wire N__37687;
    wire N__37686;
    wire N__37685;
    wire N__37684;
    wire N__37681;
    wire N__37676;
    wire N__37673;
    wire N__37668;
    wire N__37663;
    wire N__37660;
    wire N__37657;
    wire N__37654;
    wire N__37653;
    wire N__37650;
    wire N__37645;
    wire N__37642;
    wire N__37641;
    wire N__37640;
    wire N__37637;
    wire N__37634;
    wire N__37631;
    wire N__37628;
    wire N__37621;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37609;
    wire N__37606;
    wire N__37605;
    wire N__37604;
    wire N__37603;
    wire N__37600;
    wire N__37593;
    wire N__37588;
    wire N__37585;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37570;
    wire N__37567;
    wire N__37564;
    wire N__37561;
    wire N__37558;
    wire N__37555;
    wire N__37552;
    wire N__37551;
    wire N__37546;
    wire N__37545;
    wire N__37542;
    wire N__37541;
    wire N__37538;
    wire N__37535;
    wire N__37532;
    wire N__37525;
    wire N__37522;
    wire N__37519;
    wire N__37516;
    wire N__37515;
    wire N__37514;
    wire N__37513;
    wire N__37510;
    wire N__37503;
    wire N__37502;
    wire N__37501;
    wire N__37496;
    wire N__37495;
    wire N__37494;
    wire N__37489;
    wire N__37486;
    wire N__37481;
    wire N__37474;
    wire N__37473;
    wire N__37472;
    wire N__37471;
    wire N__37470;
    wire N__37469;
    wire N__37468;
    wire N__37459;
    wire N__37454;
    wire N__37451;
    wire N__37446;
    wire N__37443;
    wire N__37440;
    wire N__37435;
    wire N__37432;
    wire N__37431;
    wire N__37430;
    wire N__37429;
    wire N__37428;
    wire N__37425;
    wire N__37424;
    wire N__37415;
    wire N__37410;
    wire N__37409;
    wire N__37404;
    wire N__37401;
    wire N__37398;
    wire N__37393;
    wire N__37390;
    wire N__37389;
    wire N__37388;
    wire N__37385;
    wire N__37382;
    wire N__37377;
    wire N__37372;
    wire N__37369;
    wire N__37366;
    wire N__37363;
    wire N__37360;
    wire N__37357;
    wire N__37356;
    wire N__37353;
    wire N__37350;
    wire N__37345;
    wire N__37342;
    wire N__37339;
    wire N__37336;
    wire N__37335;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37319;
    wire N__37318;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37302;
    wire N__37297;
    wire N__37294;
    wire N__37291;
    wire N__37288;
    wire N__37285;
    wire N__37282;
    wire N__37279;
    wire N__37276;
    wire N__37273;
    wire N__37270;
    wire N__37267;
    wire N__37264;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37254;
    wire N__37251;
    wire N__37250;
    wire N__37247;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37231;
    wire N__37222;
    wire N__37221;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37207;
    wire N__37204;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37194;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37176;
    wire N__37171;
    wire N__37170;
    wire N__37167;
    wire N__37164;
    wire N__37161;
    wire N__37158;
    wire N__37155;
    wire N__37152;
    wire N__37147;
    wire N__37146;
    wire N__37143;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37135;
    wire N__37132;
    wire N__37129;
    wire N__37126;
    wire N__37123;
    wire N__37118;
    wire N__37111;
    wire N__37108;
    wire N__37105;
    wire N__37102;
    wire N__37099;
    wire N__37098;
    wire N__37095;
    wire N__37092;
    wire N__37089;
    wire N__37084;
    wire N__37083;
    wire N__37080;
    wire N__37077;
    wire N__37072;
    wire N__37071;
    wire N__37068;
    wire N__37065;
    wire N__37062;
    wire N__37061;
    wire N__37060;
    wire N__37057;
    wire N__37054;
    wire N__37051;
    wire N__37048;
    wire N__37047;
    wire N__37046;
    wire N__37043;
    wire N__37036;
    wire N__37033;
    wire N__37030;
    wire N__37025;
    wire N__37018;
    wire N__37015;
    wire N__37014;
    wire N__37011;
    wire N__37008;
    wire N__37005;
    wire N__37000;
    wire N__36997;
    wire N__36994;
    wire N__36993;
    wire N__36990;
    wire N__36987;
    wire N__36986;
    wire N__36985;
    wire N__36982;
    wire N__36979;
    wire N__36974;
    wire N__36971;
    wire N__36968;
    wire N__36961;
    wire N__36960;
    wire N__36957;
    wire N__36952;
    wire N__36949;
    wire N__36948;
    wire N__36947;
    wire N__36944;
    wire N__36941;
    wire N__36938;
    wire N__36933;
    wire N__36928;
    wire N__36925;
    wire N__36924;
    wire N__36921;
    wire N__36918;
    wire N__36915;
    wire N__36910;
    wire N__36909;
    wire N__36908;
    wire N__36907;
    wire N__36906;
    wire N__36903;
    wire N__36902;
    wire N__36901;
    wire N__36900;
    wire N__36899;
    wire N__36898;
    wire N__36897;
    wire N__36896;
    wire N__36895;
    wire N__36894;
    wire N__36891;
    wire N__36890;
    wire N__36889;
    wire N__36888;
    wire N__36887;
    wire N__36884;
    wire N__36883;
    wire N__36882;
    wire N__36877;
    wire N__36874;
    wire N__36873;
    wire N__36872;
    wire N__36871;
    wire N__36870;
    wire N__36867;
    wire N__36864;
    wire N__36863;
    wire N__36862;
    wire N__36859;
    wire N__36854;
    wire N__36849;
    wire N__36848;
    wire N__36847;
    wire N__36844;
    wire N__36841;
    wire N__36838;
    wire N__36835;
    wire N__36834;
    wire N__36833;
    wire N__36830;
    wire N__36825;
    wire N__36822;
    wire N__36819;
    wire N__36818;
    wire N__36817;
    wire N__36814;
    wire N__36809;
    wire N__36800;
    wire N__36797;
    wire N__36788;
    wire N__36783;
    wire N__36778;
    wire N__36769;
    wire N__36766;
    wire N__36765;
    wire N__36762;
    wire N__36761;
    wire N__36760;
    wire N__36759;
    wire N__36756;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36742;
    wire N__36741;
    wire N__36738;
    wire N__36733;
    wire N__36728;
    wire N__36721;
    wire N__36718;
    wire N__36715;
    wire N__36712;
    wire N__36705;
    wire N__36698;
    wire N__36695;
    wire N__36692;
    wire N__36689;
    wire N__36682;
    wire N__36679;
    wire N__36676;
    wire N__36665;
    wire N__36652;
    wire N__36649;
    wire N__36646;
    wire N__36645;
    wire N__36644;
    wire N__36643;
    wire N__36638;
    wire N__36633;
    wire N__36630;
    wire N__36625;
    wire N__36624;
    wire N__36623;
    wire N__36620;
    wire N__36617;
    wire N__36614;
    wire N__36611;
    wire N__36608;
    wire N__36605;
    wire N__36600;
    wire N__36595;
    wire N__36594;
    wire N__36591;
    wire N__36588;
    wire N__36587;
    wire N__36586;
    wire N__36583;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36571;
    wire N__36566;
    wire N__36559;
    wire N__36558;
    wire N__36557;
    wire N__36556;
    wire N__36553;
    wire N__36550;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36540;
    wire N__36537;
    wire N__36532;
    wire N__36531;
    wire N__36530;
    wire N__36527;
    wire N__36522;
    wire N__36519;
    wire N__36514;
    wire N__36505;
    wire N__36504;
    wire N__36503;
    wire N__36500;
    wire N__36499;
    wire N__36496;
    wire N__36495;
    wire N__36492;
    wire N__36489;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36477;
    wire N__36472;
    wire N__36469;
    wire N__36460;
    wire N__36459;
    wire N__36458;
    wire N__36455;
    wire N__36454;
    wire N__36451;
    wire N__36446;
    wire N__36443;
    wire N__36440;
    wire N__36433;
    wire N__36430;
    wire N__36427;
    wire N__36426;
    wire N__36425;
    wire N__36422;
    wire N__36419;
    wire N__36416;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36406;
    wire N__36403;
    wire N__36398;
    wire N__36395;
    wire N__36392;
    wire N__36389;
    wire N__36382;
    wire N__36381;
    wire N__36378;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36368;
    wire N__36367;
    wire N__36364;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36350;
    wire N__36343;
    wire N__36340;
    wire N__36337;
    wire N__36334;
    wire N__36331;
    wire N__36328;
    wire N__36325;
    wire N__36324;
    wire N__36323;
    wire N__36320;
    wire N__36315;
    wire N__36310;
    wire N__36307;
    wire N__36304;
    wire N__36301;
    wire N__36300;
    wire N__36299;
    wire N__36296;
    wire N__36291;
    wire N__36286;
    wire N__36285;
    wire N__36282;
    wire N__36279;
    wire N__36276;
    wire N__36271;
    wire N__36268;
    wire N__36265;
    wire N__36262;
    wire N__36259;
    wire N__36258;
    wire N__36257;
    wire N__36256;
    wire N__36253;
    wire N__36252;
    wire N__36249;
    wire N__36246;
    wire N__36243;
    wire N__36240;
    wire N__36237;
    wire N__36234;
    wire N__36231;
    wire N__36220;
    wire N__36217;
    wire N__36216;
    wire N__36213;
    wire N__36210;
    wire N__36207;
    wire N__36204;
    wire N__36201;
    wire N__36198;
    wire N__36197;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36185;
    wire N__36178;
    wire N__36175;
    wire N__36172;
    wire N__36169;
    wire N__36166;
    wire N__36165;
    wire N__36160;
    wire N__36159;
    wire N__36156;
    wire N__36155;
    wire N__36154;
    wire N__36151;
    wire N__36148;
    wire N__36143;
    wire N__36136;
    wire N__36133;
    wire N__36130;
    wire N__36127;
    wire N__36124;
    wire N__36123;
    wire N__36122;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36112;
    wire N__36111;
    wire N__36108;
    wire N__36105;
    wire N__36100;
    wire N__36097;
    wire N__36088;
    wire N__36085;
    wire N__36082;
    wire N__36079;
    wire N__36078;
    wire N__36075;
    wire N__36072;
    wire N__36069;
    wire N__36066;
    wire N__36063;
    wire N__36062;
    wire N__36059;
    wire N__36058;
    wire N__36057;
    wire N__36056;
    wire N__36053;
    wire N__36050;
    wire N__36047;
    wire N__36044;
    wire N__36039;
    wire N__36028;
    wire N__36027;
    wire N__36024;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36010;
    wire N__36007;
    wire N__36004;
    wire N__36001;
    wire N__35998;
    wire N__35997;
    wire N__35994;
    wire N__35993;
    wire N__35990;
    wire N__35989;
    wire N__35986;
    wire N__35983;
    wire N__35980;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35967;
    wire N__35964;
    wire N__35953;
    wire N__35950;
    wire N__35947;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35932;
    wire N__35929;
    wire N__35928;
    wire N__35925;
    wire N__35922;
    wire N__35919;
    wire N__35916;
    wire N__35911;
    wire N__35908;
    wire N__35905;
    wire N__35902;
    wire N__35899;
    wire N__35896;
    wire N__35895;
    wire N__35892;
    wire N__35891;
    wire N__35890;
    wire N__35887;
    wire N__35884;
    wire N__35881;
    wire N__35878;
    wire N__35877;
    wire N__35874;
    wire N__35873;
    wire N__35872;
    wire N__35869;
    wire N__35866;
    wire N__35861;
    wire N__35858;
    wire N__35853;
    wire N__35842;
    wire N__35839;
    wire N__35836;
    wire N__35833;
    wire N__35830;
    wire N__35827;
    wire N__35824;
    wire N__35821;
    wire N__35818;
    wire N__35815;
    wire N__35812;
    wire N__35811;
    wire N__35810;
    wire N__35807;
    wire N__35804;
    wire N__35801;
    wire N__35794;
    wire N__35791;
    wire N__35788;
    wire N__35787;
    wire N__35784;
    wire N__35781;
    wire N__35776;
    wire N__35773;
    wire N__35772;
    wire N__35769;
    wire N__35766;
    wire N__35765;
    wire N__35764;
    wire N__35763;
    wire N__35762;
    wire N__35759;
    wire N__35756;
    wire N__35753;
    wire N__35750;
    wire N__35747;
    wire N__35744;
    wire N__35739;
    wire N__35728;
    wire N__35725;
    wire N__35724;
    wire N__35723;
    wire N__35720;
    wire N__35717;
    wire N__35714;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35704;
    wire N__35703;
    wire N__35702;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35690;
    wire N__35687;
    wire N__35684;
    wire N__35681;
    wire N__35668;
    wire N__35665;
    wire N__35662;
    wire N__35659;
    wire N__35656;
    wire N__35655;
    wire N__35652;
    wire N__35649;
    wire N__35646;
    wire N__35645;
    wire N__35644;
    wire N__35641;
    wire N__35638;
    wire N__35635;
    wire N__35632;
    wire N__35629;
    wire N__35624;
    wire N__35619;
    wire N__35614;
    wire N__35611;
    wire N__35610;
    wire N__35609;
    wire N__35606;
    wire N__35605;
    wire N__35600;
    wire N__35597;
    wire N__35594;
    wire N__35591;
    wire N__35590;
    wire N__35587;
    wire N__35582;
    wire N__35579;
    wire N__35572;
    wire N__35569;
    wire N__35568;
    wire N__35565;
    wire N__35562;
    wire N__35559;
    wire N__35556;
    wire N__35553;
    wire N__35550;
    wire N__35545;
    wire N__35542;
    wire N__35539;
    wire N__35536;
    wire N__35533;
    wire N__35530;
    wire N__35529;
    wire N__35526;
    wire N__35523;
    wire N__35520;
    wire N__35519;
    wire N__35518;
    wire N__35517;
    wire N__35514;
    wire N__35511;
    wire N__35508;
    wire N__35505;
    wire N__35502;
    wire N__35499;
    wire N__35496;
    wire N__35493;
    wire N__35486;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35470;
    wire N__35467;
    wire N__35464;
    wire N__35461;
    wire N__35458;
    wire N__35455;
    wire N__35452;
    wire N__35449;
    wire N__35446;
    wire N__35445;
    wire N__35442;
    wire N__35439;
    wire N__35434;
    wire N__35431;
    wire N__35428;
    wire N__35425;
    wire N__35422;
    wire N__35419;
    wire N__35418;
    wire N__35415;
    wire N__35412;
    wire N__35409;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35391;
    wire N__35390;
    wire N__35387;
    wire N__35386;
    wire N__35385;
    wire N__35382;
    wire N__35381;
    wire N__35378;
    wire N__35375;
    wire N__35370;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35360;
    wire N__35355;
    wire N__35352;
    wire N__35341;
    wire N__35338;
    wire N__35335;
    wire N__35334;
    wire N__35331;
    wire N__35328;
    wire N__35325;
    wire N__35320;
    wire N__35317;
    wire N__35316;
    wire N__35311;
    wire N__35310;
    wire N__35309;
    wire N__35308;
    wire N__35305;
    wire N__35300;
    wire N__35297;
    wire N__35294;
    wire N__35289;
    wire N__35284;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35274;
    wire N__35271;
    wire N__35268;
    wire N__35265;
    wire N__35260;
    wire N__35257;
    wire N__35254;
    wire N__35253;
    wire N__35252;
    wire N__35249;
    wire N__35246;
    wire N__35245;
    wire N__35242;
    wire N__35239;
    wire N__35236;
    wire N__35233;
    wire N__35226;
    wire N__35221;
    wire N__35220;
    wire N__35217;
    wire N__35214;
    wire N__35213;
    wire N__35210;
    wire N__35209;
    wire N__35208;
    wire N__35205;
    wire N__35202;
    wire N__35201;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35191;
    wire N__35186;
    wire N__35181;
    wire N__35170;
    wire N__35169;
    wire N__35166;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35149;
    wire N__35146;
    wire N__35143;
    wire N__35140;
    wire N__35139;
    wire N__35136;
    wire N__35135;
    wire N__35134;
    wire N__35131;
    wire N__35128;
    wire N__35123;
    wire N__35122;
    wire N__35121;
    wire N__35120;
    wire N__35117;
    wire N__35116;
    wire N__35111;
    wire N__35108;
    wire N__35103;
    wire N__35100;
    wire N__35097;
    wire N__35094;
    wire N__35091;
    wire N__35080;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35065;
    wire N__35064;
    wire N__35061;
    wire N__35058;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35043;
    wire N__35042;
    wire N__35039;
    wire N__35036;
    wire N__35035;
    wire N__35032;
    wire N__35031;
    wire N__35030;
    wire N__35027;
    wire N__35024;
    wire N__35021;
    wire N__35016;
    wire N__35013;
    wire N__35002;
    wire N__34999;
    wire N__34998;
    wire N__34995;
    wire N__34992;
    wire N__34989;
    wire N__34984;
    wire N__34981;
    wire N__34980;
    wire N__34979;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34967;
    wire N__34966;
    wire N__34963;
    wire N__34958;
    wire N__34957;
    wire N__34954;
    wire N__34949;
    wire N__34946;
    wire N__34943;
    wire N__34940;
    wire N__34933;
    wire N__34930;
    wire N__34929;
    wire N__34928;
    wire N__34927;
    wire N__34926;
    wire N__34925;
    wire N__34922;
    wire N__34919;
    wire N__34916;
    wire N__34913;
    wire N__34908;
    wire N__34907;
    wire N__34904;
    wire N__34901;
    wire N__34898;
    wire N__34893;
    wire N__34890;
    wire N__34887;
    wire N__34884;
    wire N__34879;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34850;
    wire N__34845;
    wire N__34842;
    wire N__34839;
    wire N__34834;
    wire N__34831;
    wire N__34828;
    wire N__34827;
    wire N__34824;
    wire N__34821;
    wire N__34818;
    wire N__34817;
    wire N__34814;
    wire N__34811;
    wire N__34808;
    wire N__34801;
    wire N__34798;
    wire N__34795;
    wire N__34794;
    wire N__34793;
    wire N__34792;
    wire N__34789;
    wire N__34784;
    wire N__34781;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34756;
    wire N__34753;
    wire N__34750;
    wire N__34747;
    wire N__34744;
    wire N__34741;
    wire N__34738;
    wire N__34735;
    wire N__34732;
    wire N__34731;
    wire N__34728;
    wire N__34725;
    wire N__34722;
    wire N__34717;
    wire N__34714;
    wire N__34711;
    wire N__34710;
    wire N__34707;
    wire N__34704;
    wire N__34701;
    wire N__34696;
    wire N__34693;
    wire N__34690;
    wire N__34687;
    wire N__34684;
    wire N__34681;
    wire N__34678;
    wire N__34675;
    wire N__34672;
    wire N__34669;
    wire N__34668;
    wire N__34665;
    wire N__34662;
    wire N__34659;
    wire N__34654;
    wire N__34651;
    wire N__34648;
    wire N__34645;
    wire N__34642;
    wire N__34639;
    wire N__34636;
    wire N__34635;
    wire N__34632;
    wire N__34631;
    wire N__34628;
    wire N__34627;
    wire N__34624;
    wire N__34623;
    wire N__34622;
    wire N__34621;
    wire N__34618;
    wire N__34615;
    wire N__34612;
    wire N__34609;
    wire N__34602;
    wire N__34595;
    wire N__34588;
    wire N__34585;
    wire N__34584;
    wire N__34579;
    wire N__34576;
    wire N__34573;
    wire N__34570;
    wire N__34567;
    wire N__34566;
    wire N__34565;
    wire N__34564;
    wire N__34559;
    wire N__34556;
    wire N__34553;
    wire N__34550;
    wire N__34543;
    wire N__34542;
    wire N__34541;
    wire N__34540;
    wire N__34537;
    wire N__34534;
    wire N__34531;
    wire N__34526;
    wire N__34523;
    wire N__34516;
    wire N__34513;
    wire N__34510;
    wire N__34507;
    wire N__34504;
    wire N__34503;
    wire N__34502;
    wire N__34497;
    wire N__34494;
    wire N__34491;
    wire N__34486;
    wire N__34483;
    wire N__34480;
    wire N__34477;
    wire N__34476;
    wire N__34473;
    wire N__34470;
    wire N__34467;
    wire N__34464;
    wire N__34459;
    wire N__34456;
    wire N__34455;
    wire N__34454;
    wire N__34453;
    wire N__34452;
    wire N__34449;
    wire N__34446;
    wire N__34445;
    wire N__34438;
    wire N__34433;
    wire N__34430;
    wire N__34427;
    wire N__34426;
    wire N__34421;
    wire N__34418;
    wire N__34415;
    wire N__34412;
    wire N__34409;
    wire N__34406;
    wire N__34399;
    wire N__34398;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34388;
    wire N__34387;
    wire N__34386;
    wire N__34383;
    wire N__34380;
    wire N__34373;
    wire N__34366;
    wire N__34363;
    wire N__34362;
    wire N__34359;
    wire N__34356;
    wire N__34353;
    wire N__34348;
    wire N__34345;
    wire N__34344;
    wire N__34343;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34329;
    wire N__34326;
    wire N__34323;
    wire N__34318;
    wire N__34315;
    wire N__34312;
    wire N__34309;
    wire N__34308;
    wire N__34303;
    wire N__34302;
    wire N__34301;
    wire N__34298;
    wire N__34295;
    wire N__34292;
    wire N__34289;
    wire N__34282;
    wire N__34279;
    wire N__34278;
    wire N__34277;
    wire N__34274;
    wire N__34269;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34252;
    wire N__34249;
    wire N__34248;
    wire N__34247;
    wire N__34246;
    wire N__34241;
    wire N__34238;
    wire N__34235;
    wire N__34232;
    wire N__34229;
    wire N__34222;
    wire N__34219;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34204;
    wire N__34201;
    wire N__34198;
    wire N__34197;
    wire N__34194;
    wire N__34193;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34177;
    wire N__34172;
    wire N__34165;
    wire N__34164;
    wire N__34161;
    wire N__34158;
    wire N__34157;
    wire N__34156;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34132;
    wire N__34129;
    wire N__34126;
    wire N__34123;
    wire N__34120;
    wire N__34119;
    wire N__34116;
    wire N__34113;
    wire N__34110;
    wire N__34105;
    wire N__34102;
    wire N__34101;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34087;
    wire N__34084;
    wire N__34081;
    wire N__34080;
    wire N__34077;
    wire N__34074;
    wire N__34071;
    wire N__34066;
    wire N__34063;
    wire N__34062;
    wire N__34059;
    wire N__34056;
    wire N__34053;
    wire N__34048;
    wire N__34045;
    wire N__34042;
    wire N__34039;
    wire N__34036;
    wire N__34033;
    wire N__34030;
    wire N__34027;
    wire N__34024;
    wire N__34023;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34009;
    wire N__34006;
    wire N__34005;
    wire N__34000;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33985;
    wire N__33982;
    wire N__33979;
    wire N__33976;
    wire N__33975;
    wire N__33972;
    wire N__33971;
    wire N__33970;
    wire N__33969;
    wire N__33968;
    wire N__33967;
    wire N__33966;
    wire N__33965;
    wire N__33964;
    wire N__33963;
    wire N__33960;
    wire N__33959;
    wire N__33956;
    wire N__33949;
    wire N__33948;
    wire N__33947;
    wire N__33946;
    wire N__33945;
    wire N__33944;
    wire N__33943;
    wire N__33942;
    wire N__33939;
    wire N__33938;
    wire N__33937;
    wire N__33932;
    wire N__33927;
    wire N__33924;
    wire N__33919;
    wire N__33914;
    wire N__33907;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33889;
    wire N__33888;
    wire N__33887;
    wire N__33886;
    wire N__33883;
    wire N__33870;
    wire N__33865;
    wire N__33864;
    wire N__33863;
    wire N__33858;
    wire N__33855;
    wire N__33854;
    wire N__33845;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33823;
    wire N__33816;
    wire N__33805;
    wire N__33804;
    wire N__33801;
    wire N__33798;
    wire N__33795;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33775;
    wire N__33772;
    wire N__33771;
    wire N__33770;
    wire N__33769;
    wire N__33768;
    wire N__33767;
    wire N__33764;
    wire N__33763;
    wire N__33760;
    wire N__33757;
    wire N__33756;
    wire N__33749;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33734;
    wire N__33731;
    wire N__33722;
    wire N__33719;
    wire N__33716;
    wire N__33713;
    wire N__33706;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33693;
    wire N__33692;
    wire N__33691;
    wire N__33690;
    wire N__33689;
    wire N__33688;
    wire N__33687;
    wire N__33686;
    wire N__33685;
    wire N__33684;
    wire N__33683;
    wire N__33682;
    wire N__33681;
    wire N__33680;
    wire N__33679;
    wire N__33678;
    wire N__33677;
    wire N__33676;
    wire N__33673;
    wire N__33672;
    wire N__33669;
    wire N__33668;
    wire N__33665;
    wire N__33664;
    wire N__33663;
    wire N__33660;
    wire N__33657;
    wire N__33656;
    wire N__33653;
    wire N__33652;
    wire N__33649;
    wire N__33648;
    wire N__33645;
    wire N__33644;
    wire N__33641;
    wire N__33640;
    wire N__33637;
    wire N__33636;
    wire N__33633;
    wire N__33632;
    wire N__33629;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33619;
    wire N__33616;
    wire N__33613;
    wire N__33610;
    wire N__33607;
    wire N__33606;
    wire N__33605;
    wire N__33592;
    wire N__33587;
    wire N__33570;
    wire N__33553;
    wire N__33544;
    wire N__33535;
    wire N__33532;
    wire N__33527;
    wire N__33522;
    wire N__33517;
    wire N__33514;
    wire N__33509;
    wire N__33506;
    wire N__33499;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33489;
    wire N__33484;
    wire N__33481;
    wire N__33478;
    wire N__33475;
    wire N__33474;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33460;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33448;
    wire N__33445;
    wire N__33442;
    wire N__33439;
    wire N__33436;
    wire N__33433;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33423;
    wire N__33418;
    wire N__33415;
    wire N__33414;
    wire N__33409;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33391;
    wire N__33388;
    wire N__33387;
    wire N__33386;
    wire N__33383;
    wire N__33380;
    wire N__33377;
    wire N__33376;
    wire N__33373;
    wire N__33370;
    wire N__33367;
    wire N__33366;
    wire N__33363;
    wire N__33358;
    wire N__33355;
    wire N__33350;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33334;
    wire N__33331;
    wire N__33328;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33292;
    wire N__33289;
    wire N__33286;
    wire N__33283;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33271;
    wire N__33268;
    wire N__33265;
    wire N__33262;
    wire N__33259;
    wire N__33256;
    wire N__33253;
    wire N__33250;
    wire N__33249;
    wire N__33246;
    wire N__33245;
    wire N__33244;
    wire N__33243;
    wire N__33240;
    wire N__33237;
    wire N__33234;
    wire N__33231;
    wire N__33230;
    wire N__33227;
    wire N__33222;
    wire N__33219;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33199;
    wire N__33196;
    wire N__33193;
    wire N__33190;
    wire N__33187;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33162;
    wire N__33161;
    wire N__33160;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33085;
    wire N__33084;
    wire N__33081;
    wire N__33078;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33064;
    wire N__33061;
    wire N__33060;
    wire N__33059;
    wire N__33058;
    wire N__33057;
    wire N__33056;
    wire N__33051;
    wire N__33050;
    wire N__33043;
    wire N__33040;
    wire N__33037;
    wire N__33034;
    wire N__33031;
    wire N__33022;
    wire N__33019;
    wire N__33018;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32980;
    wire N__32979;
    wire N__32976;
    wire N__32975;
    wire N__32972;
    wire N__32969;
    wire N__32966;
    wire N__32965;
    wire N__32962;
    wire N__32959;
    wire N__32956;
    wire N__32955;
    wire N__32952;
    wire N__32945;
    wire N__32942;
    wire N__32935;
    wire N__32932;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32920;
    wire N__32919;
    wire N__32918;
    wire N__32915;
    wire N__32910;
    wire N__32905;
    wire N__32902;
    wire N__32901;
    wire N__32900;
    wire N__32897;
    wire N__32894;
    wire N__32893;
    wire N__32892;
    wire N__32889;
    wire N__32886;
    wire N__32883;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32868;
    wire N__32857;
    wire N__32856;
    wire N__32853;
    wire N__32852;
    wire N__32849;
    wire N__32846;
    wire N__32845;
    wire N__32842;
    wire N__32839;
    wire N__32836;
    wire N__32833;
    wire N__32824;
    wire N__32823;
    wire N__32820;
    wire N__32817;
    wire N__32816;
    wire N__32811;
    wire N__32808;
    wire N__32805;
    wire N__32800;
    wire N__32799;
    wire N__32796;
    wire N__32793;
    wire N__32792;
    wire N__32791;
    wire N__32790;
    wire N__32789;
    wire N__32786;
    wire N__32785;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32773;
    wire N__32770;
    wire N__32767;
    wire N__32764;
    wire N__32761;
    wire N__32758;
    wire N__32753;
    wire N__32740;
    wire N__32739;
    wire N__32738;
    wire N__32735;
    wire N__32734;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32726;
    wire N__32725;
    wire N__32724;
    wire N__32721;
    wire N__32718;
    wire N__32715;
    wire N__32712;
    wire N__32705;
    wire N__32704;
    wire N__32701;
    wire N__32700;
    wire N__32697;
    wire N__32694;
    wire N__32691;
    wire N__32688;
    wire N__32685;
    wire N__32680;
    wire N__32677;
    wire N__32670;
    wire N__32667;
    wire N__32662;
    wire N__32653;
    wire N__32650;
    wire N__32647;
    wire N__32644;
    wire N__32641;
    wire N__32638;
    wire N__32637;
    wire N__32634;
    wire N__32631;
    wire N__32626;
    wire N__32623;
    wire N__32620;
    wire N__32617;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32607;
    wire N__32604;
    wire N__32601;
    wire N__32598;
    wire N__32593;
    wire N__32592;
    wire N__32589;
    wire N__32586;
    wire N__32583;
    wire N__32580;
    wire N__32577;
    wire N__32572;
    wire N__32569;
    wire N__32566;
    wire N__32565;
    wire N__32562;
    wire N__32561;
    wire N__32558;
    wire N__32555;
    wire N__32554;
    wire N__32553;
    wire N__32552;
    wire N__32549;
    wire N__32544;
    wire N__32541;
    wire N__32538;
    wire N__32535;
    wire N__32526;
    wire N__32521;
    wire N__32518;
    wire N__32517;
    wire N__32516;
    wire N__32513;
    wire N__32512;
    wire N__32509;
    wire N__32506;
    wire N__32505;
    wire N__32502;
    wire N__32499;
    wire N__32498;
    wire N__32495;
    wire N__32494;
    wire N__32493;
    wire N__32490;
    wire N__32487;
    wire N__32482;
    wire N__32479;
    wire N__32476;
    wire N__32473;
    wire N__32470;
    wire N__32465;
    wire N__32460;
    wire N__32449;
    wire N__32448;
    wire N__32447;
    wire N__32446;
    wire N__32443;
    wire N__32442;
    wire N__32439;
    wire N__32434;
    wire N__32431;
    wire N__32428;
    wire N__32425;
    wire N__32422;
    wire N__32421;
    wire N__32420;
    wire N__32417;
    wire N__32414;
    wire N__32411;
    wire N__32408;
    wire N__32403;
    wire N__32398;
    wire N__32389;
    wire N__32386;
    wire N__32385;
    wire N__32384;
    wire N__32381;
    wire N__32380;
    wire N__32377;
    wire N__32374;
    wire N__32373;
    wire N__32372;
    wire N__32371;
    wire N__32368;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32346;
    wire N__32343;
    wire N__32334;
    wire N__32323;
    wire N__32320;
    wire N__32317;
    wire N__32314;
    wire N__32311;
    wire N__32310;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32302;
    wire N__32299;
    wire N__32296;
    wire N__32293;
    wire N__32290;
    wire N__32287;
    wire N__32286;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32274;
    wire N__32273;
    wire N__32270;
    wire N__32263;
    wire N__32260;
    wire N__32257;
    wire N__32248;
    wire N__32247;
    wire N__32246;
    wire N__32245;
    wire N__32242;
    wire N__32237;
    wire N__32234;
    wire N__32233;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32212;
    wire N__32211;
    wire N__32210;
    wire N__32207;
    wire N__32206;
    wire N__32205;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32190;
    wire N__32187;
    wire N__32186;
    wire N__32179;
    wire N__32176;
    wire N__32173;
    wire N__32170;
    wire N__32167;
    wire N__32162;
    wire N__32159;
    wire N__32152;
    wire N__32149;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32141;
    wire N__32136;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32116;
    wire N__32115;
    wire N__32114;
    wire N__32113;
    wire N__32110;
    wire N__32109;
    wire N__32106;
    wire N__32101;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32089;
    wire N__32086;
    wire N__32083;
    wire N__32080;
    wire N__32075;
    wire N__32068;
    wire N__32065;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32055;
    wire N__32050;
    wire N__32047;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32039;
    wire N__32036;
    wire N__32035;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32021;
    wire N__32014;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32002;
    wire N__31999;
    wire N__31996;
    wire N__31993;
    wire N__31990;
    wire N__31989;
    wire N__31988;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31974;
    wire N__31969;
    wire N__31968;
    wire N__31965;
    wire N__31964;
    wire N__31961;
    wire N__31958;
    wire N__31957;
    wire N__31956;
    wire N__31953;
    wire N__31948;
    wire N__31943;
    wire N__31940;
    wire N__31935;
    wire N__31930;
    wire N__31927;
    wire N__31926;
    wire N__31923;
    wire N__31922;
    wire N__31919;
    wire N__31916;
    wire N__31913;
    wire N__31912;
    wire N__31909;
    wire N__31904;
    wire N__31901;
    wire N__31894;
    wire N__31893;
    wire N__31892;
    wire N__31887;
    wire N__31886;
    wire N__31883;
    wire N__31882;
    wire N__31881;
    wire N__31878;
    wire N__31877;
    wire N__31872;
    wire N__31867;
    wire N__31864;
    wire N__31861;
    wire N__31852;
    wire N__31849;
    wire N__31846;
    wire N__31843;
    wire N__31840;
    wire N__31839;
    wire N__31838;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31824;
    wire N__31821;
    wire N__31818;
    wire N__31813;
    wire N__31810;
    wire N__31807;
    wire N__31804;
    wire N__31801;
    wire N__31798;
    wire N__31797;
    wire N__31794;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31777;
    wire N__31774;
    wire N__31771;
    wire N__31770;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31757;
    wire N__31754;
    wire N__31751;
    wire N__31748;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31729;
    wire N__31728;
    wire N__31723;
    wire N__31720;
    wire N__31719;
    wire N__31714;
    wire N__31711;
    wire N__31708;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31696;
    wire N__31693;
    wire N__31692;
    wire N__31689;
    wire N__31688;
    wire N__31687;
    wire N__31684;
    wire N__31683;
    wire N__31682;
    wire N__31679;
    wire N__31676;
    wire N__31673;
    wire N__31670;
    wire N__31667;
    wire N__31664;
    wire N__31657;
    wire N__31656;
    wire N__31653;
    wire N__31646;
    wire N__31643;
    wire N__31636;
    wire N__31635;
    wire N__31634;
    wire N__31633;
    wire N__31632;
    wire N__31631;
    wire N__31630;
    wire N__31627;
    wire N__31624;
    wire N__31623;
    wire N__31618;
    wire N__31613;
    wire N__31610;
    wire N__31607;
    wire N__31604;
    wire N__31601;
    wire N__31594;
    wire N__31587;
    wire N__31582;
    wire N__31579;
    wire N__31576;
    wire N__31573;
    wire N__31570;
    wire N__31569;
    wire N__31566;
    wire N__31565;
    wire N__31562;
    wire N__31561;
    wire N__31558;
    wire N__31555;
    wire N__31552;
    wire N__31549;
    wire N__31540;
    wire N__31537;
    wire N__31536;
    wire N__31531;
    wire N__31528;
    wire N__31527;
    wire N__31522;
    wire N__31519;
    wire N__31516;
    wire N__31515;
    wire N__31510;
    wire N__31507;
    wire N__31504;
    wire N__31501;
    wire N__31498;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31486;
    wire N__31485;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31468;
    wire N__31465;
    wire N__31462;
    wire N__31459;
    wire N__31458;
    wire N__31457;
    wire N__31454;
    wire N__31451;
    wire N__31448;
    wire N__31441;
    wire N__31438;
    wire N__31435;
    wire N__31434;
    wire N__31431;
    wire N__31428;
    wire N__31425;
    wire N__31420;
    wire N__31419;
    wire N__31418;
    wire N__31417;
    wire N__31416;
    wire N__31415;
    wire N__31412;
    wire N__31409;
    wire N__31406;
    wire N__31405;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31391;
    wire N__31386;
    wire N__31383;
    wire N__31378;
    wire N__31377;
    wire N__31374;
    wire N__31367;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31351;
    wire N__31350;
    wire N__31349;
    wire N__31348;
    wire N__31345;
    wire N__31342;
    wire N__31341;
    wire N__31338;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31325;
    wire N__31322;
    wire N__31319;
    wire N__31316;
    wire N__31313;
    wire N__31310;
    wire N__31297;
    wire N__31296;
    wire N__31295;
    wire N__31294;
    wire N__31289;
    wire N__31286;
    wire N__31285;
    wire N__31282;
    wire N__31277;
    wire N__31274;
    wire N__31273;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31263;
    wire N__31258;
    wire N__31257;
    wire N__31256;
    wire N__31253;
    wire N__31252;
    wire N__31249;
    wire N__31244;
    wire N__31241;
    wire N__31238;
    wire N__31235;
    wire N__31232;
    wire N__31219;
    wire N__31218;
    wire N__31217;
    wire N__31214;
    wire N__31213;
    wire N__31210;
    wire N__31209;
    wire N__31208;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31190;
    wire N__31185;
    wire N__31182;
    wire N__31177;
    wire N__31174;
    wire N__31171;
    wire N__31166;
    wire N__31159;
    wire N__31158;
    wire N__31153;
    wire N__31152;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31142;
    wire N__31139;
    wire N__31132;
    wire N__31131;
    wire N__31130;
    wire N__31129;
    wire N__31128;
    wire N__31123;
    wire N__31120;
    wire N__31115;
    wire N__31110;
    wire N__31107;
    wire N__31102;
    wire N__31099;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31089;
    wire N__31088;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31072;
    wire N__31071;
    wire N__31070;
    wire N__31067;
    wire N__31064;
    wire N__31061;
    wire N__31054;
    wire N__31051;
    wire N__31048;
    wire N__31047;
    wire N__31044;
    wire N__31043;
    wire N__31042;
    wire N__31039;
    wire N__31036;
    wire N__31031;
    wire N__31024;
    wire N__31021;
    wire N__31018;
    wire N__31015;
    wire N__31012;
    wire N__31009;
    wire N__31006;
    wire N__31003;
    wire N__31000;
    wire N__30997;
    wire N__30994;
    wire N__30991;
    wire N__30988;
    wire N__30985;
    wire N__30982;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30967;
    wire N__30964;
    wire N__30961;
    wire N__30958;
    wire N__30955;
    wire N__30952;
    wire N__30949;
    wire N__30946;
    wire N__30943;
    wire N__30940;
    wire N__30937;
    wire N__30934;
    wire N__30933;
    wire N__30930;
    wire N__30929;
    wire N__30926;
    wire N__30923;
    wire N__30920;
    wire N__30915;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30898;
    wire N__30897;
    wire N__30896;
    wire N__30893;
    wire N__30890;
    wire N__30887;
    wire N__30880;
    wire N__30877;
    wire N__30874;
    wire N__30871;
    wire N__30870;
    wire N__30869;
    wire N__30866;
    wire N__30863;
    wire N__30860;
    wire N__30853;
    wire N__30850;
    wire N__30847;
    wire N__30844;
    wire N__30843;
    wire N__30842;
    wire N__30839;
    wire N__30836;
    wire N__30833;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30816;
    wire N__30813;
    wire N__30810;
    wire N__30809;
    wire N__30804;
    wire N__30801;
    wire N__30798;
    wire N__30793;
    wire N__30790;
    wire N__30787;
    wire N__30784;
    wire N__30781;
    wire N__30780;
    wire N__30779;
    wire N__30778;
    wire N__30775;
    wire N__30772;
    wire N__30767;
    wire N__30760;
    wire N__30757;
    wire N__30754;
    wire N__30751;
    wire N__30748;
    wire N__30745;
    wire N__30742;
    wire N__30739;
    wire N__30736;
    wire N__30735;
    wire N__30732;
    wire N__30731;
    wire N__30730;
    wire N__30729;
    wire N__30722;
    wire N__30721;
    wire N__30720;
    wire N__30715;
    wire N__30712;
    wire N__30711;
    wire N__30708;
    wire N__30707;
    wire N__30706;
    wire N__30705;
    wire N__30704;
    wire N__30703;
    wire N__30700;
    wire N__30697;
    wire N__30694;
    wire N__30691;
    wire N__30684;
    wire N__30677;
    wire N__30664;
    wire N__30661;
    wire N__30660;
    wire N__30657;
    wire N__30654;
    wire N__30651;
    wire N__30650;
    wire N__30645;
    wire N__30644;
    wire N__30643;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30629;
    wire N__30622;
    wire N__30619;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30611;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30597;
    wire N__30592;
    wire N__30591;
    wire N__30588;
    wire N__30585;
    wire N__30580;
    wire N__30579;
    wire N__30576;
    wire N__30573;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30558;
    wire N__30557;
    wire N__30554;
    wire N__30551;
    wire N__30550;
    wire N__30547;
    wire N__30544;
    wire N__30541;
    wire N__30538;
    wire N__30535;
    wire N__30526;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30514;
    wire N__30513;
    wire N__30510;
    wire N__30505;
    wire N__30502;
    wire N__30499;
    wire N__30498;
    wire N__30495;
    wire N__30494;
    wire N__30491;
    wire N__30488;
    wire N__30485;
    wire N__30478;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30457;
    wire N__30454;
    wire N__30453;
    wire N__30452;
    wire N__30451;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30443;
    wire N__30436;
    wire N__30433;
    wire N__30432;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30409;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30388;
    wire N__30385;
    wire N__30384;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30370;
    wire N__30367;
    wire N__30366;
    wire N__30363;
    wire N__30360;
    wire N__30355;
    wire N__30352;
    wire N__30349;
    wire N__30346;
    wire N__30343;
    wire N__30340;
    wire N__30339;
    wire N__30338;
    wire N__30335;
    wire N__30332;
    wire N__30329;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30301;
    wire N__30300;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30288;
    wire N__30283;
    wire N__30280;
    wire N__30279;
    wire N__30278;
    wire N__30277;
    wire N__30274;
    wire N__30269;
    wire N__30266;
    wire N__30259;
    wire N__30256;
    wire N__30253;
    wire N__30252;
    wire N__30249;
    wire N__30246;
    wire N__30241;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30231;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30219;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30192;
    wire N__30187;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30164;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30142;
    wire N__30133;
    wire N__30130;
    wire N__30129;
    wire N__30126;
    wire N__30123;
    wire N__30120;
    wire N__30115;
    wire N__30112;
    wire N__30111;
    wire N__30108;
    wire N__30105;
    wire N__30102;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30085;
    wire N__30082;
    wire N__30079;
    wire N__30076;
    wire N__30073;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30052;
    wire N__30049;
    wire N__30046;
    wire N__30043;
    wire N__30040;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30030;
    wire N__30029;
    wire N__30026;
    wire N__30025;
    wire N__30022;
    wire N__30019;
    wire N__30016;
    wire N__30011;
    wire N__30004;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29992;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29980;
    wire N__29979;
    wire N__29978;
    wire N__29977;
    wire N__29968;
    wire N__29965;
    wire N__29962;
    wire N__29959;
    wire N__29958;
    wire N__29957;
    wire N__29954;
    wire N__29951;
    wire N__29948;
    wire N__29947;
    wire N__29944;
    wire N__29941;
    wire N__29938;
    wire N__29937;
    wire N__29934;
    wire N__29929;
    wire N__29926;
    wire N__29923;
    wire N__29914;
    wire N__29911;
    wire N__29908;
    wire N__29905;
    wire N__29902;
    wire N__29899;
    wire N__29898;
    wire N__29895;
    wire N__29892;
    wire N__29887;
    wire N__29884;
    wire N__29883;
    wire N__29880;
    wire N__29877;
    wire N__29874;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29860;
    wire N__29857;
    wire N__29854;
    wire N__29853;
    wire N__29852;
    wire N__29851;
    wire N__29850;
    wire N__29847;
    wire N__29844;
    wire N__29837;
    wire N__29830;
    wire N__29829;
    wire N__29826;
    wire N__29825;
    wire N__29824;
    wire N__29821;
    wire N__29816;
    wire N__29813;
    wire N__29806;
    wire N__29805;
    wire N__29804;
    wire N__29801;
    wire N__29796;
    wire N__29791;
    wire N__29788;
    wire N__29785;
    wire N__29782;
    wire N__29781;
    wire N__29780;
    wire N__29777;
    wire N__29772;
    wire N__29767;
    wire N__29766;
    wire N__29765;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29753;
    wire N__29746;
    wire N__29743;
    wire N__29742;
    wire N__29739;
    wire N__29736;
    wire N__29733;
    wire N__29728;
    wire N__29727;
    wire N__29722;
    wire N__29721;
    wire N__29718;
    wire N__29715;
    wire N__29710;
    wire N__29707;
    wire N__29706;
    wire N__29705;
    wire N__29702;
    wire N__29699;
    wire N__29696;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29684;
    wire N__29679;
    wire N__29676;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29664;
    wire N__29661;
    wire N__29660;
    wire N__29659;
    wire N__29656;
    wire N__29655;
    wire N__29652;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29640;
    wire N__29639;
    wire N__29636;
    wire N__29631;
    wire N__29628;
    wire N__29623;
    wire N__29618;
    wire N__29611;
    wire N__29608;
    wire N__29605;
    wire N__29602;
    wire N__29601;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29577;
    wire N__29576;
    wire N__29575;
    wire N__29570;
    wire N__29565;
    wire N__29564;
    wire N__29563;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29537;
    wire N__29530;
    wire N__29529;
    wire N__29524;
    wire N__29521;
    wire N__29520;
    wire N__29517;
    wire N__29514;
    wire N__29509;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29497;
    wire N__29494;
    wire N__29491;
    wire N__29488;
    wire N__29485;
    wire N__29482;
    wire N__29479;
    wire N__29476;
    wire N__29473;
    wire N__29470;
    wire N__29467;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29455;
    wire N__29452;
    wire N__29449;
    wire N__29446;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29424;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29416;
    wire N__29413;
    wire N__29412;
    wire N__29411;
    wire N__29408;
    wire N__29405;
    wire N__29402;
    wire N__29399;
    wire N__29394;
    wire N__29389;
    wire N__29380;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29359;
    wire N__29358;
    wire N__29355;
    wire N__29354;
    wire N__29353;
    wire N__29350;
    wire N__29347;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29327;
    wire N__29320;
    wire N__29317;
    wire N__29314;
    wire N__29311;
    wire N__29308;
    wire N__29305;
    wire N__29302;
    wire N__29299;
    wire N__29296;
    wire N__29293;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29283;
    wire N__29280;
    wire N__29277;
    wire N__29272;
    wire N__29271;
    wire N__29270;
    wire N__29267;
    wire N__29264;
    wire N__29261;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29245;
    wire N__29242;
    wire N__29239;
    wire N__29236;
    wire N__29233;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29221;
    wire N__29218;
    wire N__29215;
    wire N__29212;
    wire N__29209;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29199;
    wire N__29194;
    wire N__29193;
    wire N__29192;
    wire N__29189;
    wire N__29186;
    wire N__29183;
    wire N__29180;
    wire N__29173;
    wire N__29170;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29158;
    wire N__29155;
    wire N__29154;
    wire N__29153;
    wire N__29152;
    wire N__29149;
    wire N__29146;
    wire N__29145;
    wire N__29144;
    wire N__29139;
    wire N__29136;
    wire N__29135;
    wire N__29132;
    wire N__29127;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29108;
    wire N__29103;
    wire N__29100;
    wire N__29089;
    wire N__29088;
    wire N__29085;
    wire N__29082;
    wire N__29079;
    wire N__29074;
    wire N__29071;
    wire N__29070;
    wire N__29069;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29057;
    wire N__29050;
    wire N__29049;
    wire N__29046;
    wire N__29043;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29032;
    wire N__29029;
    wire N__29024;
    wire N__29021;
    wire N__29016;
    wire N__29011;
    wire N__29010;
    wire N__29007;
    wire N__29004;
    wire N__29001;
    wire N__28996;
    wire N__28993;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28983;
    wire N__28980;
    wire N__28977;
    wire N__28974;
    wire N__28969;
    wire N__28966;
    wire N__28965;
    wire N__28962;
    wire N__28959;
    wire N__28958;
    wire N__28955;
    wire N__28954;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28930;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28912;
    wire N__28911;
    wire N__28908;
    wire N__28905;
    wire N__28900;
    wire N__28897;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28889;
    wire N__28888;
    wire N__28885;
    wire N__28882;
    wire N__28877;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28857;
    wire N__28856;
    wire N__28849;
    wire N__28846;
    wire N__28845;
    wire N__28844;
    wire N__28843;
    wire N__28840;
    wire N__28837;
    wire N__28832;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28818;
    wire N__28815;
    wire N__28812;
    wire N__28811;
    wire N__28806;
    wire N__28803;
    wire N__28800;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28782;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28772;
    wire N__28771;
    wire N__28770;
    wire N__28767;
    wire N__28762;
    wire N__28759;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28741;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28728;
    wire N__28723;
    wire N__28722;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28708;
    wire N__28705;
    wire N__28704;
    wire N__28701;
    wire N__28698;
    wire N__28695;
    wire N__28690;
    wire N__28687;
    wire N__28684;
    wire N__28681;
    wire N__28678;
    wire N__28675;
    wire N__28672;
    wire N__28669;
    wire N__28666;
    wire N__28663;
    wire N__28660;
    wire N__28657;
    wire N__28654;
    wire N__28651;
    wire N__28648;
    wire N__28645;
    wire N__28642;
    wire N__28639;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28615;
    wire N__28612;
    wire N__28611;
    wire N__28610;
    wire N__28607;
    wire N__28606;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28591;
    wire N__28582;
    wire N__28579;
    wire N__28576;
    wire N__28573;
    wire N__28570;
    wire N__28567;
    wire N__28566;
    wire N__28563;
    wire N__28558;
    wire N__28555;
    wire N__28552;
    wire N__28549;
    wire N__28546;
    wire N__28543;
    wire N__28540;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28525;
    wire N__28522;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28512;
    wire N__28509;
    wire N__28506;
    wire N__28501;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28488;
    wire N__28487;
    wire N__28482;
    wire N__28481;
    wire N__28478;
    wire N__28475;
    wire N__28474;
    wire N__28471;
    wire N__28470;
    wire N__28467;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28447;
    wire N__28438;
    wire N__28435;
    wire N__28432;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28422;
    wire N__28419;
    wire N__28416;
    wire N__28413;
    wire N__28410;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28393;
    wire N__28392;
    wire N__28391;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28366;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28356;
    wire N__28353;
    wire N__28352;
    wire N__28349;
    wire N__28346;
    wire N__28345;
    wire N__28344;
    wire N__28339;
    wire N__28338;
    wire N__28335;
    wire N__28334;
    wire N__28329;
    wire N__28326;
    wire N__28325;
    wire N__28322;
    wire N__28321;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28311;
    wire N__28308;
    wire N__28305;
    wire N__28302;
    wire N__28299;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28273;
    wire N__28270;
    wire N__28269;
    wire N__28266;
    wire N__28263;
    wire N__28258;
    wire N__28255;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28243;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28218;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28195;
    wire N__28192;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28177;
    wire N__28174;
    wire N__28171;
    wire N__28170;
    wire N__28169;
    wire N__28166;
    wire N__28161;
    wire N__28156;
    wire N__28153;
    wire N__28150;
    wire N__28147;
    wire N__28144;
    wire N__28141;
    wire N__28138;
    wire N__28135;
    wire N__28132;
    wire N__28131;
    wire N__28126;
    wire N__28123;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28111;
    wire N__28110;
    wire N__28107;
    wire N__28104;
    wire N__28099;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28089;
    wire N__28084;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28072;
    wire N__28069;
    wire N__28066;
    wire N__28065;
    wire N__28062;
    wire N__28059;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28035;
    wire N__28032;
    wire N__28029;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28017;
    wire N__28012;
    wire N__28009;
    wire N__28006;
    wire N__28003;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27991;
    wire N__27988;
    wire N__27985;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27973;
    wire N__27972;
    wire N__27971;
    wire N__27966;
    wire N__27963;
    wire N__27958;
    wire N__27957;
    wire N__27954;
    wire N__27951;
    wire N__27946;
    wire N__27945;
    wire N__27942;
    wire N__27939;
    wire N__27934;
    wire N__27933;
    wire N__27930;
    wire N__27927;
    wire N__27924;
    wire N__27919;
    wire N__27918;
    wire N__27915;
    wire N__27912;
    wire N__27907;
    wire N__27906;
    wire N__27903;
    wire N__27900;
    wire N__27895;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27883;
    wire N__27882;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27868;
    wire N__27865;
    wire N__27864;
    wire N__27863;
    wire N__27860;
    wire N__27859;
    wire N__27858;
    wire N__27855;
    wire N__27852;
    wire N__27849;
    wire N__27844;
    wire N__27841;
    wire N__27832;
    wire N__27831;
    wire N__27826;
    wire N__27825;
    wire N__27824;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27795;
    wire N__27790;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27780;
    wire N__27777;
    wire N__27772;
    wire N__27769;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27753;
    wire N__27748;
    wire N__27747;
    wire N__27746;
    wire N__27743;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27729;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27715;
    wire N__27714;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27697;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27685;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27673;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27658;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27646;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27634;
    wire N__27633;
    wire N__27630;
    wire N__27627;
    wire N__27622;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27612;
    wire N__27607;
    wire N__27606;
    wire N__27603;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27593;
    wire N__27590;
    wire N__27583;
    wire N__27580;
    wire N__27579;
    wire N__27578;
    wire N__27575;
    wire N__27574;
    wire N__27569;
    wire N__27566;
    wire N__27563;
    wire N__27560;
    wire N__27555;
    wire N__27552;
    wire N__27549;
    wire N__27546;
    wire N__27543;
    wire N__27538;
    wire N__27535;
    wire N__27532;
    wire N__27531;
    wire N__27530;
    wire N__27527;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27510;
    wire N__27505;
    wire N__27504;
    wire N__27503;
    wire N__27496;
    wire N__27493;
    wire N__27492;
    wire N__27489;
    wire N__27486;
    wire N__27481;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27469;
    wire N__27468;
    wire N__27465;
    wire N__27462;
    wire N__27459;
    wire N__27454;
    wire N__27453;
    wire N__27450;
    wire N__27447;
    wire N__27442;
    wire N__27441;
    wire N__27438;
    wire N__27435;
    wire N__27430;
    wire N__27429;
    wire N__27426;
    wire N__27423;
    wire N__27418;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27403;
    wire N__27402;
    wire N__27399;
    wire N__27396;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27379;
    wire N__27376;
    wire N__27373;
    wire N__27372;
    wire N__27369;
    wire N__27366;
    wire N__27363;
    wire N__27358;
    wire N__27355;
    wire N__27352;
    wire N__27349;
    wire N__27346;
    wire N__27343;
    wire N__27342;
    wire N__27339;
    wire N__27338;
    wire N__27335;
    wire N__27334;
    wire N__27331;
    wire N__27330;
    wire N__27329;
    wire N__27326;
    wire N__27323;
    wire N__27322;
    wire N__27319;
    wire N__27316;
    wire N__27311;
    wire N__27310;
    wire N__27309;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27297;
    wire N__27292;
    wire N__27289;
    wire N__27286;
    wire N__27283;
    wire N__27280;
    wire N__27277;
    wire N__27272;
    wire N__27269;
    wire N__27256;
    wire N__27255;
    wire N__27250;
    wire N__27247;
    wire N__27246;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27232;
    wire N__27229;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27214;
    wire N__27211;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27160;
    wire N__27157;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27133;
    wire N__27130;
    wire N__27127;
    wire N__27124;
    wire N__27123;
    wire N__27120;
    wire N__27115;
    wire N__27112;
    wire N__27109;
    wire N__27108;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27087;
    wire N__27082;
    wire N__27079;
    wire N__27076;
    wire N__27073;
    wire N__27070;
    wire N__27067;
    wire N__27066;
    wire N__27063;
    wire N__27060;
    wire N__27055;
    wire N__27054;
    wire N__27051;
    wire N__27048;
    wire N__27043;
    wire N__27042;
    wire N__27041;
    wire N__27040;
    wire N__27037;
    wire N__27036;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27016;
    wire N__27013;
    wire N__27010;
    wire N__27009;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26997;
    wire N__26992;
    wire N__26989;
    wire N__26988;
    wire N__26987;
    wire N__26984;
    wire N__26979;
    wire N__26978;
    wire N__26975;
    wire N__26972;
    wire N__26971;
    wire N__26970;
    wire N__26967;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26938;
    wire N__26935;
    wire N__26932;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26896;
    wire N__26893;
    wire N__26890;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26875;
    wire N__26874;
    wire N__26873;
    wire N__26870;
    wire N__26867;
    wire N__26866;
    wire N__26865;
    wire N__26864;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26834;
    wire N__26831;
    wire N__26828;
    wire N__26825;
    wire N__26822;
    wire N__26819;
    wire N__26814;
    wire N__26811;
    wire N__26806;
    wire N__26797;
    wire N__26796;
    wire N__26793;
    wire N__26792;
    wire N__26791;
    wire N__26790;
    wire N__26789;
    wire N__26788;
    wire N__26785;
    wire N__26784;
    wire N__26783;
    wire N__26782;
    wire N__26781;
    wire N__26780;
    wire N__26779;
    wire N__26776;
    wire N__26771;
    wire N__26766;
    wire N__26761;
    wire N__26756;
    wire N__26749;
    wire N__26746;
    wire N__26745;
    wire N__26744;
    wire N__26743;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26733;
    wire N__26730;
    wire N__26723;
    wire N__26720;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26704;
    wire N__26701;
    wire N__26696;
    wire N__26683;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26673;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26659;
    wire N__26658;
    wire N__26655;
    wire N__26652;
    wire N__26649;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26632;
    wire N__26629;
    wire N__26626;
    wire N__26623;
    wire N__26622;
    wire N__26619;
    wire N__26616;
    wire N__26613;
    wire N__26608;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26571;
    wire N__26568;
    wire N__26565;
    wire N__26562;
    wire N__26557;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26541;
    wire N__26538;
    wire N__26535;
    wire N__26532;
    wire N__26527;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26517;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26500;
    wire N__26497;
    wire N__26494;
    wire N__26493;
    wire N__26490;
    wire N__26487;
    wire N__26482;
    wire N__26481;
    wire N__26478;
    wire N__26475;
    wire N__26472;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26460;
    wire N__26457;
    wire N__26454;
    wire N__26451;
    wire N__26446;
    wire N__26443;
    wire N__26440;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26427;
    wire N__26424;
    wire N__26423;
    wire N__26420;
    wire N__26419;
    wire N__26418;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26408;
    wire N__26403;
    wire N__26400;
    wire N__26397;
    wire N__26394;
    wire N__26389;
    wire N__26380;
    wire N__26379;
    wire N__26374;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26350;
    wire N__26347;
    wire N__26344;
    wire N__26341;
    wire N__26338;
    wire N__26335;
    wire N__26334;
    wire N__26329;
    wire N__26326;
    wire N__26325;
    wire N__26324;
    wire N__26321;
    wire N__26320;
    wire N__26315;
    wire N__26312;
    wire N__26311;
    wire N__26310;
    wire N__26307;
    wire N__26304;
    wire N__26301;
    wire N__26298;
    wire N__26295;
    wire N__26292;
    wire N__26289;
    wire N__26278;
    wire N__26275;
    wire N__26274;
    wire N__26269;
    wire N__26266;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26239;
    wire N__26238;
    wire N__26233;
    wire N__26230;
    wire N__26227;
    wire N__26224;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26212;
    wire N__26211;
    wire N__26208;
    wire N__26205;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26182;
    wire N__26179;
    wire N__26176;
    wire N__26173;
    wire N__26170;
    wire N__26167;
    wire N__26164;
    wire N__26161;
    wire N__26158;
    wire N__26155;
    wire N__26152;
    wire N__26149;
    wire N__26148;
    wire N__26145;
    wire N__26142;
    wire N__26137;
    wire N__26134;
    wire N__26131;
    wire N__26128;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26116;
    wire N__26113;
    wire N__26110;
    wire N__26107;
    wire N__26104;
    wire N__26101;
    wire N__26098;
    wire N__26095;
    wire N__26092;
    wire N__26089;
    wire N__26086;
    wire N__26085;
    wire N__26082;
    wire N__26079;
    wire N__26076;
    wire N__26071;
    wire N__26070;
    wire N__26067;
    wire N__26064;
    wire N__26059;
    wire N__26058;
    wire N__26055;
    wire N__26052;
    wire N__26049;
    wire N__26044;
    wire N__26043;
    wire N__26040;
    wire N__26037;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26020;
    wire N__26017;
    wire N__26016;
    wire N__26013;
    wire N__26010;
    wire N__26005;
    wire N__26004;
    wire N__26001;
    wire N__25998;
    wire N__25993;
    wire N__25992;
    wire N__25991;
    wire N__25988;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25974;
    wire N__25971;
    wire N__25966;
    wire N__25965;
    wire N__25960;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25929;
    wire N__25924;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25905;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25888;
    wire N__25885;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25873;
    wire N__25870;
    wire N__25867;
    wire N__25864;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25840;
    wire N__25837;
    wire N__25834;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25810;
    wire N__25807;
    wire N__25804;
    wire N__25803;
    wire N__25800;
    wire N__25797;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25780;
    wire N__25777;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25741;
    wire N__25738;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25711;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25684;
    wire N__25681;
    wire N__25678;
    wire N__25675;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25660;
    wire N__25657;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25638;
    wire N__25637;
    wire N__25636;
    wire N__25635;
    wire N__25634;
    wire N__25633;
    wire N__25630;
    wire N__25627;
    wire N__25626;
    wire N__25623;
    wire N__25620;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25607;
    wire N__25604;
    wire N__25601;
    wire N__25596;
    wire N__25591;
    wire N__25590;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25570;
    wire N__25565;
    wire N__25558;
    wire N__25549;
    wire N__25546;
    wire N__25543;
    wire N__25540;
    wire N__25539;
    wire N__25536;
    wire N__25531;
    wire N__25528;
    wire N__25525;
    wire N__25522;
    wire N__25521;
    wire N__25518;
    wire N__25515;
    wire N__25512;
    wire N__25507;
    wire N__25504;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25482;
    wire N__25479;
    wire N__25476;
    wire N__25471;
    wire N__25468;
    wire N__25465;
    wire N__25462;
    wire N__25459;
    wire N__25458;
    wire N__25453;
    wire N__25450;
    wire N__25449;
    wire N__25444;
    wire N__25441;
    wire N__25438;
    wire N__25435;
    wire N__25432;
    wire N__25429;
    wire N__25426;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25411;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25399;
    wire N__25398;
    wire N__25393;
    wire N__25390;
    wire N__25387;
    wire N__25384;
    wire N__25381;
    wire N__25378;
    wire N__25375;
    wire N__25372;
    wire N__25369;
    wire N__25366;
    wire N__25363;
    wire N__25360;
    wire N__25357;
    wire N__25354;
    wire N__25351;
    wire N__25348;
    wire N__25345;
    wire N__25342;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25330;
    wire N__25327;
    wire N__25324;
    wire N__25321;
    wire N__25320;
    wire N__25319;
    wire N__25318;
    wire N__25317;
    wire N__25316;
    wire N__25315;
    wire N__25314;
    wire N__25313;
    wire N__25312;
    wire N__25311;
    wire N__25310;
    wire N__25309;
    wire N__25308;
    wire N__25307;
    wire N__25306;
    wire N__25303;
    wire N__25302;
    wire N__25299;
    wire N__25298;
    wire N__25295;
    wire N__25294;
    wire N__25293;
    wire N__25290;
    wire N__25289;
    wire N__25286;
    wire N__25285;
    wire N__25282;
    wire N__25281;
    wire N__25278;
    wire N__25275;
    wire N__25274;
    wire N__25271;
    wire N__25270;
    wire N__25267;
    wire N__25266;
    wire N__25263;
    wire N__25262;
    wire N__25261;
    wire N__25258;
    wire N__25255;
    wire N__25252;
    wire N__25251;
    wire N__25250;
    wire N__25247;
    wire N__25246;
    wire N__25243;
    wire N__25230;
    wire N__25213;
    wire N__25196;
    wire N__25187;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25179;
    wire N__25174;
    wire N__25165;
    wire N__25162;
    wire N__25153;
    wire N__25150;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25108;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25075;
    wire N__25072;
    wire N__25069;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25045;
    wire N__25042;
    wire N__25039;
    wire N__25036;
    wire N__25033;
    wire N__25030;
    wire N__25027;
    wire N__25026;
    wire N__25025;
    wire N__25022;
    wire N__25021;
    wire N__25018;
    wire N__25011;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24997;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24976;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24961;
    wire N__24958;
    wire N__24955;
    wire N__24954;
    wire N__24953;
    wire N__24950;
    wire N__24947;
    wire N__24942;
    wire N__24939;
    wire N__24938;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24926;
    wire N__24919;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24911;
    wire N__24906;
    wire N__24903;
    wire N__24898;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24888;
    wire N__24887;
    wire N__24884;
    wire N__24881;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24859;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24844;
    wire N__24841;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24829;
    wire N__24826;
    wire N__24823;
    wire N__24820;
    wire N__24819;
    wire N__24816;
    wire N__24813;
    wire N__24808;
    wire N__24805;
    wire N__24802;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24790;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24769;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24757;
    wire N__24754;
    wire N__24751;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24736;
    wire N__24733;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24721;
    wire N__24718;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24703;
    wire N__24700;
    wire N__24699;
    wire N__24696;
    wire N__24693;
    wire N__24688;
    wire N__24685;
    wire N__24682;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24667;
    wire N__24664;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24639;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24625;
    wire N__24622;
    wire N__24621;
    wire N__24618;
    wire N__24615;
    wire N__24612;
    wire N__24607;
    wire N__24604;
    wire N__24601;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24589;
    wire N__24586;
    wire N__24583;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24562;
    wire N__24559;
    wire N__24556;
    wire N__24553;
    wire N__24552;
    wire N__24547;
    wire N__24544;
    wire N__24541;
    wire N__24538;
    wire N__24535;
    wire N__24532;
    wire N__24529;
    wire N__24526;
    wire N__24523;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24499;
    wire N__24498;
    wire N__24493;
    wire N__24490;
    wire N__24489;
    wire N__24486;
    wire N__24483;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24457;
    wire N__24454;
    wire N__24451;
    wire N__24448;
    wire N__24445;
    wire N__24442;
    wire N__24439;
    wire N__24436;
    wire N__24433;
    wire N__24430;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24403;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24334;
    wire N__24331;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24316;
    wire N__24315;
    wire N__24312;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24299;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24283;
    wire N__24282;
    wire N__24279;
    wire N__24278;
    wire N__24275;
    wire N__24272;
    wire N__24271;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24259;
    wire N__24250;
    wire N__24247;
    wire N__24244;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24224;
    wire N__24217;
    wire N__24214;
    wire N__24213;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24201;
    wire N__24198;
    wire N__24195;
    wire N__24192;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24180;
    wire N__24177;
    wire N__24174;
    wire N__24171;
    wire N__24166;
    wire N__24163;
    wire N__24160;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24150;
    wire N__24145;
    wire N__24142;
    wire N__24141;
    wire N__24138;
    wire N__24135;
    wire N__24132;
    wire N__24127;
    wire N__24124;
    wire N__24123;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24109;
    wire N__24106;
    wire N__24103;
    wire N__24102;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24088;
    wire N__24085;
    wire N__24082;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24067;
    wire N__24064;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24049;
    wire N__24046;
    wire N__24043;
    wire N__24042;
    wire N__24041;
    wire N__24038;
    wire N__24033;
    wire N__24028;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24012;
    wire N__24009;
    wire N__24006;
    wire N__24003;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23989;
    wire N__23988;
    wire N__23985;
    wire N__23982;
    wire N__23979;
    wire N__23974;
    wire N__23971;
    wire N__23970;
    wire N__23967;
    wire N__23964;
    wire N__23961;
    wire N__23956;
    wire N__23953;
    wire N__23950;
    wire N__23949;
    wire N__23946;
    wire N__23943;
    wire N__23940;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23919;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23907;
    wire N__23904;
    wire N__23901;
    wire N__23898;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23878;
    wire N__23875;
    wire N__23872;
    wire N__23871;
    wire N__23868;
    wire N__23865;
    wire N__23860;
    wire N__23857;
    wire N__23854;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23799;
    wire N__23798;
    wire N__23795;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23779;
    wire N__23778;
    wire N__23773;
    wire N__23772;
    wire N__23771;
    wire N__23768;
    wire N__23763;
    wire N__23760;
    wire N__23757;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23743;
    wire N__23740;
    wire N__23737;
    wire N__23734;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23722;
    wire N__23719;
    wire N__23716;
    wire N__23713;
    wire N__23710;
    wire N__23707;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23695;
    wire N__23692;
    wire N__23689;
    wire N__23686;
    wire N__23683;
    wire N__23680;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire VCCG0;
    wire CLK_c;
    wire tx_enable;
    wire GB_BUFFER_PIN_9_c_THRU_CO;
    wire LED_c;
    wire \quad_counter1.n26_adj_4207_cascade_ ;
    wire \quad_counter1.n25_adj_4209 ;
    wire n12907;
    wire quadB_delayed_adj_4543;
    wire PIN_13_c;
    wire n12907_cascade_;
    wire \quad_counter1.n27_adj_4208 ;
    wire \quad_counter1.n28_adj_4206 ;
    wire bfn_7_17_0_;
    wire \c0.n19612 ;
    wire \c0.n19613 ;
    wire \c0.n19614 ;
    wire \c0.n19615 ;
    wire \c0.n19616 ;
    wire \c0.n19617 ;
    wire \c0.n19618 ;
    wire n23768_cascade_;
    wire n23897_cascade_;
    wire n10_adj_4532_cascade_;
    wire \c0.n21322 ;
    wire rx_i;
    wire \quad_counter1.n27 ;
    wire \quad_counter1.n28_cascade_ ;
    wire \quad_counter1.n25 ;
    wire n9818_cascade_;
    wire b_delay_counter_0_adj_4541;
    wire n187_adj_4546;
    wire bfn_9_10_0_;
    wire \quad_counter1.b_delay_counter_1 ;
    wire \quad_counter1.n19503 ;
    wire \quad_counter1.b_delay_counter_2 ;
    wire \quad_counter1.n19504 ;
    wire \quad_counter1.b_delay_counter_3 ;
    wire \quad_counter1.n19505 ;
    wire \quad_counter1.b_delay_counter_4 ;
    wire \quad_counter1.n19506 ;
    wire \quad_counter1.b_delay_counter_5 ;
    wire \quad_counter1.n19507 ;
    wire \quad_counter1.b_delay_counter_6 ;
    wire \quad_counter1.n19508 ;
    wire \quad_counter1.b_delay_counter_7 ;
    wire \quad_counter1.n19509 ;
    wire \quad_counter1.n19510 ;
    wire \quad_counter1.b_delay_counter_8 ;
    wire bfn_9_11_0_;
    wire \quad_counter1.b_delay_counter_9 ;
    wire \quad_counter1.n19511 ;
    wire \quad_counter1.b_delay_counter_10 ;
    wire \quad_counter1.n19512 ;
    wire \quad_counter1.b_delay_counter_11 ;
    wire \quad_counter1.n19513 ;
    wire \quad_counter1.b_delay_counter_12 ;
    wire \quad_counter1.n19514 ;
    wire \quad_counter1.b_delay_counter_13 ;
    wire \quad_counter1.n19515 ;
    wire \quad_counter1.b_delay_counter_14 ;
    wire \quad_counter1.n19516 ;
    wire \quad_counter1.n19517 ;
    wire \quad_counter1.b_delay_counter_15 ;
    wire n14377;
    wire b_delay_counter_15__N_4141_adj_4548;
    wire \quad_counter1.A_delayed ;
    wire B_filtered_adj_4539;
    wire count_enable_adj_4544_cascade_;
    wire data_out_frame_10_6;
    wire n26;
    wire n24118_cascade_;
    wire \c0.n23950_cascade_ ;
    wire \c0.n24147_cascade_ ;
    wire \c0.n23882 ;
    wire n24150;
    wire n24097_cascade_;
    wire n24117;
    wire n24112;
    wire n23849_cascade_;
    wire data_out_frame_10_3;
    wire \c0.n24159_cascade_ ;
    wire \c0.n24162 ;
    wire \c0.n11_adj_4355 ;
    wire n23846;
    wire n24114_cascade_;
    wire n10;
    wire \c0.n23895 ;
    wire \c0.n24051_cascade_ ;
    wire \c0.n23844 ;
    wire \c0.n23847 ;
    wire \c0.n11_adj_4348 ;
    wire n24102;
    wire \c0.n24047 ;
    wire \c0.n5_adj_4358 ;
    wire data_out_frame_6_7;
    wire data_out_frame_0_3;
    wire \c0.n24011 ;
    wire data_out_frame_0_2;
    wire \c0.n6_adj_4521 ;
    wire \c0.n23859_cascade_ ;
    wire n23861_cascade_;
    wire n10_adj_4534;
    wire \c0.n5_adj_4522 ;
    wire data_out_frame_6_2;
    wire \c0.n24007 ;
    wire \c0.n6 ;
    wire r_Tx_Data_6;
    wire r_Tx_Data_2;
    wire b_delay_counter_15__N_4141_cascade_;
    wire bfn_10_9_0_;
    wire \quad_counter1.a_delay_counter_1 ;
    wire \quad_counter1.n19518 ;
    wire \quad_counter1.a_delay_counter_2 ;
    wire \quad_counter1.n19519 ;
    wire \quad_counter1.a_delay_counter_3 ;
    wire \quad_counter1.n19520 ;
    wire \quad_counter1.a_delay_counter_4 ;
    wire \quad_counter1.n19521 ;
    wire \quad_counter1.a_delay_counter_5 ;
    wire \quad_counter1.n19522 ;
    wire \quad_counter1.n19523 ;
    wire \quad_counter1.a_delay_counter_7 ;
    wire \quad_counter1.n19524 ;
    wire \quad_counter1.n19525 ;
    wire \quad_counter1.a_delay_counter_8 ;
    wire bfn_10_10_0_;
    wire \quad_counter1.n19526 ;
    wire \quad_counter1.a_delay_counter_10 ;
    wire \quad_counter1.n19527 ;
    wire \quad_counter1.a_delay_counter_11 ;
    wire \quad_counter1.n19528 ;
    wire \quad_counter1.n19529 ;
    wire \quad_counter1.n19530 ;
    wire \quad_counter1.a_delay_counter_14 ;
    wire \quad_counter1.n19531 ;
    wire \quad_counter1.n19532 ;
    wire \quad_counter1.a_delay_counter_15 ;
    wire data_out_frame_11_6;
    wire A_filtered_adj_4538;
    wire \quad_counter1.B_delayed ;
    wire n39_adj_4545;
    wire a_delay_counter_0_adj_4540;
    wire \c0.n22048_cascade_ ;
    wire bfn_10_13_0_;
    wire encoder1_position_0;
    wire \quad_counter1.count_direction ;
    wire n2205;
    wire \quad_counter1.n19548 ;
    wire \quad_counter1.n19549 ;
    wire n2203;
    wire \quad_counter1.n19550 ;
    wire n2202;
    wire \quad_counter1.n19551 ;
    wire \quad_counter1.n19552 ;
    wire n2200;
    wire \quad_counter1.n19553 ;
    wire n2199;
    wire \quad_counter1.n19554 ;
    wire \quad_counter1.n19555 ;
    wire bfn_10_14_0_;
    wire \quad_counter1.n19556 ;
    wire \quad_counter1.n19557 ;
    wire \quad_counter1.n19558 ;
    wire \quad_counter1.n19559 ;
    wire \quad_counter1.n19560 ;
    wire \quad_counter1.n19561 ;
    wire n2191;
    wire \quad_counter1.n19562 ;
    wire \quad_counter1.n19563 ;
    wire n2190;
    wire bfn_10_15_0_;
    wire \quad_counter1.n19564 ;
    wire \quad_counter1.n19565 ;
    wire n2187;
    wire \quad_counter1.n19566 ;
    wire \quad_counter1.n19567 ;
    wire \quad_counter1.n19568 ;
    wire \quad_counter1.n19569 ;
    wire n2183;
    wire \quad_counter1.n19570 ;
    wire \quad_counter1.n19571 ;
    wire bfn_10_16_0_;
    wire \quad_counter1.n19572 ;
    wire \quad_counter1.n19573 ;
    wire n2179;
    wire \quad_counter1.n19574 ;
    wire \quad_counter1.n19575 ;
    wire n2177;
    wire \quad_counter1.n19576 ;
    wire \quad_counter1.n19577 ;
    wire \quad_counter1.n19578 ;
    wire \quad_counter1.n19579 ;
    wire \quad_counter1.n2140 ;
    wire bfn_10_17_0_;
    wire n2174;
    wire data_out_frame_0_4;
    wire data_out_frame_13_5;
    wire data_out_frame_9_3;
    wire \c0.n24171 ;
    wire \c0.n24174 ;
    wire \c0.n23856 ;
    wire n24108;
    wire n23858_cascade_;
    wire r_Tx_Data_5;
    wire r_Tx_Data_4;
    wire n10_adj_4533;
    wire data_out_frame_9_2;
    wire \c0.n24180_cascade_ ;
    wire n24106;
    wire data_out_frame_7_0;
    wire data_out_frame_6_0;
    wire n10_adj_4536;
    wire \c0.n5_adj_4422 ;
    wire \c0.n24059 ;
    wire \c0.n23850_cascade_ ;
    wire n23852_cascade_;
    wire byte_transmit_counter_3;
    wire n10_adj_4537_cascade_;
    wire n24110;
    wire r_Tx_Data_0;
    wire n24195;
    wire n24100_cascade_;
    wire n16706;
    wire \c0.tx.n23985_cascade_ ;
    wire \c0.tx.n31_adj_4216_cascade_ ;
    wire n187;
    wire bfn_10_22_0_;
    wire \quad_counter0.n19473 ;
    wire \quad_counter0.n19474 ;
    wire \quad_counter0.n19475 ;
    wire \quad_counter0.n19476 ;
    wire \quad_counter0.n19477 ;
    wire \quad_counter0.n19478 ;
    wire \quad_counter0.n19479 ;
    wire \quad_counter0.n19480 ;
    wire bfn_10_23_0_;
    wire \quad_counter0.n19481 ;
    wire \quad_counter0.n19482 ;
    wire \quad_counter0.n19483 ;
    wire \quad_counter0.n19484 ;
    wire \quad_counter0.n19485 ;
    wire \quad_counter0.n19486 ;
    wire \quad_counter0.n19487 ;
    wire n14198;
    wire b_delay_counter_15__N_4141;
    wire bfn_10_24_0_;
    wire \quad_counter0.n19488 ;
    wire \quad_counter0.n19489 ;
    wire \quad_counter0.n19490 ;
    wire \quad_counter0.n19491 ;
    wire \quad_counter0.n19492 ;
    wire \quad_counter0.n19493 ;
    wire \quad_counter0.n19494 ;
    wire \quad_counter0.n19495 ;
    wire bfn_10_25_0_;
    wire \quad_counter0.n19496 ;
    wire \quad_counter0.n19497 ;
    wire \quad_counter0.n19498 ;
    wire \quad_counter0.n19499 ;
    wire \quad_counter0.n19500 ;
    wire \quad_counter0.n19501 ;
    wire \quad_counter0.n19502 ;
    wire \c0.n24_adj_4502 ;
    wire \c0.n18_adj_4414_cascade_ ;
    wire \c0.n13360 ;
    wire \c0.n23550_cascade_ ;
    wire \c0.n22_adj_4503_cascade_ ;
    wire \c0.n26_adj_4504 ;
    wire \c0.n26_adj_4517 ;
    wire \c0.n21305_cascade_ ;
    wire \c0.data_out_frame_28_2 ;
    wire \c0.n6_adj_4515 ;
    wire \c0.n12532_cascade_ ;
    wire \c0.n22126_cascade_ ;
    wire \c0.data_out_frame_28_4 ;
    wire \quad_counter1.a_delay_counter_12 ;
    wire \quad_counter1.a_delay_counter_13 ;
    wire \quad_counter1.a_delay_counter_9 ;
    wire \quad_counter1.a_delay_counter_6 ;
    wire \quad_counter1.n26 ;
    wire a_delay_counter_15__N_4124_adj_4547;
    wire quadA_delayed_adj_4542;
    wire PIN_12_c;
    wire a_delay_counter_15__N_4124_adj_4547_cascade_;
    wire n9818;
    wire n14228;
    wire data_out_frame_29_2;
    wire n2196;
    wire \c0.n13079_cascade_ ;
    wire \c0.n22116 ;
    wire \c0.n6_adj_4308 ;
    wire data_out_frame_13_0;
    wire \c0.n11_adj_4424 ;
    wire \c0.n6_adj_4335_cascade_ ;
    wire \c0.n21229_cascade_ ;
    wire n2193;
    wire \c0.n6_adj_4309 ;
    wire n2204;
    wire \c0.n6_adj_4310_cascade_ ;
    wire \c0.n22037 ;
    wire encoder1_position_15;
    wire data_out_frame_12_7;
    wire \c0.n11_adj_4360 ;
    wire n2197;
    wire \c0.n5_adj_4227 ;
    wire data_out_frame_7_4;
    wire \c0.data_out_frame_29__7__N_850 ;
    wire data_out_frame_11_4;
    wire \c0.n23881 ;
    wire n2189;
    wire encoder1_position_16;
    wire data_out_frame_10_4;
    wire data_out_frame_7_2;
    wire n2188;
    wire n2184;
    wire n2182;
    wire n2176;
    wire data_out_frame_29_3;
    wire data_out_frame_28_3;
    wire \c0.n26 ;
    wire n2175;
    wire data_out_frame_7_5;
    wire \c0.n5_adj_4346 ;
    wire data_out_frame_9_7;
    wire tx_o;
    wire \c0.n6_adj_4392 ;
    wire \c0.byte_transmit_counter_6 ;
    wire \c0.n23574_cascade_ ;
    wire \c0.byte_transmit_counter_7 ;
    wire \c0.n38_adj_4387_cascade_ ;
    wire data_out_frame_5_2;
    wire n23768;
    wire byte_transmit_counter_4;
    wire n23864;
    wire data_out_frame_5_6;
    wire data_out_frame_13_3;
    wire \c0.n11_adj_4218 ;
    wire data_out_frame_11_5;
    wire data_out_frame_9_5;
    wire \c0.n24141_cascade_ ;
    wire data_out_frame_8_5;
    wire \c0.n24144 ;
    wire r_Tx_Data_7;
    wire r_Tx_Data_3;
    wire r_Bit_Index_2_adj_4551;
    wire n4_adj_4554;
    wire n24189_cascade_;
    wire r_Bit_Index_1_adj_4552;
    wire n10_adj_4535;
    wire byte_transmit_counter_5;
    wire r_Tx_Data_1;
    wire data_in_0_7;
    wire data_out_frame_5_3;
    wire data_out_frame_6_3;
    wire \c0.n5 ;
    wire data_out_frame_5_5;
    wire data_out_frame_11_0;
    wire \c0.n24165_cascade_ ;
    wire \c0.n24168 ;
    wire \quad_counter0.b_delay_counter_3 ;
    wire \quad_counter0.b_delay_counter_9 ;
    wire \quad_counter0.b_delay_counter_4 ;
    wire b_delay_counter_0;
    wire PIN_8_c;
    wire quadB_delayed;
    wire B_filtered;
    wire \quad_counter0.b_delay_counter_13 ;
    wire \quad_counter0.b_delay_counter_1 ;
    wire \quad_counter0.b_delay_counter_2 ;
    wire \quad_counter0.b_delay_counter_5 ;
    wire \quad_counter0.b_delay_counter_11 ;
    wire \quad_counter0.b_delay_counter_10 ;
    wire \quad_counter0.b_delay_counter_8 ;
    wire \quad_counter0.b_delay_counter_6 ;
    wire \quad_counter0.n28_adj_4198 ;
    wire \quad_counter0.n26_adj_4199_cascade_ ;
    wire \quad_counter0.n25_adj_4201 ;
    wire n12909;
    wire \quad_counter0.A_delayed ;
    wire \quad_counter0.B_delayed ;
    wire \quad_counter0.a_delay_counter_3 ;
    wire \quad_counter0.a_delay_counter_8 ;
    wire \quad_counter0.a_delay_counter_2 ;
    wire \quad_counter0.a_delay_counter_1 ;
    wire \quad_counter0.a_delay_counter_5 ;
    wire \quad_counter0.a_delay_counter_11 ;
    wire \quad_counter0.a_delay_counter_4 ;
    wire A_filtered;
    wire PIN_7_c;
    wire quadA_delayed;
    wire n14421;
    wire a_delay_counter_15__N_4124;
    wire n39;
    wire n14421_cascade_;
    wire a_delay_counter_0;
    wire \quad_counter0.a_delay_counter_14 ;
    wire \quad_counter0.a_delay_counter_15 ;
    wire \quad_counter0.a_delay_counter_7 ;
    wire \quad_counter0.a_delay_counter_10 ;
    wire \quad_counter0.n28_adj_4202 ;
    wire \quad_counter0.n27_adj_4204_cascade_ ;
    wire \quad_counter0.n25_adj_4205 ;
    wire n9821;
    wire \quad_counter0.a_delay_counter_12 ;
    wire \quad_counter0.a_delay_counter_13 ;
    wire \quad_counter0.a_delay_counter_6 ;
    wire \quad_counter0.a_delay_counter_9 ;
    wire \quad_counter0.n26_adj_4203 ;
    wire data_out_frame_28__3__N_1881;
    wire \c0.n20257 ;
    wire \c0.n21062 ;
    wire \c0.data_out_frame_28_1 ;
    wire \c0.data_out_frame_29_1 ;
    wire \c0.n26_adj_4519 ;
    wire \c0.n12542_cascade_ ;
    wire \c0.n14_adj_4340_cascade_ ;
    wire \c0.n20320 ;
    wire \c0.n20320_cascade_ ;
    wire \c0.n22180_cascade_ ;
    wire \c0.n10498_cascade_ ;
    wire \c0.n20253_cascade_ ;
    wire \c0.n21229 ;
    wire \c0.n15_adj_4513 ;
    wire \c0.n22066 ;
    wire encoder1_position_3;
    wire \c0.n21071_cascade_ ;
    wire data_out_frame_29__2__N_1749;
    wire \c0.n17_adj_4501 ;
    wire \c0.data_out_frame_29_0 ;
    wire \c0.n26_adj_4423 ;
    wire \c0.n16_adj_4500 ;
    wire \c0.n10422 ;
    wire \c0.n6_adj_4313_cascade_ ;
    wire \c0.n21156_cascade_ ;
    wire \c0.n21175_cascade_ ;
    wire \c0.n20276_cascade_ ;
    wire \c0.n21110_cascade_ ;
    wire \c0.n14_adj_4514 ;
    wire encoder1_position_22;
    wire n2201;
    wire \c0.n22277 ;
    wire \c0.n22102_cascade_ ;
    wire \c0.n22293 ;
    wire \c0.n15_adj_4325_cascade_ ;
    wire \c0.n21041 ;
    wire \c0.n21041_cascade_ ;
    wire \c0.n22102 ;
    wire \c0.n22361_cascade_ ;
    wire \c0.n10_adj_4314 ;
    wire encoder1_position_21;
    wire \c0.n24153 ;
    wire data_out_frame_8_6;
    wire \c0.n24156 ;
    wire data_out_frame_12_6;
    wire data_out_frame_11_3;
    wire n2181;
    wire \c0.n22224 ;
    wire \c0.n22224_cascade_ ;
    wire \c0.n13349_cascade_ ;
    wire \c0.n6_adj_4334 ;
    wire n24104;
    wire \c0.n22405 ;
    wire encoder1_position_31;
    wire data_out_frame_10_7;
    wire data_out_frame_8_7;
    wire data_out_frame_11_7;
    wire data_out_frame_12_3;
    wire \c0.n7_adj_4492_cascade_ ;
    wire data_in_1_5;
    wire \c0.n9_adj_4493 ;
    wire \c0.n23600 ;
    wire data_in_0_6;
    wire data_in_2_2;
    wire data_in_0_3;
    wire \c0.n14_adj_4495_cascade_ ;
    wire \c0.n15_adj_4496 ;
    wire \c0.n10_adj_4231_cascade_ ;
    wire \c0.n14 ;
    wire n9539;
    wire data_out_frame_10_0;
    wire data_in_3_3;
    wire encoder1_position_18;
    wire data_out_frame_11_2;
    wire \c0.n24177 ;
    wire data_out_frame_5_0;
    wire encoder1_position_29;
    wire data_out_frame_10_5;
    wire \c0.tx.n16631_cascade_ ;
    wire n14442;
    wire \c0.n21370 ;
    wire \c0.n21376 ;
    wire \c0.n21362 ;
    wire \c0.n21128 ;
    wire \c0.n12_adj_4516 ;
    wire \c0.n9_adj_4339 ;
    wire \c0.n22018_cascade_ ;
    wire \c0.n21946 ;
    wire \c0.n21946_cascade_ ;
    wire \c0.n12532 ;
    wire \c0.n12491_cascade_ ;
    wire \c0.data_out_frame_28_6 ;
    wire \c0.n26_adj_4351 ;
    wire \c0.n7_adj_4307_cascade_ ;
    wire data_out_frame_29__3__N_1662;
    wire \c0.n22024 ;
    wire \c0.data_out_frame_29_4 ;
    wire \c0.n22151 ;
    wire \c0.n22151_cascade_ ;
    wire \c0.n6_adj_4397_cascade_ ;
    wire \c0.data_out_frame_28_0 ;
    wire \c0.n22018 ;
    wire \c0.data_out_frame_29_5 ;
    wire \c0.data_out_frame_28_5 ;
    wire \c0.n26_adj_4347 ;
    wire \c0.n20376 ;
    wire \c0.n6_adj_4509_cascade_ ;
    wire \c0.n22393 ;
    wire \c0.n10498 ;
    wire \c0.n22393_cascade_ ;
    wire \c0.n14_adj_4510_cascade_ ;
    wire \c0.n10462 ;
    wire \c0.n21150 ;
    wire \c0.n10_adj_4511 ;
    wire \c0.n10_adj_4330 ;
    wire \c0.n21192_cascade_ ;
    wire \c0.n20931_cascade_ ;
    wire \c0.n21175 ;
    wire \c0.n21156 ;
    wire \c0.n12554 ;
    wire \c0.n20931 ;
    wire \c0.n22991 ;
    wire \c0.n21189_cascade_ ;
    wire \c0.n21058 ;
    wire \c0.n21192 ;
    wire \c0.n13349 ;
    wire \c0.n13480_cascade_ ;
    wire \c0.n21122_cascade_ ;
    wire encoder1_position_14;
    wire \c0.n20767 ;
    wire \c0.n20767_cascade_ ;
    wire encoder1_position_24;
    wire n2195;
    wire data_out_frame_9_6;
    wire data_out_frame_13_6;
    wire n2194;
    wire \c0.n11 ;
    wire \c0.n14_adj_4329 ;
    wire n2198;
    wire n2192;
    wire n2186;
    wire encoder1_position_19;
    wire \c0.n19_adj_4319 ;
    wire \c0.n23557 ;
    wire n2180;
    wire \c0.n21914_cascade_ ;
    wire \c0.n21_adj_4320 ;
    wire data_out_frame_8_4;
    wire \c0.n23880 ;
    wire data_out_frame_9_4;
    wire n2178;
    wire encoder1_position_27;
    wire data_out_frame_10_2;
    wire data_out_frame_5_4;
    wire data_out_frame_6_4;
    wire \c0.n13003 ;
    wire \c0.n19_adj_4367 ;
    wire \c0.n20_adj_4362_cascade_ ;
    wire \c0.n23834 ;
    wire data_in_1_2;
    wire data_in_0_5;
    wire data_in_1_6;
    wire \c0.n17_adj_4479_cascade_ ;
    wire \c0.n13023 ;
    wire data_in_0_2;
    wire \c0.n13006 ;
    wire \c0.n21767 ;
    wire \c0.tx.n14296 ;
    wire data_in_1_0;
    wire data_in_0_0;
    wire data_in_0_4;
    wire data_in_1_7;
    wire \c0.n10_adj_4494 ;
    wire \c0.n16_adj_4476 ;
    wire \c0.n17_adj_4477 ;
    wire r_Bit_Index_0_adj_4553;
    wire n24192;
    wire n24198;
    wire o_Tx_Serial_N_3783_cascade_;
    wire \c0.tx.n12 ;
    wire r_SM_Main_1_adj_4550;
    wire \c0.tx.n6_adj_4214_cascade_ ;
    wire \c0.tx.n16630 ;
    wire n8_cascade_;
    wire \c0.tx.n6_cascade_ ;
    wire \c0.tx.n31 ;
    wire \c0.tx.n31_cascade_ ;
    wire \c0.tx.n47 ;
    wire \c0.tx.n10 ;
    wire \c0.tx.r_Clock_Count_0 ;
    wire \c0.tx.n23960 ;
    wire bfn_13_21_0_;
    wire \c0.tx.r_Clock_Count_1 ;
    wire \c0.tx.n23961 ;
    wire \c0.tx.n19540 ;
    wire \c0.tx.r_Clock_Count_2 ;
    wire \c0.tx.n23958 ;
    wire \c0.tx.n19541 ;
    wire \c0.tx.r_Clock_Count_3 ;
    wire \c0.tx.n23963 ;
    wire \c0.tx.n19542 ;
    wire \c0.tx.r_Clock_Count_4 ;
    wire \c0.tx.n23953 ;
    wire \c0.tx.n19543 ;
    wire r_Clock_Count_5;
    wire n316;
    wire \c0.tx.n19544 ;
    wire \c0.tx.n19545 ;
    wire r_Clock_Count_7;
    wire n314;
    wire \c0.tx.n19546 ;
    wire \c0.tx.n19547 ;
    wire bfn_13_22_0_;
    wire \c0.n12878 ;
    wire \c0.n21360 ;
    wire \c0.n21356 ;
    wire \c0.n22317 ;
    wire \c0.n6_adj_4305 ;
    wire \c0.n24119 ;
    wire \c0.n21050 ;
    wire \c0.n6_adj_4402 ;
    wire \c0.n22188 ;
    wire \c0.n20658_cascade_ ;
    wire \c0.n22166 ;
    wire \c0.n10467 ;
    wire \c0.n22180 ;
    wire \c0.n20330 ;
    wire \c0.n10434 ;
    wire \c0.n10513 ;
    wire \c0.n21189 ;
    wire \c0.n21135 ;
    wire \c0.n21219 ;
    wire \c0.n21811 ;
    wire \c0.n21135_cascade_ ;
    wire \c0.n6_adj_4497_cascade_ ;
    wire \c0.n20151 ;
    wire \c0.data_out_frame_29_6 ;
    wire \c0.n21848 ;
    wire \c0.n20253 ;
    wire \c0.n21852_cascade_ ;
    wire \c0.n22346 ;
    wire \c0.n22126 ;
    wire \c0.n20298 ;
    wire \c0.n10_adj_4512_cascade_ ;
    wire \c0.n10496 ;
    wire \c0.n20274 ;
    wire \c0.n21231 ;
    wire \c0.n22736 ;
    wire \c0.n21162_cascade_ ;
    wire \c0.n12526 ;
    wire \c0.n20201 ;
    wire \c0.n21876 ;
    wire data_out_frame_13_7;
    wire \c0.n21056 ;
    wire \c0.n22177 ;
    wire \c0.n22072 ;
    wire \c0.n22072_cascade_ ;
    wire \c0.n22073 ;
    wire \c0.n20175 ;
    wire \c0.n20249_cascade_ ;
    wire \c0.n12528 ;
    wire \c0.n21065 ;
    wire \c0.n21842 ;
    wire \c0.n20230 ;
    wire \c0.n6_adj_4394 ;
    wire encoder1_position_5;
    wire \c0.n22163_cascade_ ;
    wire \c0.n20_adj_4505 ;
    wire \c0.n19_adj_4506_cascade_ ;
    wire \c0.n21283 ;
    wire \c0.n6_adj_4508 ;
    wire \c0.n21116 ;
    wire \c0.n20819 ;
    wire \c0.n21_adj_4507 ;
    wire \c0.n20276 ;
    wire \c0.n21122 ;
    wire \c0.n21166 ;
    wire \c0.n13480 ;
    wire \c0.n22078 ;
    wire encoder1_position_9;
    wire \c0.n21112 ;
    wire \c0.n21253 ;
    wire \c0.n20180_cascade_ ;
    wire \c0.data_out_frame_29__7__N_1144 ;
    wire \c0.n20465 ;
    wire \c0.n21943 ;
    wire \c0.n21196 ;
    wire encoder1_position_25;
    wire encoder1_position_11;
    wire \c0.n20232_cascade_ ;
    wire \c0.n21146 ;
    wire \c0.n21146_cascade_ ;
    wire encoder1_position_23;
    wire \c0.n20232 ;
    wire \c0.n20744 ;
    wire encoder1_position_1;
    wire \c0.n20160 ;
    wire bfn_14_14_0_;
    wire \quad_counter0.count_direction ;
    wire \quad_counter0.n19580 ;
    wire n2270;
    wire \quad_counter0.n19581 ;
    wire n2269;
    wire \quad_counter0.n19582 ;
    wire n2268;
    wire \quad_counter0.n19583 ;
    wire \quad_counter0.n19584 ;
    wire \quad_counter0.n19585 ;
    wire \quad_counter0.n19586 ;
    wire \quad_counter0.n19587 ;
    wire encoder0_position_7;
    wire n2264;
    wire bfn_14_15_0_;
    wire \quad_counter0.n19588 ;
    wire \quad_counter0.n19589 ;
    wire \quad_counter0.n19590 ;
    wire \quad_counter0.n19591 ;
    wire \quad_counter0.n19592 ;
    wire n2258;
    wire \quad_counter0.n19593 ;
    wire n2257;
    wire \quad_counter0.n19594 ;
    wire \quad_counter0.n19595 ;
    wire bfn_14_16_0_;
    wire \quad_counter0.n19596 ;
    wire \quad_counter0.n19597 ;
    wire \quad_counter0.n19598 ;
    wire n2252;
    wire \quad_counter0.n19599 ;
    wire n2251;
    wire \quad_counter0.n19600 ;
    wire \quad_counter0.n19601 ;
    wire \quad_counter0.n19602 ;
    wire \quad_counter0.n19603 ;
    wire bfn_14_17_0_;
    wire \quad_counter0.n19604 ;
    wire \quad_counter0.n19605 ;
    wire \quad_counter0.n19606 ;
    wire encoder0_position_27;
    wire n2244;
    wire \quad_counter0.n19607 ;
    wire \quad_counter0.n19608 ;
    wire \quad_counter0.n19609 ;
    wire n2241;
    wire \quad_counter0.n19610 ;
    wire \quad_counter0.n19611 ;
    wire \quad_counter0.n2227 ;
    wire bfn_14_18_0_;
    wire \c0.n14474_cascade_ ;
    wire data_out_frame_9_1;
    wire data_out_frame_8_1;
    wire \c0.n24186 ;
    wire n2248;
    wire n2240;
    wire data_out_frame_7_7;
    wire data_out_frame_5_1;
    wire data_out_frame_8_0;
    wire data_out_frame_7_1;
    wire \c0.n24093 ;
    wire \c0.n5_adj_4518_cascade_ ;
    wire \c0.n23862 ;
    wire \c0.byte_transmit_counter_2 ;
    wire data_out_frame_5_7;
    wire \c0.n24054 ;
    wire \c0.tx.r_SM_Main_0 ;
    wire \c0.tx.n7086 ;
    wire data_in_2_3;
    wire data_in_2_1;
    wire \c0.n13_adj_4388_cascade_ ;
    wire \c0.n23135 ;
    wire \quad_counter0.b_delay_counter_14 ;
    wire \quad_counter0.b_delay_counter_7 ;
    wire \quad_counter0.b_delay_counter_12 ;
    wire \quad_counter0.b_delay_counter_15 ;
    wire \quad_counter0.n27_adj_4200 ;
    wire \c0.n14457 ;
    wire \c0.FRAME_MATCHER_state_22 ;
    wire \c0.n14457_cascade_ ;
    wire \c0.FRAME_MATCHER_state_27 ;
    wire \c0.n21330 ;
    wire \c0.n30_adj_4411_cascade_ ;
    wire \c0.FRAME_MATCHER_state_8 ;
    wire \c0.n21344 ;
    wire \c0.n21336 ;
    wire \c0.n44_adj_4412 ;
    wire \c0.FRAME_MATCHER_state_14 ;
    wire \c0.FRAME_MATCHER_state_21 ;
    wire \c0.n21368 ;
    wire \c0.FRAME_MATCHER_state_29 ;
    wire \c0.n21326 ;
    wire \c0.n20658 ;
    wire \c0.n21152 ;
    wire \c0.n21168 ;
    wire \c0.n12542 ;
    wire \c0.n20180 ;
    wire \c0.n23260 ;
    wire \c0.n16_adj_4498_cascade_ ;
    wire \c0.n21998 ;
    wire \c0.n21852 ;
    wire \c0.n20249 ;
    wire \c0.n21210 ;
    wire \c0.n17_adj_4499 ;
    wire \c0.data_out_frame_29_7 ;
    wire \c0.data_out_frame_28_7 ;
    wire \c0.n26_adj_4359 ;
    wire data_out_frame_13_1;
    wire data_out_frame_12_1;
    wire \c0.n11_adj_4520 ;
    wire data_out_frame_8_3;
    wire \c0.n11_adj_4303 ;
    wire encoder1_position_12;
    wire data_out_frame_12_4;
    wire encoder1_position_8;
    wire data_out_frame_12_0;
    wire \c0.n13079 ;
    wire \c0.n22174 ;
    wire data_in_3_5;
    wire encoder1_position_10;
    wire data_out_frame_12_2;
    wire \c0.n21918 ;
    wire encoder1_position_4;
    wire data_out_frame_13_4;
    wire encoder1_position_2;
    wire data_out_frame_13_2;
    wire encoder1_position_6;
    wire encoder1_position_7;
    wire \c0.n21896 ;
    wire encoder1_position_26;
    wire \c0.n20236 ;
    wire \c0.n22449 ;
    wire \c0.n22474 ;
    wire \c0.n22483 ;
    wire encoder1_position_30;
    wire \c0.n16_adj_4321_cascade_ ;
    wire \c0.n18_adj_4322_cascade_ ;
    wire \c0.n17_adj_4323 ;
    wire \c0.n14_adj_4324 ;
    wire \c0.n22376 ;
    wire \c0.n13619 ;
    wire \c0.n13619_cascade_ ;
    wire \c0.n22412 ;
    wire \c0.n13524_cascade_ ;
    wire \c0.n10_adj_4317 ;
    wire \c0.n20328 ;
    wire encoder0_position_14;
    wire \c0.n20328_cascade_ ;
    wire \c0.n22367 ;
    wire \c0.n22367_cascade_ ;
    wire \c0.n23569 ;
    wire n2271;
    wire \c0.n10_adj_4331 ;
    wire \c0.n22230 ;
    wire encoder0_position_1;
    wire \c0.n22461_cascade_ ;
    wire encoder0_position_13;
    wire \c0.n20_adj_4318 ;
    wire n2265;
    wire encoder0_position_6;
    wire encoder0_position_20;
    wire n2266;
    wire encoder0_position_5;
    wire \c0.n21808 ;
    wire n2250;
    wire encoder0_position_21;
    wire n2262;
    wire n2260;
    wire n2254;
    wire \c0.n10394 ;
    wire encoder0_position_17;
    wire encoder1_position_28;
    wire \c0.n13338 ;
    wire data_in_2_5;
    wire data_in_1_3;
    wire \c0.n16_adj_4478 ;
    wire data_in_1_1;
    wire data_in_0_1;
    wire data_out_frame_6_5;
    wire n2256;
    wire encoder0_position_15;
    wire data_in_2_0;
    wire n2247;
    wire n2242;
    wire data_in_3_6;
    wire data_in_2_6;
    wire data_out_frame_10_1;
    wire \c0.byte_transmit_counter_1 ;
    wire \c0.n24183 ;
    wire data_in_3_7;
    wire data_in_2_7;
    wire data_in_3_2;
    wire encoder1_position_17;
    wire data_out_frame_11_1;
    wire \c0.n9_adj_4415_cascade_ ;
    wire n14252;
    wire \c0.n38_adj_4387 ;
    wire \c0.tx_active ;
    wire \c0.n22651 ;
    wire n22661_cascade_;
    wire data_out_frame_7_3;
    wire data_out_frame_6_1;
    wire encoder0_position_0;
    wire data_out_frame_9_0;
    wire \c0.n21789 ;
    wire \c0.n12996_cascade_ ;
    wire \c0.n13020_cascade_ ;
    wire \c0.data_out_frame_29_7_N_1483_1_cascade_ ;
    wire \c0.n6650 ;
    wire \c0.n6650_cascade_ ;
    wire \c0.n6_adj_4270 ;
    wire \c0.n117 ;
    wire \c0.n63_adj_4301 ;
    wire \c0.n16958_cascade_ ;
    wire \c0.n63 ;
    wire \c0.n22695_cascade_ ;
    wire \c0.FRAME_MATCHER_state_2 ;
    wire \c0.n13_adj_4388 ;
    wire \c0.n9207 ;
    wire \c0.n14_adj_4337 ;
    wire \c0.n7_adj_4352_cascade_ ;
    wire \c0.FRAME_MATCHER_state_26 ;
    wire \c0.n48_cascade_ ;
    wire \c0.n45_adj_4413 ;
    wire \c0.FRAME_MATCHER_state_23 ;
    wire \c0.n14_adj_4316 ;
    wire \c0.FRAME_MATCHER_state_24 ;
    wire \c0.n21372 ;
    wire \c0.n21346 ;
    wire \c0.n21364 ;
    wire \c0.FRAME_MATCHER_state_9 ;
    wire \c0.n46 ;
    wire \c0.n20_adj_4482 ;
    wire \c0.n21_adj_4480_cascade_ ;
    wire \c0.n19_adj_4481 ;
    wire \c0.n14789 ;
    wire \c0.FRAME_MATCHER_state_18 ;
    wire \c0.FRAME_MATCHER_state_16 ;
    wire \c0.FRAME_MATCHER_state_17 ;
    wire \c0.n21682 ;
    wire \c0.FRAME_MATCHER_state_4 ;
    wire \c0.n47 ;
    wire \c0.FRAME_MATCHER_state_25 ;
    wire \c0.n21374 ;
    wire \c0.FRAME_MATCHER_state_10 ;
    wire \c0.n21348 ;
    wire \c0.FRAME_MATCHER_state_7 ;
    wire \c0.n21342 ;
    wire \c0.FRAME_MATCHER_state_11 ;
    wire \c0.n21350 ;
    wire encoder1_position_13;
    wire data_out_frame_12_5;
    wire \c0.n14_adj_4364 ;
    wire \c0.n13 ;
    wire \c0.n13_adj_4366_cascade_ ;
    wire \c0.n14_adj_4365 ;
    wire \c0.n14_adj_4400 ;
    wire \c0.n17600_cascade_ ;
    wire \c0.data_in_frame_10_4 ;
    wire \c0.n21908 ;
    wire count_enable_adj_4544;
    wire n2185;
    wire \c0.n13839 ;
    wire \c0.n22015 ;
    wire encoder0_position_29;
    wire \c0.data_out_frame_29__7__N_856 ;
    wire \c0.n22382 ;
    wire \c0.n6_adj_4311 ;
    wire \c0.n22427 ;
    wire encoder0_position_19;
    wire \c0.n21885 ;
    wire \c0.n22200 ;
    wire \c0.n22200_cascade_ ;
    wire \c0.n21970 ;
    wire \c0.n13705 ;
    wire n2259;
    wire n2267;
    wire n2261;
    wire n2255;
    wire encoder0_position_16;
    wire \c0.n22408 ;
    wire encoder0_position_4;
    wire \c0.n22227_cascade_ ;
    wire \c0.n22128 ;
    wire \c0.n10444 ;
    wire encoder1_position_20;
    wire \c0.n6_adj_4312 ;
    wire encoder0_position_12;
    wire \c0.n22477 ;
    wire \c0.n22477_cascade_ ;
    wire \c0.n6_adj_4333 ;
    wire n2243;
    wire encoder0_position_28;
    wire encoder0_position_9;
    wire \c0.n6_adj_4315_cascade_ ;
    wire \c0.n20171 ;
    wire \c0.data_out_frame_29__7__N_847 ;
    wire \c0.data_out_frame_29__7__N_847_cascade_ ;
    wire encoder0_position_11;
    wire \c0.n10_adj_4332 ;
    wire encoder0_position_24;
    wire \c0.n21931 ;
    wire \c0.r_SM_Main_2_N_3755_0 ;
    wire \c0.n14322 ;
    wire \c0.n14322_cascade_ ;
    wire \c0.n14871 ;
    wire \c0.tx_transmit_N_3651 ;
    wire \c0.n23975 ;
    wire \c0.n18_adj_4403 ;
    wire \c0.n20875 ;
    wire \c0.n17602 ;
    wire \c0.n17602_cascade_ ;
    wire \c0.n8_adj_4417 ;
    wire n2245;
    wire encoder0_position_26;
    wire n2263;
    wire encoder0_position_10;
    wire data_out_frame_8_2;
    wire n2246;
    wire encoder0_position_25;
    wire data_out_frame_7_6;
    wire \c0.byte_transmit_counter_0 ;
    wire \c0.n5_adj_4350 ;
    wire control_mode_2;
    wire encoder0_position_23;
    wire encoder0_position_8;
    wire \c0.n22032 ;
    wire data_in_3_0;
    wire control_mode_5;
    wire \c0.n23215_cascade_ ;
    wire data_out_frame_29_7_N_1483_2;
    wire \c0.n6_adj_4338 ;
    wire \c0.data_out_frame_0__7__N_2568_cascade_ ;
    wire \c0.n1220_cascade_ ;
    wire \c0.n4_adj_4373 ;
    wire \c0.n5024_cascade_ ;
    wire \c0.n21773 ;
    wire \c0.n21773_cascade_ ;
    wire \c0.data_out_frame_29_7_N_1483_1 ;
    wire \c0.n4_adj_4328_cascade_ ;
    wire \c0.data_out_frame_0__7__N_2568 ;
    wire \c0.FRAME_MATCHER_state_1 ;
    wire \c0.n4_adj_4391 ;
    wire \c0.n38_adj_4390 ;
    wire \c0.n8107 ;
    wire \c0.n49 ;
    wire \c0.n50 ;
    wire \c0.n54 ;
    wire \c0.n22665 ;
    wire \c0.n3239 ;
    wire \c0.n63_adj_4293_cascade_ ;
    wire \c0.n13020 ;
    wire \c0.n4_adj_4345 ;
    wire \c0.n84_cascade_ ;
    wire \c0.n12990 ;
    wire \c0.n7_adj_4344 ;
    wire \c0.n12967 ;
    wire \c0.FRAME_MATCHER_state_0 ;
    wire \c0.n12996 ;
    wire \c0.n4_adj_4419 ;
    wire \c0.FRAME_MATCHER_state_30 ;
    wire \c0.n8_adj_4396 ;
    wire \c0.n21737_cascade_ ;
    wire \c0.FRAME_MATCHER_state_6 ;
    wire \c0.n21340 ;
    wire \c0.FRAME_MATCHER_state_19 ;
    wire \c0.n8_adj_4398 ;
    wire \c0.FRAME_MATCHER_state_5 ;
    wire \c0.n21338 ;
    wire \c0.n38_adj_4407_cascade_ ;
    wire \c0.n23836 ;
    wire \c0.n43_adj_4410_cascade_ ;
    wire \c0.n22443_cascade_ ;
    wire \c0.n21986_cascade_ ;
    wire data_in_frame_6_0;
    wire \c0.n6_adj_4393_cascade_ ;
    wire \c0.n13086_cascade_ ;
    wire \c0.n25_adj_4408 ;
    wire \c0.n23648 ;
    wire \c0.n16_adj_4401 ;
    wire \c0.n21893 ;
    wire \c0.n44_adj_4409 ;
    wire \c0.data_in_frame_20_6 ;
    wire n21744_cascade_;
    wire data_in_frame_6_3;
    wire n2253;
    wire \c0.n21816 ;
    wire \c0.n21740_cascade_ ;
    wire encoder0_position_18;
    wire encoder0_position_3;
    wire encoder0_position_31;
    wire \c0.n21813 ;
    wire data_in_frame_6_5;
    wire \c0.tx.n23987 ;
    wire \c0.tx.r_Clock_Count_6 ;
    wire n313;
    wire r_SM_Main_2_adj_4549;
    wire n8;
    wire r_Clock_Count_8;
    wire n2249;
    wire count_enable;
    wire encoder0_position_22;
    wire data_in_2_4;
    wire data_in_1_4;
    wire \c0.FRAME_MATCHER_rx_data_ready_prev ;
    wire \c0.n17790_cascade_ ;
    wire \c0.n21775_cascade_ ;
    wire data_in_3_4;
    wire control_mode_1;
    wire control_mode_3;
    wire control_mode_4;
    wire control_mode_7;
    wire n23726_cascade_;
    wire control_mode_6;
    wire \c0.n12876 ;
    wire \c0.n21022 ;
    wire \c0.n12991 ;
    wire \c0.n5024 ;
    wire \c0.n5_adj_4342_cascade_ ;
    wire \c0.n21686 ;
    wire \c0.FRAME_MATCHER_state_3 ;
    wire \c0.n21686_cascade_ ;
    wire \c0.n21334 ;
    wire \c0.n44_adj_4336 ;
    wire \c0.n1_adj_4349 ;
    wire \c0.n21734 ;
    wire \c0.n13021 ;
    wire \c0.n23965 ;
    wire \c0.n22575 ;
    wire \c0.n45_adj_4389 ;
    wire rx_data_ready;
    wire data_in_3_1;
    wire \c0.n1 ;
    wire \c0.n19783 ;
    wire \c0.n937 ;
    wire \c0.FRAME_MATCHER_state_12 ;
    wire \c0.n21352 ;
    wire \c0.n20_adj_4327 ;
    wire \c0.n12992 ;
    wire \c0.n9668 ;
    wire \c0.n7_adj_4356 ;
    wire \c0.FRAME_MATCHER_state_28 ;
    wire \c0.n21378 ;
    wire \c0.FRAME_MATCHER_state_31 ;
    wire \c0.n21332 ;
    wire \c0.FRAME_MATCHER_state_13 ;
    wire \c0.n21354 ;
    wire \c0.FRAME_MATCHER_state_15 ;
    wire \c0.n21358 ;
    wire \c0.n21957 ;
    wire \c0.n21957_cascade_ ;
    wire \c0.n22287 ;
    wire \c0.data_in_frame_3_3 ;
    wire \c0.data_in_frame_5_4 ;
    wire \c0.n23838 ;
    wire \c0.n21902_cascade_ ;
    wire \c0.data_in_frame_3_0 ;
    wire \c0.n21902 ;
    wire \c0.data_in_frame_5_2 ;
    wire \c0.n21879_cascade_ ;
    wire \c0.data_in_frame_3_4 ;
    wire \c0.n22290 ;
    wire \c0.n22258 ;
    wire \c0.n22258_cascade_ ;
    wire \c0.n29_adj_4374 ;
    wire \c0.n27_adj_4377_cascade_ ;
    wire \c0.n14072_cascade_ ;
    wire \c0.n14072 ;
    wire \c0.n6_adj_4385_cascade_ ;
    wire \c0.n21803 ;
    wire \c0.n18_adj_4370 ;
    wire \c0.n22194 ;
    wire \c0.n21803_cascade_ ;
    wire \c0.n30_adj_4371 ;
    wire \c0.data_in_frame_0_1 ;
    wire \c0.data_in_frame_0_0 ;
    wire \c0.n13376_cascade_ ;
    wire \c0.n13376 ;
    wire data_in_frame_1_6;
    wire data_in_frame_6_2;
    wire \c0.n13386_cascade_ ;
    wire \c0.data_in_frame_4_4 ;
    wire \c0.n22261 ;
    wire \c0.data_in_frame_2_1 ;
    wire \c0.n22261_cascade_ ;
    wire \c0.n22320 ;
    wire \c0.n28_adj_4372 ;
    wire \c0.data_in_frame_3_6 ;
    wire \c0.data_in_frame_4_1 ;
    wire \c0.n22218 ;
    wire \c0.n21928_cascade_ ;
    wire \c0.data_in_frame_2_3 ;
    wire \c0.n21791 ;
    wire \c0.n21882_cascade_ ;
    wire \c0.data_out_frame_0__7__N_2744 ;
    wire \c0.data_out_frame_0__7__N_2744_cascade_ ;
    wire \c0.n6_adj_4272_cascade_ ;
    wire \c0.data_in_frame_3_7 ;
    wire \c0.data_in_frame_4_7 ;
    wire \c0.data_in_frame_5_1 ;
    wire \c0.n21992 ;
    wire \c0.data_in_frame_2_2 ;
    wire data_in_frame_1_7;
    wire \c0.n39_adj_4406 ;
    wire data_in_frame_6_7;
    wire \c0.n21882 ;
    wire \c0.n21928 ;
    wire \c0.n14037_cascade_ ;
    wire \c0.n6_adj_4369 ;
    wire \c0.n5_adj_4368 ;
    wire \c0.data_out_frame_29__7__N_1474 ;
    wire data_in_frame_6_6;
    wire \c0.data_in_frame_0_2 ;
    wire \c0.data_in_frame_2_4 ;
    wire \c0.data_in_frame_5_0 ;
    wire \c0.data_in_frame_2_0 ;
    wire data_in_frame_6_1;
    wire n4_cascade_;
    wire \c0.data_in_frame_4_6 ;
    wire n4;
    wire \c0.n21758_cascade_ ;
    wire \c0.n17790 ;
    wire data_in_frame_1_0;
    wire n23726;
    wire control_mode_0;
    wire \c0.data_in_frame_29_4 ;
    wire \c0.n10_adj_4286_cascade_ ;
    wire \c0.data_in_frame_28_2 ;
    wire \c0.data_in_frame_29_0 ;
    wire \c0.n17600 ;
    wire \c0.n19_cascade_ ;
    wire \c0.n23389 ;
    wire \c0.n32_adj_4295_cascade_ ;
    wire \c0.n23523 ;
    wire \c0.n34 ;
    wire \c0.data_in_frame_29_2 ;
    wire \c0.data_in_frame_29_1 ;
    wire \c0.n23388_cascade_ ;
    wire \c0.n30_adj_4299 ;
    wire \c0.n15_adj_4376_cascade_ ;
    wire \c0.n17_adj_4378 ;
    wire \c0.n18_adj_4379_cascade_ ;
    wire \c0.n27_adj_4383 ;
    wire \c0.n30_adj_4380_cascade_ ;
    wire \c0.n28_adj_4381 ;
    wire \c0.n13000 ;
    wire data_in_frame_22_1;
    wire \c0.rx.n22611_cascade_ ;
    wire \c0.rx.n8_cascade_ ;
    wire \c0.n29_adj_4382 ;
    wire \c0.n161 ;
    wire bfn_19_1_0_;
    wire \c0.n3 ;
    wire \c0.n19442 ;
    wire \c0.n19442_THRU_CRY_0_THRU_CO ;
    wire \c0.n19442_THRU_CRY_1_THRU_CO ;
    wire \c0.n19442_THRU_CRY_2_THRU_CO ;
    wire \c0.n19442_THRU_CRY_3_THRU_CO ;
    wire \c0.n19442_THRU_CRY_4_THRU_CO ;
    wire \c0.n19442_THRU_CRY_5_THRU_CO ;
    wire \c0.n19442_THRU_CRY_6_THRU_CO ;
    wire bfn_19_2_0_;
    wire \c0.n19443 ;
    wire \c0.n19443_THRU_CRY_0_THRU_CO ;
    wire \c0.n19443_THRU_CRY_1_THRU_CO ;
    wire \c0.n19443_THRU_CRY_2_THRU_CO ;
    wire \c0.n19443_THRU_CRY_3_THRU_CO ;
    wire \c0.n19443_THRU_CRY_4_THRU_CO ;
    wire \c0.n19443_THRU_CRY_5_THRU_CO ;
    wire \c0.n19443_THRU_CRY_6_THRU_CO ;
    wire bfn_19_3_0_;
    wire \c0.n19444 ;
    wire \c0.n19444_THRU_CRY_0_THRU_CO ;
    wire \c0.n19444_THRU_CRY_1_THRU_CO ;
    wire \c0.n19444_THRU_CRY_2_THRU_CO ;
    wire \c0.n19444_THRU_CRY_3_THRU_CO ;
    wire \c0.n19444_THRU_CRY_4_THRU_CO ;
    wire \c0.n19444_THRU_CRY_5_THRU_CO ;
    wire \c0.n19444_THRU_CRY_6_THRU_CO ;
    wire bfn_19_4_0_;
    wire \c0.n19445 ;
    wire \c0.n19445_THRU_CRY_0_THRU_CO ;
    wire \c0.n19445_THRU_CRY_1_THRU_CO ;
    wire \c0.n19445_THRU_CRY_2_THRU_CO ;
    wire \c0.n19445_THRU_CRY_3_THRU_CO ;
    wire \c0.n19445_THRU_CRY_4_THRU_CO ;
    wire \c0.n19445_THRU_CRY_5_THRU_CO ;
    wire \c0.n19445_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_4 ;
    wire bfn_19_5_0_;
    wire \c0.n3_adj_4470 ;
    wire \c0.n19446 ;
    wire \c0.n19446_THRU_CRY_0_THRU_CO ;
    wire \c0.n19446_THRU_CRY_1_THRU_CO ;
    wire \c0.n19446_THRU_CRY_2_THRU_CO ;
    wire \c0.n19446_THRU_CRY_3_THRU_CO ;
    wire \c0.n19446_THRU_CRY_4_THRU_CO ;
    wire \c0.n19446_THRU_CRY_5_THRU_CO ;
    wire \c0.n19446_THRU_CRY_6_THRU_CO ;
    wire bfn_19_6_0_;
    wire \c0.n3_adj_4468 ;
    wire \c0.n19447 ;
    wire \c0.n19447_THRU_CRY_0_THRU_CO ;
    wire \c0.n19447_THRU_CRY_1_THRU_CO ;
    wire \c0.n19447_THRU_CRY_2_THRU_CO ;
    wire \c0.n19447_THRU_CRY_3_THRU_CO ;
    wire \c0.n19447_THRU_CRY_4_THRU_CO ;
    wire \c0.n19447_THRU_CRY_5_THRU_CO ;
    wire \c0.n19447_THRU_CRY_6_THRU_CO ;
    wire bfn_19_7_0_;
    wire \c0.n3_adj_4467 ;
    wire \c0.n19448 ;
    wire \c0.n19448_THRU_CRY_0_THRU_CO ;
    wire \c0.n19448_THRU_CRY_1_THRU_CO ;
    wire \c0.n19448_THRU_CRY_2_THRU_CO ;
    wire \c0.n19448_THRU_CRY_3_THRU_CO ;
    wire \c0.n19448_THRU_CRY_4_THRU_CO ;
    wire \c0.n19448_THRU_CRY_5_THRU_CO ;
    wire \c0.n19448_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_7 ;
    wire bfn_19_8_0_;
    wire \c0.n3_adj_4465 ;
    wire \c0.n19449 ;
    wire \c0.n19449_THRU_CRY_0_THRU_CO ;
    wire \c0.n19449_THRU_CRY_1_THRU_CO ;
    wire \c0.n19449_THRU_CRY_2_THRU_CO ;
    wire \c0.n19449_THRU_CRY_3_THRU_CO ;
    wire \c0.n19449_THRU_CRY_4_THRU_CO ;
    wire \c0.n19449_THRU_CRY_5_THRU_CO ;
    wire \c0.n19449_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_8 ;
    wire bfn_19_9_0_;
    wire \c0.n3_adj_4463 ;
    wire \c0.n19450 ;
    wire \c0.n19450_THRU_CRY_0_THRU_CO ;
    wire \c0.n19450_THRU_CRY_1_THRU_CO ;
    wire \c0.n19450_THRU_CRY_2_THRU_CO ;
    wire \c0.n19450_THRU_CRY_3_THRU_CO ;
    wire \c0.n19450_THRU_CRY_4_THRU_CO ;
    wire \c0.n19450_THRU_CRY_5_THRU_CO ;
    wire \c0.n19450_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_9 ;
    wire bfn_19_10_0_;
    wire \c0.n3_adj_4462 ;
    wire \c0.n19451 ;
    wire \c0.n19451_THRU_CRY_0_THRU_CO ;
    wire \c0.n19451_THRU_CRY_1_THRU_CO ;
    wire \c0.n19451_THRU_CRY_2_THRU_CO ;
    wire \c0.n19451_THRU_CRY_3_THRU_CO ;
    wire \c0.n19451_THRU_CRY_4_THRU_CO ;
    wire \c0.n19451_THRU_CRY_5_THRU_CO ;
    wire \c0.n19451_THRU_CRY_6_THRU_CO ;
    wire bfn_19_11_0_;
    wire \c0.n19452 ;
    wire \c0.n19452_THRU_CRY_0_THRU_CO ;
    wire \c0.n19452_THRU_CRY_1_THRU_CO ;
    wire \c0.n19452_THRU_CRY_2_THRU_CO ;
    wire \c0.n19452_THRU_CRY_3_THRU_CO ;
    wire \c0.n19452_THRU_CRY_4_THRU_CO ;
    wire \c0.n19452_THRU_CRY_5_THRU_CO ;
    wire \c0.n19452_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_11 ;
    wire bfn_19_12_0_;
    wire \c0.n3_adj_4458 ;
    wire \c0.n19453 ;
    wire \c0.n19453_THRU_CRY_0_THRU_CO ;
    wire \c0.n19453_THRU_CRY_1_THRU_CO ;
    wire \c0.n19453_THRU_CRY_2_THRU_CO ;
    wire \c0.n19453_THRU_CRY_3_THRU_CO ;
    wire \c0.n19453_THRU_CRY_4_THRU_CO ;
    wire \c0.n19453_THRU_CRY_5_THRU_CO ;
    wire \c0.n19453_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_12 ;
    wire bfn_19_13_0_;
    wire \c0.n3_adj_4456 ;
    wire \c0.n19454 ;
    wire \c0.n19454_THRU_CRY_0_THRU_CO ;
    wire \c0.n19454_THRU_CRY_1_THRU_CO ;
    wire \c0.n19454_THRU_CRY_2_THRU_CO ;
    wire \c0.n19454_THRU_CRY_3_THRU_CO ;
    wire \c0.n19454_THRU_CRY_4_THRU_CO ;
    wire \c0.n19454_THRU_CRY_5_THRU_CO ;
    wire \c0.n19454_THRU_CRY_6_THRU_CO ;
    wire bfn_19_14_0_;
    wire \c0.n19455 ;
    wire \c0.n19455_THRU_CRY_0_THRU_CO ;
    wire \c0.n19455_THRU_CRY_1_THRU_CO ;
    wire \c0.n19455_THRU_CRY_2_THRU_CO ;
    wire \c0.n19455_THRU_CRY_3_THRU_CO ;
    wire \c0.n19455_THRU_CRY_4_THRU_CO ;
    wire \c0.n19455_THRU_CRY_5_THRU_CO ;
    wire \c0.n19455_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_14 ;
    wire bfn_19_15_0_;
    wire \c0.n3_adj_4453 ;
    wire \c0.n19456 ;
    wire \c0.n19456_THRU_CRY_0_THRU_CO ;
    wire \c0.n19456_THRU_CRY_1_THRU_CO ;
    wire \c0.n19456_THRU_CRY_2_THRU_CO ;
    wire \c0.n19456_THRU_CRY_3_THRU_CO ;
    wire \c0.n19456_THRU_CRY_4_THRU_CO ;
    wire \c0.n19456_THRU_CRY_5_THRU_CO ;
    wire \c0.n19456_THRU_CRY_6_THRU_CO ;
    wire bfn_19_16_0_;
    wire \c0.n19457 ;
    wire \c0.n19457_THRU_CRY_0_THRU_CO ;
    wire \c0.n19457_THRU_CRY_1_THRU_CO ;
    wire \c0.n19457_THRU_CRY_2_THRU_CO ;
    wire \c0.n19457_THRU_CRY_3_THRU_CO ;
    wire \c0.n19457_THRU_CRY_4_THRU_CO ;
    wire \c0.n19457_THRU_CRY_5_THRU_CO ;
    wire \c0.n19457_THRU_CRY_6_THRU_CO ;
    wire bfn_19_17_0_;
    wire \c0.n3_adj_4450 ;
    wire \c0.n19458 ;
    wire \c0.n19458_THRU_CRY_0_THRU_CO ;
    wire \c0.n19458_THRU_CRY_1_THRU_CO ;
    wire \c0.n19458_THRU_CRY_2_THRU_CO ;
    wire \c0.n19458_THRU_CRY_3_THRU_CO ;
    wire \c0.n19458_THRU_CRY_4_THRU_CO ;
    wire \c0.n19458_THRU_CRY_5_THRU_CO ;
    wire \c0.n19458_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_17 ;
    wire bfn_19_18_0_;
    wire \c0.n3_adj_4448 ;
    wire \c0.n19459 ;
    wire \c0.n19459_THRU_CRY_0_THRU_CO ;
    wire \c0.n19459_THRU_CRY_1_THRU_CO ;
    wire \c0.n19459_THRU_CRY_2_THRU_CO ;
    wire \c0.n19459_THRU_CRY_3_THRU_CO ;
    wire \c0.n19459_THRU_CRY_4_THRU_CO ;
    wire \c0.n19459_THRU_CRY_5_THRU_CO ;
    wire \c0.n19459_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_18 ;
    wire bfn_19_19_0_;
    wire \c0.n3_adj_4446 ;
    wire \c0.n19460 ;
    wire \c0.n19460_THRU_CRY_0_THRU_CO ;
    wire \c0.n19460_THRU_CRY_1_THRU_CO ;
    wire \c0.n19460_THRU_CRY_2_THRU_CO ;
    wire \c0.n19460_THRU_CRY_3_THRU_CO ;
    wire \c0.n19460_THRU_CRY_4_THRU_CO ;
    wire \c0.n19460_THRU_CRY_5_THRU_CO ;
    wire \c0.n19460_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_19 ;
    wire bfn_19_20_0_;
    wire \c0.n3_adj_4444 ;
    wire \c0.n19461 ;
    wire \c0.n19461_THRU_CRY_0_THRU_CO ;
    wire \c0.n19461_THRU_CRY_1_THRU_CO ;
    wire \c0.n19461_THRU_CRY_2_THRU_CO ;
    wire \c0.n19461_THRU_CRY_3_THRU_CO ;
    wire \c0.n19461_THRU_CRY_4_THRU_CO ;
    wire \c0.n19461_THRU_CRY_5_THRU_CO ;
    wire \c0.n19461_THRU_CRY_6_THRU_CO ;
    wire bfn_19_21_0_;
    wire \c0.n19462 ;
    wire \c0.n19462_THRU_CRY_0_THRU_CO ;
    wire \c0.n19462_THRU_CRY_1_THRU_CO ;
    wire \c0.n19462_THRU_CRY_2_THRU_CO ;
    wire \c0.n19462_THRU_CRY_3_THRU_CO ;
    wire \c0.n19462_THRU_CRY_4_THRU_CO ;
    wire \c0.n19462_THRU_CRY_5_THRU_CO ;
    wire \c0.n19462_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_21 ;
    wire bfn_19_22_0_;
    wire \c0.n3_adj_4440 ;
    wire \c0.n19463 ;
    wire \c0.n19463_THRU_CRY_0_THRU_CO ;
    wire \c0.n19463_THRU_CRY_1_THRU_CO ;
    wire \c0.n19463_THRU_CRY_2_THRU_CO ;
    wire \c0.n19463_THRU_CRY_3_THRU_CO ;
    wire \c0.n19463_THRU_CRY_4_THRU_CO ;
    wire \c0.n19463_THRU_CRY_5_THRU_CO ;
    wire \c0.n19463_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_22 ;
    wire bfn_19_23_0_;
    wire \c0.n3_adj_4438 ;
    wire \c0.n19464 ;
    wire \c0.n19464_THRU_CRY_0_THRU_CO ;
    wire \c0.n19464_THRU_CRY_1_THRU_CO ;
    wire \c0.n19464_THRU_CRY_2_THRU_CO ;
    wire \c0.n19464_THRU_CRY_3_THRU_CO ;
    wire \c0.n19464_THRU_CRY_4_THRU_CO ;
    wire \c0.n19464_THRU_CRY_5_THRU_CO ;
    wire \c0.n19464_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_23 ;
    wire bfn_19_24_0_;
    wire \c0.n3_adj_4436 ;
    wire \c0.n19465 ;
    wire \c0.n19465_THRU_CRY_0_THRU_CO ;
    wire \c0.n19465_THRU_CRY_1_THRU_CO ;
    wire \c0.n19465_THRU_CRY_2_THRU_CO ;
    wire \c0.n19465_THRU_CRY_3_THRU_CO ;
    wire \c0.n19465_THRU_CRY_4_THRU_CO ;
    wire \c0.n19465_THRU_CRY_5_THRU_CO ;
    wire \c0.n19465_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_24 ;
    wire bfn_19_25_0_;
    wire \c0.n3_adj_4435 ;
    wire \c0.n19466 ;
    wire \c0.n19466_THRU_CRY_0_THRU_CO ;
    wire \c0.n19466_THRU_CRY_1_THRU_CO ;
    wire \c0.n19466_THRU_CRY_2_THRU_CO ;
    wire \c0.n19466_THRU_CRY_3_THRU_CO ;
    wire \c0.n19466_THRU_CRY_4_THRU_CO ;
    wire \c0.n19466_THRU_CRY_5_THRU_CO ;
    wire \c0.n19466_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_25 ;
    wire bfn_19_26_0_;
    wire \c0.n3_adj_4434 ;
    wire \c0.n19467 ;
    wire \c0.n19467_THRU_CRY_0_THRU_CO ;
    wire \c0.n19467_THRU_CRY_1_THRU_CO ;
    wire \c0.n19467_THRU_CRY_2_THRU_CO ;
    wire \c0.n19467_THRU_CRY_3_THRU_CO ;
    wire \c0.n19467_THRU_CRY_4_THRU_CO ;
    wire \c0.n19467_THRU_CRY_5_THRU_CO ;
    wire \c0.n19467_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_26 ;
    wire bfn_19_27_0_;
    wire \c0.n3_adj_4433 ;
    wire \c0.n19468 ;
    wire \c0.n19468_THRU_CRY_0_THRU_CO ;
    wire \c0.n19468_THRU_CRY_1_THRU_CO ;
    wire \c0.n19468_THRU_CRY_2_THRU_CO ;
    wire \c0.n19468_THRU_CRY_3_THRU_CO ;
    wire \c0.n19468_THRU_CRY_4_THRU_CO ;
    wire \c0.n19468_THRU_CRY_5_THRU_CO ;
    wire \c0.n19468_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_27 ;
    wire bfn_19_28_0_;
    wire \c0.n3_adj_4432 ;
    wire \c0.n19469 ;
    wire \c0.n19469_THRU_CRY_0_THRU_CO ;
    wire \c0.n19469_THRU_CRY_1_THRU_CO ;
    wire \c0.n19469_THRU_CRY_2_THRU_CO ;
    wire \c0.n19469_THRU_CRY_3_THRU_CO ;
    wire \c0.n19469_THRU_CRY_4_THRU_CO ;
    wire \c0.n19469_THRU_CRY_5_THRU_CO ;
    wire \c0.n19469_THRU_CRY_6_THRU_CO ;
    wire bfn_19_29_0_;
    wire \c0.n19470 ;
    wire \c0.n19470_THRU_CRY_0_THRU_CO ;
    wire \c0.n19470_THRU_CRY_1_THRU_CO ;
    wire \c0.n19470_THRU_CRY_2_THRU_CO ;
    wire \c0.n19470_THRU_CRY_3_THRU_CO ;
    wire \c0.n19470_THRU_CRY_4_THRU_CO ;
    wire \c0.n19470_THRU_CRY_5_THRU_CO ;
    wire \c0.n19470_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_29 ;
    wire bfn_19_30_0_;
    wire \c0.n3_adj_4428 ;
    wire \c0.n19471 ;
    wire \c0.n19471_THRU_CRY_0_THRU_CO ;
    wire \c0.n19471_THRU_CRY_1_THRU_CO ;
    wire \c0.n19471_THRU_CRY_2_THRU_CO ;
    wire \c0.n19471_THRU_CRY_3_THRU_CO ;
    wire \c0.n19471_THRU_CRY_4_THRU_CO ;
    wire \c0.n19471_THRU_CRY_5_THRU_CO ;
    wire \c0.n19471_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_30 ;
    wire bfn_19_31_0_;
    wire \c0.n3_adj_4426 ;
    wire \c0.n19472 ;
    wire \c0.n19472_THRU_CRY_0_THRU_CO ;
    wire \c0.n19472_THRU_CRY_1_THRU_CO ;
    wire \c0.n19472_THRU_CRY_2_THRU_CO ;
    wire \c0.n19472_THRU_CRY_3_THRU_CO ;
    wire \c0.n19472_THRU_CRY_4_THRU_CO ;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire \c0.n19472_THRU_CRY_5_THRU_CO ;
    wire \c0.n19472_THRU_CRY_6_THRU_CO ;
    wire bfn_19_32_0_;
    wire \c0.FRAME_MATCHER_i_31 ;
    wire \c0.n3_adj_4421 ;
    wire \c0.n3_adj_4475 ;
    wire \c0.FRAME_MATCHER_i_3 ;
    wire \c0.n3_adj_4472 ;
    wire \c0.n3_adj_4474 ;
    wire \c0.FRAME_MATCHER_i_5 ;
    wire \c0.FRAME_MATCHER_i_6 ;
    wire \c0.n11_adj_4326 ;
    wire \c0.n10_adj_4399 ;
    wire \c0.n13033 ;
    wire \c0.data_in_frame_2_7 ;
    wire \c0.data_in_frame_0_7 ;
    wire \c0.data_in_frame_8_4 ;
    wire \c0.n21861_cascade_ ;
    wire \c0.n6_adj_4258 ;
    wire \c0.data_in_frame_9_5 ;
    wire \c0.n8_adj_4254_cascade_ ;
    wire \c0.n4_adj_4255 ;
    wire \c0.data_in_frame_5_5 ;
    wire \c0.data_in_frame_3_1 ;
    wire \c0.data_in_frame_3_2 ;
    wire \c0.n6_adj_4395 ;
    wire data_in_frame_1_1;
    wire data_in_frame_1_5;
    wire \c0.n21986 ;
    wire \c0.n13848_cascade_ ;
    wire \c0.n13_adj_4405 ;
    wire \c0.data_in_frame_2_5 ;
    wire \c0.data_in_frame_0_3 ;
    wire \c0.n13398 ;
    wire data_in_frame_1_3;
    wire \c0.data_in_frame_3_5 ;
    wire \c0.n13398_cascade_ ;
    wire \c0.n13852 ;
    wire \c0.n21794 ;
    wire \c0.data_in_frame_8_2 ;
    wire \c0.n21794_cascade_ ;
    wire \c0.data_in_frame_5_7 ;
    wire \c0.n6_adj_4257_cascade_ ;
    wire \c0.n21825 ;
    wire \c0.n13771_cascade_ ;
    wire \c0.n22239 ;
    wire \c0.n4_cascade_ ;
    wire \c0.n37 ;
    wire \c0.n6_adj_4220 ;
    wire \c0.data_in_frame_8_3 ;
    wire \c0.n13652 ;
    wire \c0.n13771 ;
    wire \c0.data_in_frame_10_3 ;
    wire \c0.n21964 ;
    wire \c0.n22280 ;
    wire \c0.n21964_cascade_ ;
    wire \c0.n14113 ;
    wire \c0.n6_adj_4241 ;
    wire \c0.n13086 ;
    wire \c0.data_in_frame_8_5 ;
    wire \c0.n22415_cascade_ ;
    wire \c0.data_in_frame_10_5 ;
    wire \c0.n35 ;
    wire n21744;
    wire \c0.n6_adj_4386 ;
    wire \c0.data_in_frame_4_3 ;
    wire data_in_frame_6_4;
    wire \c0.data_in_frame_4_2 ;
    wire FRAME_MATCHER_state_31_N_2976_2;
    wire n22661;
    wire encoder0_position_30;
    wire data_out_frame_6_6;
    wire \c0.n13697 ;
    wire \c0.n22440_cascade_ ;
    wire \c0.data_in_frame_10_7 ;
    wire \c0.n10_adj_4229_cascade_ ;
    wire \c0.n5943_cascade_ ;
    wire \c0.n22081_cascade_ ;
    wire \c0.n22349_cascade_ ;
    wire \c0.n21858_cascade_ ;
    wire \c0.FRAME_MATCHER_i_16 ;
    wire \c0.n16_adj_4375 ;
    wire \c0.FRAME_MATCHER_i_13 ;
    wire \c0.n3_adj_4454 ;
    wire \c0.FRAME_MATCHER_i_15 ;
    wire \c0.n3_adj_4452 ;
    wire \c0.FRAME_MATCHER_i_20 ;
    wire \c0.n3_adj_4442 ;
    wire \c0.data_in_frame_28_1 ;
    wire \c0.n21870_cascade_ ;
    wire \c0.data_in_frame_21_3 ;
    wire \c0.data_in_frame_23_5 ;
    wire \c0.data_in_frame_23_4 ;
    wire \c0.n10_adj_4287_cascade_ ;
    wire \c0.n22_adj_4298 ;
    wire \c0.n13266 ;
    wire \c0.data_in_frame_29_7 ;
    wire \c0.n21233_cascade_ ;
    wire \c0.n23506 ;
    wire \c0.data_in_frame_27_1 ;
    wire \c0.FRAME_MATCHER_i_10 ;
    wire \c0.n3_adj_4460 ;
    wire n18678;
    wire \c0.rx.n18655_cascade_ ;
    wire \c0.rx.n21704_cascade_ ;
    wire \c0.rx.n22573_cascade_ ;
    wire \c0.rx.n12_cascade_ ;
    wire bfn_20_24_0_;
    wire \c0.rx.r_Clock_Count_1 ;
    wire \c0.rx.n19533 ;
    wire \c0.rx.r_Clock_Count_2 ;
    wire \c0.rx.n19534 ;
    wire \c0.rx.r_Clock_Count_3 ;
    wire \c0.rx.n19535 ;
    wire \c0.rx.n19536 ;
    wire \c0.rx.n19537 ;
    wire \c0.rx.n19538 ;
    wire \c0.rx.n19539 ;
    wire \c0.rx.n14391 ;
    wire \c0.rx.n17411 ;
    wire \c0.data_out_frame_29_7_N_1483_0 ;
    wire \c0.n1220 ;
    wire \c0.FRAME_MATCHER_i_28 ;
    wire \c0.n31_adj_4271 ;
    wire \c0.n3_adj_4430 ;
    wire \c0.data_in_frame_7_4 ;
    wire \c0.n13555_cascade_ ;
    wire \c0.n13555 ;
    wire \c0.n22043_cascade_ ;
    wire \c0.data_in_frame_2_6 ;
    wire \c0.data_in_frame_0_4 ;
    wire \c0.n10_adj_4363 ;
    wire \c0.n22283 ;
    wire \c0.n13488_cascade_ ;
    wire \c0.n13180 ;
    wire \c0.data_in_frame_0_5 ;
    wire \c0.data_in_frame_0_6 ;
    wire \c0.n23827 ;
    wire \c0.data_in_frame_5_3 ;
    wire \c0.data_in_frame_7_5 ;
    wire \c0.n12484 ;
    wire \c0.n20368_cascade_ ;
    wire \c0.data_in_frame_10_1 ;
    wire \c0.n22133_cascade_ ;
    wire \c0.n21925 ;
    wire \c0.n20927_cascade_ ;
    wire \c0.n22133 ;
    wire \c0.n36 ;
    wire data_in_frame_1_2;
    wire \c0.n22334 ;
    wire \c0.n22334_cascade_ ;
    wire \c0.n22051 ;
    wire \c0.n15_adj_4404 ;
    wire \c0.data_in_frame_8_0 ;
    wire \c0.data_in_frame_7_7 ;
    wire \c0.n6_adj_4259 ;
    wire \c0.n39_adj_4263 ;
    wire \c0.n40_adj_4261 ;
    wire \c0.n22060_cascade_ ;
    wire \c0.n44_adj_4262 ;
    wire \c0.n11_adj_4266_cascade_ ;
    wire \c0.n13425 ;
    wire \c0.n22842_cascade_ ;
    wire \c0.data_in_frame_5_6 ;
    wire \c0.n22245 ;
    wire \c0.n22379 ;
    wire \c0.n38_adj_4260 ;
    wire \c0.n6_adj_4256 ;
    wire \c0.data_in_frame_7_3 ;
    wire \c0.n13488 ;
    wire \c0.n22139_cascade_ ;
    wire \c0.data_in_frame_9_0 ;
    wire \c0.n13605 ;
    wire \c0.n13043 ;
    wire \c0.data_in_frame_8_6 ;
    wire \c0.n21822_cascade_ ;
    wire \c0.n22443 ;
    wire \c0.n10_adj_4242_cascade_ ;
    wire \c0.data_in_frame_8_1 ;
    wire \c0.data_in_frame_16_6 ;
    wire \c0.n13786_cascade_ ;
    wire \c0.n21170 ;
    wire \c0.n13974 ;
    wire \c0.data_in_frame_10_2 ;
    wire \c0.n20402_cascade_ ;
    wire \c0.data_in_frame_9_6 ;
    wire \c0.data_in_frame_9_4 ;
    wire \c0.n21873 ;
    wire \c0.n13287 ;
    wire \c0.n13190 ;
    wire \c0.n18_adj_4222_cascade_ ;
    wire \c0.n22270 ;
    wire \c0.n6_adj_4221 ;
    wire \c0.n22308 ;
    wire \c0.n22003_cascade_ ;
    wire \c0.n5943 ;
    wire \c0.n6221_cascade_ ;
    wire \c0.n22003 ;
    wire \c0.data_in_frame_20_1 ;
    wire \c0.n6_adj_4226_cascade_ ;
    wire \c0.n23615_cascade_ ;
    wire \c0.n22100_cascade_ ;
    wire \c0.n22081 ;
    wire \c0.n6_adj_4224 ;
    wire \c0.n21737 ;
    wire \c0.n6_adj_4353 ;
    wire \c0.n5_adj_4342 ;
    wire \c0.FRAME_MATCHER_state_20 ;
    wire \c0.n21366 ;
    wire \c0.n21855 ;
    wire encoder0_position_2;
    wire \c0.n22248 ;
    wire \c0.n13379 ;
    wire \c0.data_in_frame_20_7 ;
    wire \c0.n28_cascade_ ;
    wire \c0.n23640_cascade_ ;
    wire \c0.n22305_cascade_ ;
    wire \c0.data_in_frame_21_1 ;
    wire \c0.n23640 ;
    wire \c0.n22305 ;
    wire \c0.n6_adj_4219_cascade_ ;
    wire \c0.data_in_frame_21_2 ;
    wire \c0.n22197 ;
    wire \c0.n21949_cascade_ ;
    wire \c0.n20137 ;
    wire \c0.n22157_cascade_ ;
    wire \c0.n20846 ;
    wire \c0.n20846_cascade_ ;
    wire \c0.data_in_frame_25_4 ;
    wire \c0.data_in_frame_25_2 ;
    wire \c0.data_in_frame_25_3 ;
    wire \c0.data_in_frame_25_5 ;
    wire \c0.n22370 ;
    wire \c0.n12_adj_4491 ;
    wire \c0.n23009 ;
    wire \c0.n22370_cascade_ ;
    wire \c0.n23356 ;
    wire \c0.n13761 ;
    wire \c0.n22145 ;
    wire \c0.n21949 ;
    wire \c0.n22145_cascade_ ;
    wire \c0.n10_adj_4297 ;
    wire \c0.n23335_cascade_ ;
    wire \c0.n21_adj_4300 ;
    wire \c0.data_in_frame_29_3 ;
    wire \c0.data_in_frame_28_0 ;
    wire \c0.n6404 ;
    wire \c0.n21834 ;
    wire \c0.n22040 ;
    wire \c0.n22040_cascade_ ;
    wire \c0.n21208 ;
    wire \c0.n21099 ;
    wire \c0.n22119 ;
    wire \c0.n21099_cascade_ ;
    wire \c0.n21160 ;
    wire \c0.data_in_frame_29_6 ;
    wire \c0.n63_adj_4293 ;
    wire \c0.n22148_cascade_ ;
    wire \c0.n21233 ;
    wire \c0.n26_adj_4294 ;
    wire \c0.rx.n12862_cascade_ ;
    wire \c0.rx.r_Clock_Count_7 ;
    wire \c0.rx.r_Clock_Count_5 ;
    wire \c0.rx.r_Clock_Count_6 ;
    wire \c0.rx.n80_cascade_ ;
    wire r_SM_Main_2_N_3681_2_cascade_;
    wire n14283;
    wire \c0.rx.r_Clock_Count_4 ;
    wire \c0.rx.n18655 ;
    wire \c0.rx.r_Clock_Count_0 ;
    wire \c0.rx.n80 ;
    wire \c0.rx.n21783 ;
    wire \c0.rx.r_Rx_Data_R ;
    wire \c0.data_in_frame_12_6 ;
    wire \c0.data_in_frame_15_3 ;
    wire \c0.n20927 ;
    wire \c0.n22060 ;
    wire \c0.n6_adj_4244_cascade_ ;
    wire \c0.n21097 ;
    wire \c0.n20240_cascade_ ;
    wire \c0.data_in_frame_15_0 ;
    wire \c0.n22385_cascade_ ;
    wire data_in_frame_14_5;
    wire data_in_frame_14_3;
    wire \c0.data_in_frame_4_0 ;
    wire data_in_frame_1_4;
    wire \c0.n21797 ;
    wire \c0.n13237 ;
    wire \c0.data_in_frame_7_6 ;
    wire \c0.data_in_frame_10_0 ;
    wire \c0.n10_adj_4245_cascade_ ;
    wire \c0.n13099 ;
    wire \c0.data_in_frame_9_1 ;
    wire \c0.n14037 ;
    wire \c0.n22233 ;
    wire \c0.data_in_frame_11_3 ;
    wire \c0.n10_adj_4274 ;
    wire \c0.n22108 ;
    wire \c0.n4_adj_4240_cascade_ ;
    wire \c0.data_in_frame_7_1 ;
    wire \c0.n6_adj_4273 ;
    wire \c0.n22139 ;
    wire \c0.n6_adj_4243 ;
    wire \c0.n13861 ;
    wire \c0.n5813_cascade_ ;
    wire \c0.n21967 ;
    wire \c0.n20222_cascade_ ;
    wire \c0.n13677 ;
    wire \c0.n28_adj_4232_cascade_ ;
    wire \c0.n32_cascade_ ;
    wire \c0.n29_adj_4234 ;
    wire \c0.n13681 ;
    wire \c0.n21238_cascade_ ;
    wire \c0.n21989 ;
    wire \c0.n21238 ;
    wire \c0.n22430 ;
    wire \c0.n5810 ;
    wire \c0.n13719_cascade_ ;
    wire \c0.n22221 ;
    wire \c0.n13786 ;
    wire data_in_frame_14_6;
    wire data_in_frame_14_7;
    wire \c0.n5996 ;
    wire \c0.n7_adj_4235 ;
    wire \c0.n8_adj_4236 ;
    wire \c0.n20203_cascade_ ;
    wire \c0.n21120 ;
    wire \c0.data_in_frame_15_2 ;
    wire \c0.n22242 ;
    wire \c0.n20402 ;
    wire \c0.n20196 ;
    wire \c0.n22100 ;
    wire \c0.n21054_cascade_ ;
    wire \c0.n21043 ;
    wire \c0.data_in_frame_17_3 ;
    wire \c0.data_in_frame_17_4 ;
    wire \c0.n22480 ;
    wire \c0.data_in_frame_17_5 ;
    wire \c0.n13719 ;
    wire \c0.n18 ;
    wire \c0.n22349 ;
    wire \c0.n30 ;
    wire \c0.n22 ;
    wire \c0.n22355 ;
    wire \c0.n23062_cascade_ ;
    wire \c0.data_in_frame_21_0 ;
    wire \c0.n23062 ;
    wire \c0.n8 ;
    wire \c0.n27 ;
    wire \c0.n22296 ;
    wire \c0.n21831 ;
    wire \c0.data_in_frame_17_0 ;
    wire \c0.n16_adj_4223_cascade_ ;
    wire \c0.n17 ;
    wire \c0.n21187 ;
    wire \c0.n22211_cascade_ ;
    wire \c0.n21140 ;
    wire \c0.n22311 ;
    wire \c0.n22211 ;
    wire \c0.n23298 ;
    wire \c0.n7 ;
    wire \c0.n23298_cascade_ ;
    wire \c0.n45_adj_4486 ;
    wire \c0.data_in_frame_27_4 ;
    wire \c0.n52_cascade_ ;
    wire \c0.n13872 ;
    wire \c0.n12420 ;
    wire \c0.n23615 ;
    wire \c0.n44_adj_4490 ;
    wire \c0.n48_adj_4485_cascade_ ;
    wire \c0.n12_adj_4290 ;
    wire \c0.data_in_frame_25_1 ;
    wire \c0.n49_adj_4488 ;
    wire \c0.n55 ;
    wire \c0.n53 ;
    wire \c0.n23416 ;
    wire \c0.n23416_cascade_ ;
    wire \c0.n12_adj_4296 ;
    wire \c0.data_in_frame_27_2 ;
    wire \c0.n36_adj_4489 ;
    wire \c0.data_in_frame_19_2 ;
    wire \c0.n6221 ;
    wire \c0.n21037 ;
    wire \c0.data_in_frame_23_6 ;
    wire \c0.n21037_cascade_ ;
    wire \c0.data_in_frame_19_4 ;
    wire \c0.n13282 ;
    wire \c0.n20370 ;
    wire \c0.data_in_frame_29_5 ;
    wire \c0.n22157 ;
    wire \c0.data_in_frame_27_3 ;
    wire \c0.n22719 ;
    wire \c0.n8_adj_4291_cascade_ ;
    wire \c0.n22148 ;
    wire \c0.n23811 ;
    wire n12977;
    wire \c0.rx.n21704 ;
    wire n14436_cascade_;
    wire \c0.rx.n12862 ;
    wire n19619;
    wire r_Bit_Index_2;
    wire n91_cascade_;
    wire r_SM_Main_2_N_3681_2;
    wire r_SM_Main_2;
    wire r_SM_Main_1;
    wire \c0.rx.n14_cascade_ ;
    wire \c0.rx.n36 ;
    wire r_SM_Main_0;
    wire n21755_cascade_;
    wire data_in_frame_14_1;
    wire \c0.FRAME_MATCHER_i_0 ;
    wire \c0.FRAME_MATCHER_i_1 ;
    wire \c0.FRAME_MATCHER_i_2 ;
    wire \c0.n22043 ;
    wire \c0.data_in_frame_9_7 ;
    wire \c0.n22471 ;
    wire \c0.data_in_frame_16_4 ;
    wire \c0.n20240 ;
    wire \c0.n22446 ;
    wire \c0.n22328 ;
    wire \c0.n22446_cascade_ ;
    wire \c0.n22424 ;
    wire \c0.n30_adj_4233 ;
    wire data_in_frame_14_2;
    wire \c0.n22340 ;
    wire n21755;
    wire data_in_frame_14_4;
    wire \c0.n15_adj_4269 ;
    wire \c0.n22464_cascade_ ;
    wire \c0.n22415 ;
    wire \c0.n13728 ;
    wire \c0.n14053 ;
    wire \c0.data_in_frame_18_1 ;
    wire \c0.n14053_cascade_ ;
    wire \c0.data_in_frame_17_7 ;
    wire \c0.n23586_cascade_ ;
    wire \c0.data_in_frame_9_3 ;
    wire \c0.n13210_cascade_ ;
    wire \c0.data_in_frame_8_7 ;
    wire \c0.n21822 ;
    wire \c0.n7_adj_4277_cascade_ ;
    wire \c0.data_in_frame_11_5 ;
    wire \c0.n10_adj_4264_cascade_ ;
    wire \c0.n16_adj_4265 ;
    wire \c0.data_in_frame_11_6 ;
    wire \c0.data_in_frame_11_2 ;
    wire \c0.n20135 ;
    wire \c0.n22464 ;
    wire \c0.n21867 ;
    wire \c0.n6_adj_4225 ;
    wire \c0.n21982 ;
    wire data_in_frame_14_0;
    wire \c0.n13865 ;
    wire \c0.data_in_frame_15_6 ;
    wire \c0.n4_adj_4240 ;
    wire \c0.n22352_cascade_ ;
    wire \c0.n22000_cascade_ ;
    wire \c0.n31 ;
    wire \c0.data_in_frame_15_7 ;
    wire \c0.data_in_frame_18_2 ;
    wire \c0.n22000 ;
    wire \c0.n12_cascade_ ;
    wire \c0.n10_adj_4239 ;
    wire \c0.data_in_frame_18_0 ;
    wire \c0.n14_adj_4238 ;
    wire \c0.n22352 ;
    wire \c0.data_in_frame_18_4 ;
    wire \c0.n13598 ;
    wire \c0.n20374 ;
    wire \c0.data_in_frame_16_5 ;
    wire \c0.data_in_frame_16_3 ;
    wire \c0.data_in_frame_16_2 ;
    wire \c0.n10_adj_4230 ;
    wire \c0.data_in_frame_13_4 ;
    wire \c0.data_in_frame_15_5 ;
    wire \c0.data_in_frame_26_3 ;
    wire \c0.n20266 ;
    wire \c0.n22402_cascade_ ;
    wire \c0.n33 ;
    wire \c0.n21054 ;
    wire \c0.n6_adj_4292_cascade_ ;
    wire \c0.data_in_frame_28_5 ;
    wire \c0.n23073 ;
    wire \c0.data_in_frame_21_4 ;
    wire \c0.n21905 ;
    wire \c0.n21905_cascade_ ;
    wire \c0.n21069 ;
    wire \c0.n22113 ;
    wire \c0.data_in_frame_20_3 ;
    wire \c0.n20203 ;
    wire \c0.n21870 ;
    wire \c0.n18_adj_4249_cascade_ ;
    wire \c0.n24_adj_4248 ;
    wire \c0.n26_adj_4250 ;
    wire \c0.data_in_frame_15_4 ;
    wire \c0.n23072 ;
    wire \c0.n13457 ;
    wire \c0.n23072_cascade_ ;
    wire \c0.n21067 ;
    wire \c0.n14_adj_4251 ;
    wire \c0.data_in_frame_19_5 ;
    wire \c0.data_in_frame_26_1 ;
    wire \c0.n21039 ;
    wire \c0.n24_adj_4282_cascade_ ;
    wire \c0.n22711 ;
    wire \c0.n22711_cascade_ ;
    wire \c0.n21200 ;
    wire \c0.n12596 ;
    wire \c0.n6707 ;
    wire \c0.n15_adj_4284_cascade_ ;
    wire \c0.n14_adj_4283 ;
    wire \c0.n22437 ;
    wire \c0.data_in_frame_25_0 ;
    wire \c0.data_in_frame_25_6 ;
    wire \c0.n22437_cascade_ ;
    wire \c0.n50_adj_4487 ;
    wire \c0.n22323 ;
    wire \c0.n10_adj_4483 ;
    wire \c0.n20537_cascade_ ;
    wire \c0.n14_adj_4484 ;
    wire \c0.n21890 ;
    wire \c0.n21087 ;
    wire \c0.n13320_cascade_ ;
    wire \c0.n22468 ;
    wire \c0.n10_cascade_ ;
    wire \c0.n20537 ;
    wire \c0.n22314 ;
    wire \c0.data_in_frame_24_3 ;
    wire \c0.n22142 ;
    wire \c0.data_in_frame_24_4 ;
    wire \c0.n22028 ;
    wire \c0.n22337_cascade_ ;
    wire \c0.n22020 ;
    wire \c0.n21095 ;
    wire \c0.n6_adj_4418 ;
    wire \c0.data_in_frame_26_4 ;
    wire \c0.n22337 ;
    wire \c0.n10_adj_4285_cascade_ ;
    wire \c0.n22995 ;
    wire \c0.data_in_frame_26_6 ;
    wire \c0.n22054 ;
    wire \c0.data_in_frame_24_6 ;
    wire \c0.n22434 ;
    wire \c0.data_in_frame_20_0 ;
    wire data_in_frame_22_2;
    wire \c0.n12594 ;
    wire \c0.n20596 ;
    wire \c0.data_in_frame_11_7 ;
    wire n21760;
    wire \c0.data_in_frame_26_2 ;
    wire \c0.n13993 ;
    wire n91;
    wire n12973;
    wire n14917;
    wire n14436;
    wire r_Bit_Index_1;
    wire data_in_frame_22_4;
    wire \c0.n22191 ;
    wire \c0.n25 ;
    wire r_Bit_Index_0;
    wire r_Rx_Data;
    wire n12970;
    wire \c0.data_in_frame_12_0 ;
    wire \c0.data_in_frame_24_7 ;
    wire \c0.data_in_frame_12_1 ;
    wire \c0.data_in_frame_12_2 ;
    wire \c0.data_in_frame_13_2 ;
    wire \c0.data_in_frame_13_1 ;
    wire \c0.data_in_frame_11_0 ;
    wire \c0.n22274 ;
    wire \c0.data_in_frame_10_6 ;
    wire \c0.n13999_cascade_ ;
    wire \c0.n21940 ;
    wire \c0.n13233 ;
    wire \c0.data_in_frame_9_2 ;
    wire \c0.n21845 ;
    wire \c0.n22781 ;
    wire \c0.data_in_frame_11_1 ;
    wire \c0.data_in_frame_23_3 ;
    wire \c0.n22236 ;
    wire \c0.n4 ;
    wire \c0.n5965 ;
    wire \c0.n8_adj_4275 ;
    wire \c0.n8_adj_4276 ;
    wire \c0.data_in_frame_13_0 ;
    wire \c0.data_in_frame_12_7 ;
    wire \c0.data_in_frame_23_1 ;
    wire data_in_frame_22_7;
    wire \c0.n21995 ;
    wire \c0.data_in_frame_21_7 ;
    wire \c0.n13210 ;
    wire \c0.n22091 ;
    wire \c0.n21934 ;
    wire \c0.data_in_frame_4_5 ;
    wire \c0.n13421 ;
    wire \c0.data_in_frame_11_4 ;
    wire \c0.n13421_cascade_ ;
    wire \c0.n22069 ;
    wire \c0.n10_adj_4252 ;
    wire \c0.data_in_frame_7_2 ;
    wire \c0.n22343 ;
    wire \c0.n10_adj_4267 ;
    wire \c0.data_in_frame_12_5 ;
    wire \c0.n16_adj_4268 ;
    wire \c0.n21740 ;
    wire \c0.data_in_frame_7_0 ;
    wire \c0.data_in_frame_16_1 ;
    wire \c0.data_in_frame_12_3 ;
    wire \c0.n21975 ;
    wire \c0.data_in_frame_17_2 ;
    wire \c0.data_in_frame_15_1 ;
    wire \c0.data_in_frame_12_4 ;
    wire \c0.data_in_frame_13_3 ;
    wire \c0.data_in_frame_13_5 ;
    wire \c0.n14081 ;
    wire \c0.data_in_frame_16_0 ;
    wire \c0.data_in_frame_20_4 ;
    wire data_in_frame_22_6;
    wire \c0.n20246 ;
    wire \c0.data_in_frame_13_6 ;
    wire \c0.data_in_frame_26_5 ;
    wire \c0.data_in_frame_21_6 ;
    wire \c0.n21749 ;
    wire \c0.n9_adj_4237 ;
    wire \c0.data_in_frame_13_7 ;
    wire \c0.n22388 ;
    wire \c0.data_in_frame_17_6 ;
    wire \c0.n20_adj_4247 ;
    wire \c0.data_in_frame_20_2 ;
    wire \c0.n13544 ;
    wire data_in_frame_22_3;
    wire \c0.n23426 ;
    wire \c0.n22007 ;
    wire \c0.data_in_frame_19_6 ;
    wire \c0.data_in_frame_18_5 ;
    wire \c0.n22385 ;
    wire \c0.n21126 ;
    wire \c0.data_in_frame_19_1 ;
    wire \c0.n22084 ;
    wire \c0.n22364 ;
    wire \c0.data_in_frame_19_7 ;
    wire \c0.n15 ;
    wire \c0.data_in_frame_20_5 ;
    wire \c0.data_in_frame_23_0 ;
    wire \c0.n26_adj_4281 ;
    wire rx_data_4;
    wire \c0.data_in_frame_18_3 ;
    wire \c0.n22095 ;
    wire \c0.n21124 ;
    wire \c0.n22095_cascade_ ;
    wire \c0.n14143 ;
    wire \c0.n29 ;
    wire data_in_frame_22_0;
    wire \c0.n22267 ;
    wire \c0.n22105 ;
    wire \c0.n22849 ;
    wire \c0.n20406 ;
    wire \c0.n5813 ;
    wire \c0.n21864 ;
    wire \c0.n13768 ;
    wire \c0.n22458 ;
    wire \c0.n21114 ;
    wire \c0.n18_adj_4246 ;
    wire \c0.n21_cascade_ ;
    wire \c0.n22399 ;
    wire \c0.n24 ;
    wire \c0.n20 ;
    wire \c0.data_in_frame_17_1 ;
    wire \c0.n16 ;
    wire \c0.n21979 ;
    wire \c0.n23287 ;
    wire \c0.n23287_cascade_ ;
    wire \c0.data_in_frame_19_3 ;
    wire \c0.n21921 ;
    wire rx_data_1;
    wire \c0.data_in_frame_24_0 ;
    wire \c0.data_in_frame_24_5 ;
    wire \c0.n13320 ;
    wire data_in_frame_22_5;
    wire \c0.n22255 ;
    wire \c0.data_in_frame_23_7 ;
    wire \c0.n22396 ;
    wire \c0.n20288 ;
    wire \c0.n23 ;
    wire \c0.data_in_frame_24_2 ;
    wire \c0.n13443 ;
    wire \c0.n22358 ;
    wire \c0.n22099 ;
    wire \c0.data_in_frame_24_1 ;
    wire \c0.n22057 ;
    wire \c0.n22373 ;
    wire \c0.n8_adj_4288_cascade_ ;
    wire \c0.n24_adj_4289 ;
    wire \c0.n22215 ;
    wire \c0.n22402 ;
    wire \c0.data_in_frame_28_4 ;
    wire \c0.n22455 ;
    wire \c0.n22997 ;
    wire rx_data_3;
    wire \c0.data_in_frame_28_3 ;
    wire \c0.data_in_frame_28_7 ;
    wire \c0.n9_adj_4217 ;
    wire \c0.data_in_frame_28_6 ;
    wire \c0.data_in_frame_27_7 ;
    wire \c0.data_in_frame_27_6 ;
    wire \c0.data_in_frame_27_0 ;
    wire \c0.n6268 ;
    wire \c0.n9_adj_4278 ;
    wire \c0.data_in_frame_16_7 ;
    wire \c0.data_in_frame_19_0 ;
    wire rx_data_6;
    wire \c0.data_in_frame_18_6 ;
    wire \c0.data_in_frame_18_7 ;
    wire \c0.data_in_frame_21_5 ;
    wire \c0.n22123 ;
    wire \c0.n9_adj_4302 ;
    wire \c0.data_in_frame_25_7 ;
    wire rx_data_0;
    wire \c0.data_in_frame_26_0 ;
    wire \c0.n9_adj_4341 ;
    wire rx_data_7;
    wire \c0.data_in_frame_26_7 ;
    wire \c0.n17596 ;
    wire rx_data_2;
    wire \c0.n21758 ;
    wire \c0.data_in_frame_23_2 ;
    wire \c0.n21775 ;
    wire \c0.n9 ;
    wire rx_data_5;
    wire \c0.data_in_frame_27_5 ;
    wire PIN_9_c;
    wire _gnd_net_;

    defparam \pll32MHz_inst.pll20MHz_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll32MHz_inst.pll20MHz_inst .TEST_MODE=1'b0;
    defparam \pll32MHz_inst.pll20MHz_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll32MHz_inst.pll20MHz_inst .PLLOUT_SELECT="SHIFTREG_0deg";
    defparam \pll32MHz_inst.pll20MHz_inst .FILTER_RANGE=3'b001;
    defparam \pll32MHz_inst.pll20MHz_inst .FEEDBACK_PATH="PHASE_AND_DELAY";
    defparam \pll32MHz_inst.pll20MHz_inst .FDA_RELATIVE=4'b0000;
    defparam \pll32MHz_inst.pll20MHz_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll32MHz_inst.pll20MHz_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll32MHz_inst.pll20MHz_inst .DIVR=4'b0000;
    defparam \pll32MHz_inst.pll20MHz_inst .DIVQ=3'b011;
    defparam \pll32MHz_inst.pll20MHz_inst .DIVF=7'b0000001;
    defparam \pll32MHz_inst.pll20MHz_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll32MHz_inst.pll20MHz_inst  (
            .BYPASS(GNDG0),
            .DYNAMICDELAY({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7}),
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .LOCK(),
            .PLLOUTCORE(),
            .PLLOUTGLOBAL(PIN_9_c),
            .REFERENCECLK(N__23719),
            .RESETB(N__47218),
            .SCLK(),
            .SDI(),
            .SDO());
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__70064),
            .DIN(N__70063),
            .DOUT(N__70062),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__70064),
            .PADOUT(N__70063),
            .PADIN(N__70062),
            .CLOCKENABLE(),
            .DIN0(CLK_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__70055),
            .DIN(N__70054),
            .DOUT(N__70053),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__70055),
            .PADOUT(N__70054),
            .PADIN(N__70053),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__23683),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_12_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_12_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_12_pad_iopad (
            .OE(N__70046),
            .DIN(N__70045),
            .DOUT(N__70044),
            .PACKAGEPIN(PIN_12));
    defparam PIN_12_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_12_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_12_pad_preio (
            .PADOEN(N__70046),
            .PADOUT(N__70045),
            .PADIN(N__70044),
            .CLOCKENABLE(),
            .DIN0(PIN_12_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_13_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_13_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_13_pad_iopad (
            .OE(N__70037),
            .DIN(N__70036),
            .DOUT(N__70035),
            .PACKAGEPIN(PIN_13));
    defparam PIN_13_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_13_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_13_pad_preio (
            .PADOEN(N__70037),
            .PADOUT(N__70036),
            .PADIN(N__70035),
            .CLOCKENABLE(),
            .DIN0(PIN_13_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_1_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_1_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_1_pad_iopad (
            .OE(N__70028),
            .DIN(N__70027),
            .DOUT(N__70026),
            .PACKAGEPIN(PIN_1));
    defparam PIN_1_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_1_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_1_pad_preio (
            .PADOEN(N__70028),
            .PADOUT(N__70027),
            .PADIN(N__70026),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_22_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_22_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_22_pad_iopad (
            .OE(N__70019),
            .DIN(N__70018),
            .DOUT(N__70017),
            .PACKAGEPIN(PIN_22));
    defparam PIN_22_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_22_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_22_pad_preio (
            .PADOEN(N__70019),
            .PADOUT(N__70018),
            .PADIN(N__70017),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_23_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_23_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_23_pad_iopad (
            .OE(N__70010),
            .DIN(N__70009),
            .DOUT(N__70008),
            .PACKAGEPIN(PIN_23));
    defparam PIN_23_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_23_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_23_pad_preio (
            .PADOEN(N__70010),
            .PADOUT(N__70009),
            .PADIN(N__70008),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_24_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_24_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_24_pad_iopad (
            .OE(N__70001),
            .DIN(N__70000),
            .DOUT(N__69999),
            .PACKAGEPIN(PIN_24));
    defparam PIN_24_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_24_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_24_pad_preio (
            .PADOEN(N__70001),
            .PADOUT(N__70000),
            .PADIN(N__69999),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_2_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_2_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_2_pad_iopad (
            .OE(N__69992),
            .DIN(N__69991),
            .DOUT(N__69990),
            .PACKAGEPIN(PIN_2));
    defparam PIN_2_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_2_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_2_pad_preio (
            .PADOEN(N__69992),
            .PADOUT(N__69991),
            .PADIN(N__69990),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_3_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_3_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_3_pad_iopad (
            .OE(N__69983),
            .DIN(N__69982),
            .DOUT(N__69981),
            .PACKAGEPIN(PIN_3));
    defparam PIN_3_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_3_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_3_pad_preio (
            .PADOEN(N__69983),
            .PADOUT(N__69982),
            .PADIN(N__69981),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_7_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_7_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_7_pad_iopad (
            .OE(N__69974),
            .DIN(N__69973),
            .DOUT(N__69972),
            .PACKAGEPIN(PIN_7));
    defparam PIN_7_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_7_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_7_pad_preio (
            .PADOEN(N__69974),
            .PADOUT(N__69973),
            .PADIN(N__69972),
            .CLOCKENABLE(),
            .DIN0(PIN_7_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_8_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_8_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_8_pad_iopad (
            .OE(N__69965),
            .DIN(N__69964),
            .DOUT(N__69963),
            .PACKAGEPIN(PIN_8));
    defparam PIN_8_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_8_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_8_pad_preio (
            .PADOEN(N__69965),
            .PADOUT(N__69964),
            .PADIN(N__69963),
            .CLOCKENABLE(),
            .DIN0(PIN_8_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_9_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_9_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_9_pad_iopad (
            .OE(N__69956),
            .DIN(N__69955),
            .DOUT(N__69954),
            .PACKAGEPIN(PIN_9));
    defparam PIN_9_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_9_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_9_pad_preio (
            .PADOEN(N__69956),
            .PADOUT(N__69955),
            .PADIN(N__69954),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__23689),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__69947),
            .DIN(N__69946),
            .DOUT(N__69945),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__69947),
            .PADOUT(N__69946),
            .PADIN(N__69945),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall1_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall1_input_iopad.PULLUP=1'b1;
    IO_PAD hall1_input_iopad (
            .OE(N__69938),
            .DIN(N__69937),
            .DOUT(N__69936),
            .PACKAGEPIN(PIN_4));
    defparam hall1_input_preio.PIN_TYPE=6'b000001;
    defparam hall1_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall1_input_preio (
            .PADOEN(N__69938),
            .PADOUT(N__69937),
            .PADIN(N__69936),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall2_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall2_input_iopad.PULLUP=1'b1;
    IO_PAD hall2_input_iopad (
            .OE(N__69929),
            .DIN(N__69928),
            .DOUT(N__69927),
            .PACKAGEPIN(PIN_5));
    defparam hall2_input_preio.PIN_TYPE=6'b000001;
    defparam hall2_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall2_input_preio (
            .PADOEN(N__69929),
            .PADOUT(N__69928),
            .PADIN(N__69927),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall3_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall3_input_iopad.PULLUP=1'b1;
    IO_PAD hall3_input_iopad (
            .OE(N__69920),
            .DIN(N__69919),
            .DOUT(N__69918),
            .PACKAGEPIN(PIN_6));
    defparam hall3_input_preio.PIN_TYPE=6'b000001;
    defparam hall3_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall3_input_preio (
            .PADOEN(N__69920),
            .PADOUT(N__69919),
            .PADIN(N__69918),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rx_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_input_iopad.PULLUP=1'b1;
    IO_PAD rx_input_iopad (
            .OE(N__69911),
            .DIN(N__69910),
            .DOUT(N__69909),
            .PACKAGEPIN(PIN_11));
    defparam rx_input_preio.PIN_TYPE=6'b000001;
    defparam rx_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_input_preio (
            .PADOEN(N__69911),
            .PADOUT(N__69910),
            .PADIN(N__69909),
            .CLOCKENABLE(),
            .DIN0(rx_i),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam tx_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_output_iopad.PULLUP=1'b1;
    IO_PAD tx_output_iopad (
            .OE(N__69902),
            .DIN(N__69901),
            .DOUT(N__69900),
            .PACKAGEPIN(PIN_10));
    defparam tx_output_preio.PIN_TYPE=6'b101001;
    defparam tx_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_output_preio (
            .PADOEN(N__69902),
            .PADOUT(N__69901),
            .PADIN(N__69900),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__26524),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__23695));
    InMux I__17391 (
            .O(N__69883),
            .I(N__69873));
    CascadeMux I__17390 (
            .O(N__69882),
            .I(N__69868));
    CascadeMux I__17389 (
            .O(N__69881),
            .I(N__69861));
    InMux I__17388 (
            .O(N__69880),
            .I(N__69857));
    InMux I__17387 (
            .O(N__69879),
            .I(N__69854));
    CascadeMux I__17386 (
            .O(N__69878),
            .I(N__69851));
    CascadeMux I__17385 (
            .O(N__69877),
            .I(N__69848));
    CascadeMux I__17384 (
            .O(N__69876),
            .I(N__69841));
    LocalMux I__17383 (
            .O(N__69873),
            .I(N__69836));
    InMux I__17382 (
            .O(N__69872),
            .I(N__69833));
    InMux I__17381 (
            .O(N__69871),
            .I(N__69830));
    InMux I__17380 (
            .O(N__69868),
            .I(N__69827));
    InMux I__17379 (
            .O(N__69867),
            .I(N__69824));
    CascadeMux I__17378 (
            .O(N__69866),
            .I(N__69821));
    InMux I__17377 (
            .O(N__69865),
            .I(N__69818));
    InMux I__17376 (
            .O(N__69864),
            .I(N__69815));
    InMux I__17375 (
            .O(N__69861),
            .I(N__69810));
    InMux I__17374 (
            .O(N__69860),
            .I(N__69810));
    LocalMux I__17373 (
            .O(N__69857),
            .I(N__69807));
    LocalMux I__17372 (
            .O(N__69854),
            .I(N__69803));
    InMux I__17371 (
            .O(N__69851),
            .I(N__69798));
    InMux I__17370 (
            .O(N__69848),
            .I(N__69795));
    InMux I__17369 (
            .O(N__69847),
            .I(N__69791));
    InMux I__17368 (
            .O(N__69846),
            .I(N__69784));
    InMux I__17367 (
            .O(N__69845),
            .I(N__69784));
    InMux I__17366 (
            .O(N__69844),
            .I(N__69784));
    InMux I__17365 (
            .O(N__69841),
            .I(N__69781));
    InMux I__17364 (
            .O(N__69840),
            .I(N__69778));
    InMux I__17363 (
            .O(N__69839),
            .I(N__69774));
    Span4Mux_v I__17362 (
            .O(N__69836),
            .I(N__69771));
    LocalMux I__17361 (
            .O(N__69833),
            .I(N__69766));
    LocalMux I__17360 (
            .O(N__69830),
            .I(N__69766));
    LocalMux I__17359 (
            .O(N__69827),
            .I(N__69761));
    LocalMux I__17358 (
            .O(N__69824),
            .I(N__69761));
    InMux I__17357 (
            .O(N__69821),
            .I(N__69758));
    LocalMux I__17356 (
            .O(N__69818),
            .I(N__69751));
    LocalMux I__17355 (
            .O(N__69815),
            .I(N__69751));
    LocalMux I__17354 (
            .O(N__69810),
            .I(N__69751));
    Span4Mux_h I__17353 (
            .O(N__69807),
            .I(N__69747));
    InMux I__17352 (
            .O(N__69806),
            .I(N__69744));
    Span4Mux_v I__17351 (
            .O(N__69803),
            .I(N__69741));
    InMux I__17350 (
            .O(N__69802),
            .I(N__69736));
    InMux I__17349 (
            .O(N__69801),
            .I(N__69736));
    LocalMux I__17348 (
            .O(N__69798),
            .I(N__69731));
    LocalMux I__17347 (
            .O(N__69795),
            .I(N__69731));
    CascadeMux I__17346 (
            .O(N__69794),
            .I(N__69727));
    LocalMux I__17345 (
            .O(N__69791),
            .I(N__69720));
    LocalMux I__17344 (
            .O(N__69784),
            .I(N__69720));
    LocalMux I__17343 (
            .O(N__69781),
            .I(N__69720));
    LocalMux I__17342 (
            .O(N__69778),
            .I(N__69717));
    CascadeMux I__17341 (
            .O(N__69777),
            .I(N__69713));
    LocalMux I__17340 (
            .O(N__69774),
            .I(N__69710));
    Span4Mux_h I__17339 (
            .O(N__69771),
            .I(N__69703));
    Span4Mux_v I__17338 (
            .O(N__69766),
            .I(N__69703));
    Span4Mux_v I__17337 (
            .O(N__69761),
            .I(N__69703));
    LocalMux I__17336 (
            .O(N__69758),
            .I(N__69698));
    Span4Mux_v I__17335 (
            .O(N__69751),
            .I(N__69698));
    InMux I__17334 (
            .O(N__69750),
            .I(N__69692));
    Span4Mux_h I__17333 (
            .O(N__69747),
            .I(N__69687));
    LocalMux I__17332 (
            .O(N__69744),
            .I(N__69687));
    Span4Mux_h I__17331 (
            .O(N__69741),
            .I(N__69680));
    LocalMux I__17330 (
            .O(N__69736),
            .I(N__69680));
    Span4Mux_h I__17329 (
            .O(N__69731),
            .I(N__69680));
    InMux I__17328 (
            .O(N__69730),
            .I(N__69677));
    InMux I__17327 (
            .O(N__69727),
            .I(N__69674));
    Span4Mux_v I__17326 (
            .O(N__69720),
            .I(N__69669));
    Span4Mux_v I__17325 (
            .O(N__69717),
            .I(N__69669));
    InMux I__17324 (
            .O(N__69716),
            .I(N__69666));
    InMux I__17323 (
            .O(N__69713),
            .I(N__69663));
    Span4Mux_h I__17322 (
            .O(N__69710),
            .I(N__69656));
    Span4Mux_h I__17321 (
            .O(N__69703),
            .I(N__69656));
    Span4Mux_v I__17320 (
            .O(N__69698),
            .I(N__69656));
    InMux I__17319 (
            .O(N__69697),
            .I(N__69649));
    InMux I__17318 (
            .O(N__69696),
            .I(N__69649));
    InMux I__17317 (
            .O(N__69695),
            .I(N__69649));
    LocalMux I__17316 (
            .O(N__69692),
            .I(N__69646));
    Span4Mux_v I__17315 (
            .O(N__69687),
            .I(N__69641));
    Span4Mux_v I__17314 (
            .O(N__69680),
            .I(N__69641));
    LocalMux I__17313 (
            .O(N__69677),
            .I(N__69638));
    LocalMux I__17312 (
            .O(N__69674),
            .I(N__69633));
    Span4Mux_v I__17311 (
            .O(N__69669),
            .I(N__69633));
    LocalMux I__17310 (
            .O(N__69666),
            .I(N__69630));
    LocalMux I__17309 (
            .O(N__69663),
            .I(N__69625));
    Span4Mux_v I__17308 (
            .O(N__69656),
            .I(N__69625));
    LocalMux I__17307 (
            .O(N__69649),
            .I(N__69616));
    Sp12to4 I__17306 (
            .O(N__69646),
            .I(N__69616));
    Sp12to4 I__17305 (
            .O(N__69641),
            .I(N__69616));
    Span12Mux_v I__17304 (
            .O(N__69638),
            .I(N__69616));
    Span4Mux_v I__17303 (
            .O(N__69633),
            .I(N__69613));
    Span4Mux_v I__17302 (
            .O(N__69630),
            .I(N__69608));
    Span4Mux_v I__17301 (
            .O(N__69625),
            .I(N__69608));
    Span12Mux_v I__17300 (
            .O(N__69616),
            .I(N__69605));
    Span4Mux_v I__17299 (
            .O(N__69613),
            .I(N__69602));
    Odrv4 I__17298 (
            .O(N__69608),
            .I(\c0.n9_adj_4302 ));
    Odrv12 I__17297 (
            .O(N__69605),
            .I(\c0.n9_adj_4302 ));
    Odrv4 I__17296 (
            .O(N__69602),
            .I(\c0.n9_adj_4302 ));
    InMux I__17295 (
            .O(N__69595),
            .I(N__69591));
    CascadeMux I__17294 (
            .O(N__69594),
            .I(N__69588));
    LocalMux I__17293 (
            .O(N__69591),
            .I(N__69585));
    InMux I__17292 (
            .O(N__69588),
            .I(N__69581));
    Span4Mux_v I__17291 (
            .O(N__69585),
            .I(N__69578));
    InMux I__17290 (
            .O(N__69584),
            .I(N__69575));
    LocalMux I__17289 (
            .O(N__69581),
            .I(\c0.data_in_frame_25_7 ));
    Odrv4 I__17288 (
            .O(N__69578),
            .I(\c0.data_in_frame_25_7 ));
    LocalMux I__17287 (
            .O(N__69575),
            .I(\c0.data_in_frame_25_7 ));
    InMux I__17286 (
            .O(N__69568),
            .I(N__69552));
    InMux I__17285 (
            .O(N__69567),
            .I(N__69549));
    InMux I__17284 (
            .O(N__69566),
            .I(N__69545));
    InMux I__17283 (
            .O(N__69565),
            .I(N__69542));
    InMux I__17282 (
            .O(N__69564),
            .I(N__69539));
    InMux I__17281 (
            .O(N__69563),
            .I(N__69534));
    InMux I__17280 (
            .O(N__69562),
            .I(N__69529));
    InMux I__17279 (
            .O(N__69561),
            .I(N__69529));
    InMux I__17278 (
            .O(N__69560),
            .I(N__69526));
    InMux I__17277 (
            .O(N__69559),
            .I(N__69521));
    InMux I__17276 (
            .O(N__69558),
            .I(N__69521));
    InMux I__17275 (
            .O(N__69557),
            .I(N__69518));
    InMux I__17274 (
            .O(N__69556),
            .I(N__69513));
    InMux I__17273 (
            .O(N__69555),
            .I(N__69513));
    LocalMux I__17272 (
            .O(N__69552),
            .I(N__69510));
    LocalMux I__17271 (
            .O(N__69549),
            .I(N__69507));
    InMux I__17270 (
            .O(N__69548),
            .I(N__69504));
    LocalMux I__17269 (
            .O(N__69545),
            .I(N__69497));
    LocalMux I__17268 (
            .O(N__69542),
            .I(N__69497));
    LocalMux I__17267 (
            .O(N__69539),
            .I(N__69494));
    InMux I__17266 (
            .O(N__69538),
            .I(N__69488));
    InMux I__17265 (
            .O(N__69537),
            .I(N__69483));
    LocalMux I__17264 (
            .O(N__69534),
            .I(N__69477));
    LocalMux I__17263 (
            .O(N__69529),
            .I(N__69474));
    LocalMux I__17262 (
            .O(N__69526),
            .I(N__69471));
    LocalMux I__17261 (
            .O(N__69521),
            .I(N__69468));
    LocalMux I__17260 (
            .O(N__69518),
            .I(N__69465));
    LocalMux I__17259 (
            .O(N__69513),
            .I(N__69456));
    Span4Mux_h I__17258 (
            .O(N__69510),
            .I(N__69456));
    Span4Mux_v I__17257 (
            .O(N__69507),
            .I(N__69456));
    LocalMux I__17256 (
            .O(N__69504),
            .I(N__69456));
    InMux I__17255 (
            .O(N__69503),
            .I(N__69453));
    InMux I__17254 (
            .O(N__69502),
            .I(N__69447));
    Span4Mux_v I__17253 (
            .O(N__69497),
            .I(N__69442));
    Span4Mux_h I__17252 (
            .O(N__69494),
            .I(N__69442));
    InMux I__17251 (
            .O(N__69493),
            .I(N__69439));
    InMux I__17250 (
            .O(N__69492),
            .I(N__69436));
    InMux I__17249 (
            .O(N__69491),
            .I(N__69433));
    LocalMux I__17248 (
            .O(N__69488),
            .I(N__69430));
    InMux I__17247 (
            .O(N__69487),
            .I(N__69427));
    InMux I__17246 (
            .O(N__69486),
            .I(N__69424));
    LocalMux I__17245 (
            .O(N__69483),
            .I(N__69421));
    InMux I__17244 (
            .O(N__69482),
            .I(N__69418));
    InMux I__17243 (
            .O(N__69481),
            .I(N__69413));
    InMux I__17242 (
            .O(N__69480),
            .I(N__69413));
    Span4Mux_h I__17241 (
            .O(N__69477),
            .I(N__69410));
    Span4Mux_h I__17240 (
            .O(N__69474),
            .I(N__69405));
    Span4Mux_v I__17239 (
            .O(N__69471),
            .I(N__69405));
    Span4Mux_v I__17238 (
            .O(N__69468),
            .I(N__69400));
    Span4Mux_h I__17237 (
            .O(N__69465),
            .I(N__69400));
    Span4Mux_h I__17236 (
            .O(N__69456),
            .I(N__69397));
    LocalMux I__17235 (
            .O(N__69453),
            .I(N__69394));
    InMux I__17234 (
            .O(N__69452),
            .I(N__69391));
    InMux I__17233 (
            .O(N__69451),
            .I(N__69388));
    InMux I__17232 (
            .O(N__69450),
            .I(N__69385));
    LocalMux I__17231 (
            .O(N__69447),
            .I(N__69376));
    Span4Mux_h I__17230 (
            .O(N__69442),
            .I(N__69376));
    LocalMux I__17229 (
            .O(N__69439),
            .I(N__69376));
    LocalMux I__17228 (
            .O(N__69436),
            .I(N__69376));
    LocalMux I__17227 (
            .O(N__69433),
            .I(N__69371));
    Span4Mux_h I__17226 (
            .O(N__69430),
            .I(N__69368));
    LocalMux I__17225 (
            .O(N__69427),
            .I(N__69365));
    LocalMux I__17224 (
            .O(N__69424),
            .I(N__69360));
    Span4Mux_h I__17223 (
            .O(N__69421),
            .I(N__69360));
    LocalMux I__17222 (
            .O(N__69418),
            .I(N__69355));
    LocalMux I__17221 (
            .O(N__69413),
            .I(N__69355));
    Span4Mux_v I__17220 (
            .O(N__69410),
            .I(N__69352));
    Span4Mux_h I__17219 (
            .O(N__69405),
            .I(N__69349));
    Span4Mux_h I__17218 (
            .O(N__69400),
            .I(N__69344));
    Span4Mux_v I__17217 (
            .O(N__69397),
            .I(N__69344));
    Span4Mux_v I__17216 (
            .O(N__69394),
            .I(N__69341));
    LocalMux I__17215 (
            .O(N__69391),
            .I(N__69338));
    LocalMux I__17214 (
            .O(N__69388),
            .I(N__69335));
    LocalMux I__17213 (
            .O(N__69385),
            .I(N__69330));
    Sp12to4 I__17212 (
            .O(N__69376),
            .I(N__69330));
    InMux I__17211 (
            .O(N__69375),
            .I(N__69327));
    InMux I__17210 (
            .O(N__69374),
            .I(N__69324));
    Span4Mux_h I__17209 (
            .O(N__69371),
            .I(N__69319));
    Span4Mux_h I__17208 (
            .O(N__69368),
            .I(N__69319));
    Span4Mux_h I__17207 (
            .O(N__69365),
            .I(N__69314));
    Span4Mux_h I__17206 (
            .O(N__69360),
            .I(N__69314));
    Span12Mux_h I__17205 (
            .O(N__69355),
            .I(N__69309));
    Sp12to4 I__17204 (
            .O(N__69352),
            .I(N__69309));
    Span4Mux_h I__17203 (
            .O(N__69349),
            .I(N__69304));
    Span4Mux_v I__17202 (
            .O(N__69344),
            .I(N__69304));
    Sp12to4 I__17201 (
            .O(N__69341),
            .I(N__69295));
    Span12Mux_v I__17200 (
            .O(N__69338),
            .I(N__69295));
    Span12Mux_s8_h I__17199 (
            .O(N__69335),
            .I(N__69295));
    Span12Mux_v I__17198 (
            .O(N__69330),
            .I(N__69295));
    LocalMux I__17197 (
            .O(N__69327),
            .I(rx_data_0));
    LocalMux I__17196 (
            .O(N__69324),
            .I(rx_data_0));
    Odrv4 I__17195 (
            .O(N__69319),
            .I(rx_data_0));
    Odrv4 I__17194 (
            .O(N__69314),
            .I(rx_data_0));
    Odrv12 I__17193 (
            .O(N__69309),
            .I(rx_data_0));
    Odrv4 I__17192 (
            .O(N__69304),
            .I(rx_data_0));
    Odrv12 I__17191 (
            .O(N__69295),
            .I(rx_data_0));
    InMux I__17190 (
            .O(N__69280),
            .I(N__69276));
    CascadeMux I__17189 (
            .O(N__69279),
            .I(N__69273));
    LocalMux I__17188 (
            .O(N__69276),
            .I(N__69270));
    InMux I__17187 (
            .O(N__69273),
            .I(N__69266));
    Span4Mux_h I__17186 (
            .O(N__69270),
            .I(N__69263));
    InMux I__17185 (
            .O(N__69269),
            .I(N__69260));
    LocalMux I__17184 (
            .O(N__69266),
            .I(\c0.data_in_frame_26_0 ));
    Odrv4 I__17183 (
            .O(N__69263),
            .I(\c0.data_in_frame_26_0 ));
    LocalMux I__17182 (
            .O(N__69260),
            .I(\c0.data_in_frame_26_0 ));
    CascadeMux I__17181 (
            .O(N__69253),
            .I(N__69250));
    InMux I__17180 (
            .O(N__69250),
            .I(N__69246));
    InMux I__17179 (
            .O(N__69249),
            .I(N__69241));
    LocalMux I__17178 (
            .O(N__69246),
            .I(N__69238));
    CascadeMux I__17177 (
            .O(N__69245),
            .I(N__69235));
    CascadeMux I__17176 (
            .O(N__69244),
            .I(N__69228));
    LocalMux I__17175 (
            .O(N__69241),
            .I(N__69223));
    Span4Mux_h I__17174 (
            .O(N__69238),
            .I(N__69220));
    InMux I__17173 (
            .O(N__69235),
            .I(N__69217));
    CascadeMux I__17172 (
            .O(N__69234),
            .I(N__69214));
    CascadeMux I__17171 (
            .O(N__69233),
            .I(N__69207));
    CascadeMux I__17170 (
            .O(N__69232),
            .I(N__69200));
    InMux I__17169 (
            .O(N__69231),
            .I(N__69194));
    InMux I__17168 (
            .O(N__69228),
            .I(N__69184));
    InMux I__17167 (
            .O(N__69227),
            .I(N__69184));
    InMux I__17166 (
            .O(N__69226),
            .I(N__69184));
    Span4Mux_h I__17165 (
            .O(N__69223),
            .I(N__69177));
    Span4Mux_h I__17164 (
            .O(N__69220),
            .I(N__69177));
    LocalMux I__17163 (
            .O(N__69217),
            .I(N__69177));
    InMux I__17162 (
            .O(N__69214),
            .I(N__69174));
    InMux I__17161 (
            .O(N__69213),
            .I(N__69169));
    InMux I__17160 (
            .O(N__69212),
            .I(N__69169));
    InMux I__17159 (
            .O(N__69211),
            .I(N__69165));
    InMux I__17158 (
            .O(N__69210),
            .I(N__69162));
    InMux I__17157 (
            .O(N__69207),
            .I(N__69155));
    InMux I__17156 (
            .O(N__69206),
            .I(N__69155));
    InMux I__17155 (
            .O(N__69205),
            .I(N__69155));
    InMux I__17154 (
            .O(N__69204),
            .I(N__69152));
    InMux I__17153 (
            .O(N__69203),
            .I(N__69148));
    InMux I__17152 (
            .O(N__69200),
            .I(N__69143));
    InMux I__17151 (
            .O(N__69199),
            .I(N__69143));
    InMux I__17150 (
            .O(N__69198),
            .I(N__69138));
    InMux I__17149 (
            .O(N__69197),
            .I(N__69138));
    LocalMux I__17148 (
            .O(N__69194),
            .I(N__69135));
    CascadeMux I__17147 (
            .O(N__69193),
            .I(N__69132));
    CascadeMux I__17146 (
            .O(N__69192),
            .I(N__69129));
    CascadeMux I__17145 (
            .O(N__69191),
            .I(N__69126));
    LocalMux I__17144 (
            .O(N__69184),
            .I(N__69119));
    Span4Mux_v I__17143 (
            .O(N__69177),
            .I(N__69119));
    LocalMux I__17142 (
            .O(N__69174),
            .I(N__69116));
    LocalMux I__17141 (
            .O(N__69169),
            .I(N__69113));
    InMux I__17140 (
            .O(N__69168),
            .I(N__69110));
    LocalMux I__17139 (
            .O(N__69165),
            .I(N__69107));
    LocalMux I__17138 (
            .O(N__69162),
            .I(N__69100));
    LocalMux I__17137 (
            .O(N__69155),
            .I(N__69100));
    LocalMux I__17136 (
            .O(N__69152),
            .I(N__69100));
    InMux I__17135 (
            .O(N__69151),
            .I(N__69097));
    LocalMux I__17134 (
            .O(N__69148),
            .I(N__69094));
    LocalMux I__17133 (
            .O(N__69143),
            .I(N__69089));
    LocalMux I__17132 (
            .O(N__69138),
            .I(N__69089));
    Span4Mux_v I__17131 (
            .O(N__69135),
            .I(N__69086));
    InMux I__17130 (
            .O(N__69132),
            .I(N__69081));
    InMux I__17129 (
            .O(N__69129),
            .I(N__69081));
    InMux I__17128 (
            .O(N__69126),
            .I(N__69078));
    InMux I__17127 (
            .O(N__69125),
            .I(N__69075));
    InMux I__17126 (
            .O(N__69124),
            .I(N__69072));
    Sp12to4 I__17125 (
            .O(N__69119),
            .I(N__69069));
    Span4Mux_h I__17124 (
            .O(N__69116),
            .I(N__69066));
    Span4Mux_h I__17123 (
            .O(N__69113),
            .I(N__69059));
    LocalMux I__17122 (
            .O(N__69110),
            .I(N__69056));
    Span4Mux_h I__17121 (
            .O(N__69107),
            .I(N__69053));
    Span4Mux_v I__17120 (
            .O(N__69100),
            .I(N__69050));
    LocalMux I__17119 (
            .O(N__69097),
            .I(N__69043));
    Sp12to4 I__17118 (
            .O(N__69094),
            .I(N__69043));
    Span12Mux_v I__17117 (
            .O(N__69089),
            .I(N__69043));
    Span4Mux_h I__17116 (
            .O(N__69086),
            .I(N__69034));
    LocalMux I__17115 (
            .O(N__69081),
            .I(N__69034));
    LocalMux I__17114 (
            .O(N__69078),
            .I(N__69034));
    LocalMux I__17113 (
            .O(N__69075),
            .I(N__69034));
    LocalMux I__17112 (
            .O(N__69072),
            .I(N__69027));
    Span12Mux_h I__17111 (
            .O(N__69069),
            .I(N__69027));
    Sp12to4 I__17110 (
            .O(N__69066),
            .I(N__69027));
    InMux I__17109 (
            .O(N__69065),
            .I(N__69018));
    InMux I__17108 (
            .O(N__69064),
            .I(N__69018));
    InMux I__17107 (
            .O(N__69063),
            .I(N__69018));
    InMux I__17106 (
            .O(N__69062),
            .I(N__69018));
    Span4Mux_v I__17105 (
            .O(N__69059),
            .I(N__69015));
    Span4Mux_v I__17104 (
            .O(N__69056),
            .I(N__69008));
    Span4Mux_v I__17103 (
            .O(N__69053),
            .I(N__69008));
    Span4Mux_v I__17102 (
            .O(N__69050),
            .I(N__69008));
    Span12Mux_v I__17101 (
            .O(N__69043),
            .I(N__69005));
    Sp12to4 I__17100 (
            .O(N__69034),
            .I(N__69000));
    Span12Mux_v I__17099 (
            .O(N__69027),
            .I(N__69000));
    LocalMux I__17098 (
            .O(N__69018),
            .I(\c0.n9_adj_4341 ));
    Odrv4 I__17097 (
            .O(N__69015),
            .I(\c0.n9_adj_4341 ));
    Odrv4 I__17096 (
            .O(N__69008),
            .I(\c0.n9_adj_4341 ));
    Odrv12 I__17095 (
            .O(N__69005),
            .I(\c0.n9_adj_4341 ));
    Odrv12 I__17094 (
            .O(N__69000),
            .I(\c0.n9_adj_4341 ));
    InMux I__17093 (
            .O(N__68989),
            .I(N__68984));
    InMux I__17092 (
            .O(N__68988),
            .I(N__68981));
    InMux I__17091 (
            .O(N__68987),
            .I(N__68976));
    LocalMux I__17090 (
            .O(N__68984),
            .I(N__68965));
    LocalMux I__17089 (
            .O(N__68981),
            .I(N__68965));
    InMux I__17088 (
            .O(N__68980),
            .I(N__68962));
    InMux I__17087 (
            .O(N__68979),
            .I(N__68959));
    LocalMux I__17086 (
            .O(N__68976),
            .I(N__68951));
    InMux I__17085 (
            .O(N__68975),
            .I(N__68948));
    InMux I__17084 (
            .O(N__68974),
            .I(N__68945));
    CascadeMux I__17083 (
            .O(N__68973),
            .I(N__68941));
    InMux I__17082 (
            .O(N__68972),
            .I(N__68935));
    InMux I__17081 (
            .O(N__68971),
            .I(N__68932));
    InMux I__17080 (
            .O(N__68970),
            .I(N__68929));
    Span4Mux_v I__17079 (
            .O(N__68965),
            .I(N__68926));
    LocalMux I__17078 (
            .O(N__68962),
            .I(N__68921));
    LocalMux I__17077 (
            .O(N__68959),
            .I(N__68921));
    InMux I__17076 (
            .O(N__68958),
            .I(N__68916));
    InMux I__17075 (
            .O(N__68957),
            .I(N__68916));
    InMux I__17074 (
            .O(N__68956),
            .I(N__68913));
    InMux I__17073 (
            .O(N__68955),
            .I(N__68910));
    InMux I__17072 (
            .O(N__68954),
            .I(N__68905));
    Span4Mux_v I__17071 (
            .O(N__68951),
            .I(N__68900));
    LocalMux I__17070 (
            .O(N__68948),
            .I(N__68900));
    LocalMux I__17069 (
            .O(N__68945),
            .I(N__68897));
    InMux I__17068 (
            .O(N__68944),
            .I(N__68894));
    InMux I__17067 (
            .O(N__68941),
            .I(N__68889));
    InMux I__17066 (
            .O(N__68940),
            .I(N__68889));
    InMux I__17065 (
            .O(N__68939),
            .I(N__68884));
    InMux I__17064 (
            .O(N__68938),
            .I(N__68884));
    LocalMux I__17063 (
            .O(N__68935),
            .I(N__68877));
    LocalMux I__17062 (
            .O(N__68932),
            .I(N__68873));
    LocalMux I__17061 (
            .O(N__68929),
            .I(N__68868));
    Span4Mux_h I__17060 (
            .O(N__68926),
            .I(N__68868));
    Span4Mux_v I__17059 (
            .O(N__68921),
            .I(N__68862));
    LocalMux I__17058 (
            .O(N__68916),
            .I(N__68855));
    LocalMux I__17057 (
            .O(N__68913),
            .I(N__68855));
    LocalMux I__17056 (
            .O(N__68910),
            .I(N__68855));
    InMux I__17055 (
            .O(N__68909),
            .I(N__68852));
    InMux I__17054 (
            .O(N__68908),
            .I(N__68849));
    LocalMux I__17053 (
            .O(N__68905),
            .I(N__68846));
    Span4Mux_h I__17052 (
            .O(N__68900),
            .I(N__68837));
    Span4Mux_h I__17051 (
            .O(N__68897),
            .I(N__68837));
    LocalMux I__17050 (
            .O(N__68894),
            .I(N__68837));
    LocalMux I__17049 (
            .O(N__68889),
            .I(N__68837));
    LocalMux I__17048 (
            .O(N__68884),
            .I(N__68834));
    InMux I__17047 (
            .O(N__68883),
            .I(N__68831));
    InMux I__17046 (
            .O(N__68882),
            .I(N__68826));
    InMux I__17045 (
            .O(N__68881),
            .I(N__68826));
    InMux I__17044 (
            .O(N__68880),
            .I(N__68823));
    Span4Mux_h I__17043 (
            .O(N__68877),
            .I(N__68820));
    InMux I__17042 (
            .O(N__68876),
            .I(N__68817));
    Span4Mux_v I__17041 (
            .O(N__68873),
            .I(N__68812));
    Span4Mux_v I__17040 (
            .O(N__68868),
            .I(N__68812));
    InMux I__17039 (
            .O(N__68867),
            .I(N__68809));
    InMux I__17038 (
            .O(N__68866),
            .I(N__68806));
    InMux I__17037 (
            .O(N__68865),
            .I(N__68803));
    Span4Mux_h I__17036 (
            .O(N__68862),
            .I(N__68800));
    Span4Mux_v I__17035 (
            .O(N__68855),
            .I(N__68797));
    LocalMux I__17034 (
            .O(N__68852),
            .I(N__68792));
    LocalMux I__17033 (
            .O(N__68849),
            .I(N__68792));
    Span4Mux_h I__17032 (
            .O(N__68846),
            .I(N__68789));
    Span4Mux_v I__17031 (
            .O(N__68837),
            .I(N__68786));
    Span4Mux_v I__17030 (
            .O(N__68834),
            .I(N__68781));
    LocalMux I__17029 (
            .O(N__68831),
            .I(N__68776));
    LocalMux I__17028 (
            .O(N__68826),
            .I(N__68776));
    LocalMux I__17027 (
            .O(N__68823),
            .I(N__68771));
    Span4Mux_v I__17026 (
            .O(N__68820),
            .I(N__68771));
    LocalMux I__17025 (
            .O(N__68817),
            .I(N__68766));
    Span4Mux_v I__17024 (
            .O(N__68812),
            .I(N__68766));
    LocalMux I__17023 (
            .O(N__68809),
            .I(N__68763));
    LocalMux I__17022 (
            .O(N__68806),
            .I(N__68756));
    LocalMux I__17021 (
            .O(N__68803),
            .I(N__68756));
    Sp12to4 I__17020 (
            .O(N__68800),
            .I(N__68756));
    Sp12to4 I__17019 (
            .O(N__68797),
            .I(N__68753));
    Span4Mux_h I__17018 (
            .O(N__68792),
            .I(N__68746));
    Span4Mux_v I__17017 (
            .O(N__68789),
            .I(N__68746));
    Span4Mux_h I__17016 (
            .O(N__68786),
            .I(N__68746));
    InMux I__17015 (
            .O(N__68785),
            .I(N__68743));
    InMux I__17014 (
            .O(N__68784),
            .I(N__68740));
    Span4Mux_h I__17013 (
            .O(N__68781),
            .I(N__68731));
    Span4Mux_v I__17012 (
            .O(N__68776),
            .I(N__68731));
    Span4Mux_h I__17011 (
            .O(N__68771),
            .I(N__68731));
    Span4Mux_v I__17010 (
            .O(N__68766),
            .I(N__68731));
    Span12Mux_s11_v I__17009 (
            .O(N__68763),
            .I(N__68722));
    Span12Mux_s10_h I__17008 (
            .O(N__68756),
            .I(N__68722));
    Span12Mux_h I__17007 (
            .O(N__68753),
            .I(N__68722));
    Sp12to4 I__17006 (
            .O(N__68746),
            .I(N__68722));
    LocalMux I__17005 (
            .O(N__68743),
            .I(rx_data_7));
    LocalMux I__17004 (
            .O(N__68740),
            .I(rx_data_7));
    Odrv4 I__17003 (
            .O(N__68731),
            .I(rx_data_7));
    Odrv12 I__17002 (
            .O(N__68722),
            .I(rx_data_7));
    CascadeMux I__17001 (
            .O(N__68713),
            .I(N__68709));
    InMux I__17000 (
            .O(N__68712),
            .I(N__68706));
    InMux I__16999 (
            .O(N__68709),
            .I(N__68702));
    LocalMux I__16998 (
            .O(N__68706),
            .I(N__68699));
    CascadeMux I__16997 (
            .O(N__68705),
            .I(N__68696));
    LocalMux I__16996 (
            .O(N__68702),
            .I(N__68690));
    Span4Mux_h I__16995 (
            .O(N__68699),
            .I(N__68690));
    InMux I__16994 (
            .O(N__68696),
            .I(N__68685));
    InMux I__16993 (
            .O(N__68695),
            .I(N__68685));
    Odrv4 I__16992 (
            .O(N__68690),
            .I(\c0.data_in_frame_26_7 ));
    LocalMux I__16991 (
            .O(N__68685),
            .I(\c0.data_in_frame_26_7 ));
    CascadeMux I__16990 (
            .O(N__68680),
            .I(N__68675));
    CascadeMux I__16989 (
            .O(N__68679),
            .I(N__68666));
    InMux I__16988 (
            .O(N__68678),
            .I(N__68663));
    InMux I__16987 (
            .O(N__68675),
            .I(N__68660));
    InMux I__16986 (
            .O(N__68674),
            .I(N__68655));
    InMux I__16985 (
            .O(N__68673),
            .I(N__68650));
    InMux I__16984 (
            .O(N__68672),
            .I(N__68650));
    CascadeMux I__16983 (
            .O(N__68671),
            .I(N__68647));
    InMux I__16982 (
            .O(N__68670),
            .I(N__68644));
    InMux I__16981 (
            .O(N__68669),
            .I(N__68639));
    InMux I__16980 (
            .O(N__68666),
            .I(N__68639));
    LocalMux I__16979 (
            .O(N__68663),
            .I(N__68633));
    LocalMux I__16978 (
            .O(N__68660),
            .I(N__68633));
    CascadeMux I__16977 (
            .O(N__68659),
            .I(N__68629));
    CascadeMux I__16976 (
            .O(N__68658),
            .I(N__68625));
    LocalMux I__16975 (
            .O(N__68655),
            .I(N__68620));
    LocalMux I__16974 (
            .O(N__68650),
            .I(N__68620));
    InMux I__16973 (
            .O(N__68647),
            .I(N__68617));
    LocalMux I__16972 (
            .O(N__68644),
            .I(N__68614));
    LocalMux I__16971 (
            .O(N__68639),
            .I(N__68611));
    InMux I__16970 (
            .O(N__68638),
            .I(N__68608));
    Span4Mux_v I__16969 (
            .O(N__68633),
            .I(N__68605));
    InMux I__16968 (
            .O(N__68632),
            .I(N__68602));
    InMux I__16967 (
            .O(N__68629),
            .I(N__68595));
    InMux I__16966 (
            .O(N__68628),
            .I(N__68595));
    InMux I__16965 (
            .O(N__68625),
            .I(N__68592));
    Span4Mux_h I__16964 (
            .O(N__68620),
            .I(N__68584));
    LocalMux I__16963 (
            .O(N__68617),
            .I(N__68584));
    Span4Mux_h I__16962 (
            .O(N__68614),
            .I(N__68579));
    Span4Mux_v I__16961 (
            .O(N__68611),
            .I(N__68579));
    LocalMux I__16960 (
            .O(N__68608),
            .I(N__68576));
    Span4Mux_h I__16959 (
            .O(N__68605),
            .I(N__68571));
    LocalMux I__16958 (
            .O(N__68602),
            .I(N__68571));
    InMux I__16957 (
            .O(N__68601),
            .I(N__68565));
    InMux I__16956 (
            .O(N__68600),
            .I(N__68562));
    LocalMux I__16955 (
            .O(N__68595),
            .I(N__68557));
    LocalMux I__16954 (
            .O(N__68592),
            .I(N__68557));
    InMux I__16953 (
            .O(N__68591),
            .I(N__68554));
    CascadeMux I__16952 (
            .O(N__68590),
            .I(N__68549));
    InMux I__16951 (
            .O(N__68589),
            .I(N__68546));
    Span4Mux_h I__16950 (
            .O(N__68584),
            .I(N__68542));
    Span4Mux_h I__16949 (
            .O(N__68579),
            .I(N__68539));
    Span4Mux_h I__16948 (
            .O(N__68576),
            .I(N__68536));
    Span4Mux_v I__16947 (
            .O(N__68571),
            .I(N__68533));
    InMux I__16946 (
            .O(N__68570),
            .I(N__68530));
    InMux I__16945 (
            .O(N__68569),
            .I(N__68527));
    InMux I__16944 (
            .O(N__68568),
            .I(N__68524));
    LocalMux I__16943 (
            .O(N__68565),
            .I(N__68517));
    LocalMux I__16942 (
            .O(N__68562),
            .I(N__68517));
    Span4Mux_v I__16941 (
            .O(N__68557),
            .I(N__68517));
    LocalMux I__16940 (
            .O(N__68554),
            .I(N__68513));
    InMux I__16939 (
            .O(N__68553),
            .I(N__68506));
    InMux I__16938 (
            .O(N__68552),
            .I(N__68506));
    InMux I__16937 (
            .O(N__68549),
            .I(N__68506));
    LocalMux I__16936 (
            .O(N__68546),
            .I(N__68503));
    InMux I__16935 (
            .O(N__68545),
            .I(N__68500));
    Span4Mux_h I__16934 (
            .O(N__68542),
            .I(N__68493));
    Span4Mux_h I__16933 (
            .O(N__68539),
            .I(N__68493));
    Span4Mux_v I__16932 (
            .O(N__68536),
            .I(N__68493));
    Sp12to4 I__16931 (
            .O(N__68533),
            .I(N__68488));
    LocalMux I__16930 (
            .O(N__68530),
            .I(N__68488));
    LocalMux I__16929 (
            .O(N__68527),
            .I(N__68485));
    LocalMux I__16928 (
            .O(N__68524),
            .I(N__68480));
    Span4Mux_v I__16927 (
            .O(N__68517),
            .I(N__68480));
    InMux I__16926 (
            .O(N__68516),
            .I(N__68477));
    Sp12to4 I__16925 (
            .O(N__68513),
            .I(N__68468));
    LocalMux I__16924 (
            .O(N__68506),
            .I(N__68468));
    Span12Mux_v I__16923 (
            .O(N__68503),
            .I(N__68468));
    LocalMux I__16922 (
            .O(N__68500),
            .I(N__68468));
    Sp12to4 I__16921 (
            .O(N__68493),
            .I(N__68463));
    Span12Mux_h I__16920 (
            .O(N__68488),
            .I(N__68463));
    Span4Mux_v I__16919 (
            .O(N__68485),
            .I(N__68460));
    Span4Mux_h I__16918 (
            .O(N__68480),
            .I(N__68457));
    LocalMux I__16917 (
            .O(N__68477),
            .I(N__68450));
    Span12Mux_v I__16916 (
            .O(N__68468),
            .I(N__68450));
    Span12Mux_v I__16915 (
            .O(N__68463),
            .I(N__68450));
    Odrv4 I__16914 (
            .O(N__68460),
            .I(\c0.n17596 ));
    Odrv4 I__16913 (
            .O(N__68457),
            .I(\c0.n17596 ));
    Odrv12 I__16912 (
            .O(N__68450),
            .I(\c0.n17596 ));
    InMux I__16911 (
            .O(N__68443),
            .I(N__68438));
    CascadeMux I__16910 (
            .O(N__68442),
            .I(N__68430));
    CascadeMux I__16909 (
            .O(N__68441),
            .I(N__68427));
    LocalMux I__16908 (
            .O(N__68438),
            .I(N__68423));
    InMux I__16907 (
            .O(N__68437),
            .I(N__68420));
    CascadeMux I__16906 (
            .O(N__68436),
            .I(N__68413));
    InMux I__16905 (
            .O(N__68435),
            .I(N__68407));
    InMux I__16904 (
            .O(N__68434),
            .I(N__68404));
    InMux I__16903 (
            .O(N__68433),
            .I(N__68399));
    InMux I__16902 (
            .O(N__68430),
            .I(N__68399));
    InMux I__16901 (
            .O(N__68427),
            .I(N__68396));
    InMux I__16900 (
            .O(N__68426),
            .I(N__68390));
    Span4Mux_v I__16899 (
            .O(N__68423),
            .I(N__68385));
    LocalMux I__16898 (
            .O(N__68420),
            .I(N__68385));
    InMux I__16897 (
            .O(N__68419),
            .I(N__68378));
    InMux I__16896 (
            .O(N__68418),
            .I(N__68378));
    InMux I__16895 (
            .O(N__68417),
            .I(N__68378));
    InMux I__16894 (
            .O(N__68416),
            .I(N__68374));
    InMux I__16893 (
            .O(N__68413),
            .I(N__68370));
    InMux I__16892 (
            .O(N__68412),
            .I(N__68366));
    CascadeMux I__16891 (
            .O(N__68411),
            .I(N__68363));
    InMux I__16890 (
            .O(N__68410),
            .I(N__68360));
    LocalMux I__16889 (
            .O(N__68407),
            .I(N__68349));
    LocalMux I__16888 (
            .O(N__68404),
            .I(N__68346));
    LocalMux I__16887 (
            .O(N__68399),
            .I(N__68341));
    LocalMux I__16886 (
            .O(N__68396),
            .I(N__68341));
    InMux I__16885 (
            .O(N__68395),
            .I(N__68338));
    InMux I__16884 (
            .O(N__68394),
            .I(N__68333));
    InMux I__16883 (
            .O(N__68393),
            .I(N__68333));
    LocalMux I__16882 (
            .O(N__68390),
            .I(N__68330));
    Span4Mux_h I__16881 (
            .O(N__68385),
            .I(N__68325));
    LocalMux I__16880 (
            .O(N__68378),
            .I(N__68325));
    InMux I__16879 (
            .O(N__68377),
            .I(N__68322));
    LocalMux I__16878 (
            .O(N__68374),
            .I(N__68319));
    InMux I__16877 (
            .O(N__68373),
            .I(N__68316));
    LocalMux I__16876 (
            .O(N__68370),
            .I(N__68313));
    InMux I__16875 (
            .O(N__68369),
            .I(N__68310));
    LocalMux I__16874 (
            .O(N__68366),
            .I(N__68307));
    InMux I__16873 (
            .O(N__68363),
            .I(N__68304));
    LocalMux I__16872 (
            .O(N__68360),
            .I(N__68301));
    InMux I__16871 (
            .O(N__68359),
            .I(N__68296));
    InMux I__16870 (
            .O(N__68358),
            .I(N__68296));
    InMux I__16869 (
            .O(N__68357),
            .I(N__68293));
    InMux I__16868 (
            .O(N__68356),
            .I(N__68290));
    InMux I__16867 (
            .O(N__68355),
            .I(N__68285));
    InMux I__16866 (
            .O(N__68354),
            .I(N__68280));
    InMux I__16865 (
            .O(N__68353),
            .I(N__68280));
    InMux I__16864 (
            .O(N__68352),
            .I(N__68277));
    Span4Mux_v I__16863 (
            .O(N__68349),
            .I(N__68274));
    Span4Mux_h I__16862 (
            .O(N__68346),
            .I(N__68269));
    Span4Mux_v I__16861 (
            .O(N__68341),
            .I(N__68269));
    LocalMux I__16860 (
            .O(N__68338),
            .I(N__68262));
    LocalMux I__16859 (
            .O(N__68333),
            .I(N__68262));
    Span4Mux_v I__16858 (
            .O(N__68330),
            .I(N__68262));
    Span4Mux_v I__16857 (
            .O(N__68325),
            .I(N__68259));
    LocalMux I__16856 (
            .O(N__68322),
            .I(N__68256));
    Span4Mux_h I__16855 (
            .O(N__68319),
            .I(N__68251));
    LocalMux I__16854 (
            .O(N__68316),
            .I(N__68251));
    Span4Mux_v I__16853 (
            .O(N__68313),
            .I(N__68248));
    LocalMux I__16852 (
            .O(N__68310),
            .I(N__68243));
    Span4Mux_v I__16851 (
            .O(N__68307),
            .I(N__68243));
    LocalMux I__16850 (
            .O(N__68304),
            .I(N__68238));
    Span4Mux_v I__16849 (
            .O(N__68301),
            .I(N__68238));
    LocalMux I__16848 (
            .O(N__68296),
            .I(N__68235));
    LocalMux I__16847 (
            .O(N__68293),
            .I(N__68230));
    LocalMux I__16846 (
            .O(N__68290),
            .I(N__68230));
    InMux I__16845 (
            .O(N__68289),
            .I(N__68227));
    InMux I__16844 (
            .O(N__68288),
            .I(N__68224));
    LocalMux I__16843 (
            .O(N__68285),
            .I(N__68219));
    LocalMux I__16842 (
            .O(N__68280),
            .I(N__68219));
    LocalMux I__16841 (
            .O(N__68277),
            .I(N__68216));
    Span4Mux_v I__16840 (
            .O(N__68274),
            .I(N__68211));
    Span4Mux_v I__16839 (
            .O(N__68269),
            .I(N__68211));
    Span4Mux_v I__16838 (
            .O(N__68262),
            .I(N__68208));
    Span4Mux_h I__16837 (
            .O(N__68259),
            .I(N__68205));
    Span4Mux_v I__16836 (
            .O(N__68256),
            .I(N__68196));
    Span4Mux_v I__16835 (
            .O(N__68251),
            .I(N__68196));
    Span4Mux_h I__16834 (
            .O(N__68248),
            .I(N__68196));
    Span4Mux_v I__16833 (
            .O(N__68243),
            .I(N__68196));
    Span4Mux_v I__16832 (
            .O(N__68238),
            .I(N__68189));
    Span4Mux_v I__16831 (
            .O(N__68235),
            .I(N__68189));
    Span4Mux_h I__16830 (
            .O(N__68230),
            .I(N__68189));
    LocalMux I__16829 (
            .O(N__68227),
            .I(N__68178));
    LocalMux I__16828 (
            .O(N__68224),
            .I(N__68178));
    Span12Mux_v I__16827 (
            .O(N__68219),
            .I(N__68178));
    Span12Mux_v I__16826 (
            .O(N__68216),
            .I(N__68178));
    Sp12to4 I__16825 (
            .O(N__68211),
            .I(N__68178));
    Odrv4 I__16824 (
            .O(N__68208),
            .I(rx_data_2));
    Odrv4 I__16823 (
            .O(N__68205),
            .I(rx_data_2));
    Odrv4 I__16822 (
            .O(N__68196),
            .I(rx_data_2));
    Odrv4 I__16821 (
            .O(N__68189),
            .I(rx_data_2));
    Odrv12 I__16820 (
            .O(N__68178),
            .I(rx_data_2));
    InMux I__16819 (
            .O(N__68167),
            .I(N__68152));
    InMux I__16818 (
            .O(N__68166),
            .I(N__68149));
    InMux I__16817 (
            .O(N__68165),
            .I(N__68132));
    CascadeMux I__16816 (
            .O(N__68164),
            .I(N__68129));
    InMux I__16815 (
            .O(N__68163),
            .I(N__68122));
    InMux I__16814 (
            .O(N__68162),
            .I(N__68122));
    InMux I__16813 (
            .O(N__68161),
            .I(N__68122));
    InMux I__16812 (
            .O(N__68160),
            .I(N__68117));
    InMux I__16811 (
            .O(N__68159),
            .I(N__68117));
    InMux I__16810 (
            .O(N__68158),
            .I(N__68112));
    InMux I__16809 (
            .O(N__68157),
            .I(N__68112));
    InMux I__16808 (
            .O(N__68156),
            .I(N__68104));
    InMux I__16807 (
            .O(N__68155),
            .I(N__68104));
    LocalMux I__16806 (
            .O(N__68152),
            .I(N__68101));
    LocalMux I__16805 (
            .O(N__68149),
            .I(N__68098));
    InMux I__16804 (
            .O(N__68148),
            .I(N__68088));
    CascadeMux I__16803 (
            .O(N__68147),
            .I(N__68083));
    InMux I__16802 (
            .O(N__68146),
            .I(N__68078));
    InMux I__16801 (
            .O(N__68145),
            .I(N__68078));
    InMux I__16800 (
            .O(N__68144),
            .I(N__68071));
    InMux I__16799 (
            .O(N__68143),
            .I(N__68071));
    InMux I__16798 (
            .O(N__68142),
            .I(N__68071));
    InMux I__16797 (
            .O(N__68141),
            .I(N__68062));
    InMux I__16796 (
            .O(N__68140),
            .I(N__68057));
    InMux I__16795 (
            .O(N__68139),
            .I(N__68057));
    InMux I__16794 (
            .O(N__68138),
            .I(N__68048));
    InMux I__16793 (
            .O(N__68137),
            .I(N__68048));
    InMux I__16792 (
            .O(N__68136),
            .I(N__68048));
    InMux I__16791 (
            .O(N__68135),
            .I(N__68048));
    LocalMux I__16790 (
            .O(N__68132),
            .I(N__68045));
    InMux I__16789 (
            .O(N__68129),
            .I(N__68039));
    LocalMux I__16788 (
            .O(N__68122),
            .I(N__68036));
    LocalMux I__16787 (
            .O(N__68117),
            .I(N__68033));
    LocalMux I__16786 (
            .O(N__68112),
            .I(N__68030));
    InMux I__16785 (
            .O(N__68111),
            .I(N__68023));
    InMux I__16784 (
            .O(N__68110),
            .I(N__68023));
    InMux I__16783 (
            .O(N__68109),
            .I(N__68023));
    LocalMux I__16782 (
            .O(N__68104),
            .I(N__68020));
    Span4Mux_v I__16781 (
            .O(N__68101),
            .I(N__68012));
    Span4Mux_h I__16780 (
            .O(N__68098),
            .I(N__68012));
    InMux I__16779 (
            .O(N__68097),
            .I(N__68009));
    InMux I__16778 (
            .O(N__68096),
            .I(N__68003));
    InMux I__16777 (
            .O(N__68095),
            .I(N__68000));
    InMux I__16776 (
            .O(N__68094),
            .I(N__67995));
    InMux I__16775 (
            .O(N__68093),
            .I(N__67995));
    InMux I__16774 (
            .O(N__68092),
            .I(N__67990));
    InMux I__16773 (
            .O(N__68091),
            .I(N__67990));
    LocalMux I__16772 (
            .O(N__68088),
            .I(N__67987));
    InMux I__16771 (
            .O(N__68087),
            .I(N__67984));
    InMux I__16770 (
            .O(N__68086),
            .I(N__67979));
    InMux I__16769 (
            .O(N__68083),
            .I(N__67979));
    LocalMux I__16768 (
            .O(N__68078),
            .I(N__67974));
    LocalMux I__16767 (
            .O(N__68071),
            .I(N__67974));
    InMux I__16766 (
            .O(N__68070),
            .I(N__67971));
    InMux I__16765 (
            .O(N__68069),
            .I(N__67966));
    InMux I__16764 (
            .O(N__68068),
            .I(N__67966));
    InMux I__16763 (
            .O(N__68067),
            .I(N__67959));
    InMux I__16762 (
            .O(N__68066),
            .I(N__67959));
    InMux I__16761 (
            .O(N__68065),
            .I(N__67959));
    LocalMux I__16760 (
            .O(N__68062),
            .I(N__67954));
    LocalMux I__16759 (
            .O(N__68057),
            .I(N__67954));
    LocalMux I__16758 (
            .O(N__68048),
            .I(N__67949));
    Span4Mux_v I__16757 (
            .O(N__68045),
            .I(N__67949));
    CascadeMux I__16756 (
            .O(N__68044),
            .I(N__67946));
    InMux I__16755 (
            .O(N__68043),
            .I(N__67941));
    InMux I__16754 (
            .O(N__68042),
            .I(N__67941));
    LocalMux I__16753 (
            .O(N__68039),
            .I(N__67938));
    Span4Mux_v I__16752 (
            .O(N__68036),
            .I(N__67933));
    Span4Mux_v I__16751 (
            .O(N__68033),
            .I(N__67933));
    Span4Mux_h I__16750 (
            .O(N__68030),
            .I(N__67926));
    LocalMux I__16749 (
            .O(N__68023),
            .I(N__67926));
    Span4Mux_v I__16748 (
            .O(N__68020),
            .I(N__67926));
    InMux I__16747 (
            .O(N__68019),
            .I(N__67919));
    InMux I__16746 (
            .O(N__68018),
            .I(N__67919));
    InMux I__16745 (
            .O(N__68017),
            .I(N__67919));
    Span4Mux_h I__16744 (
            .O(N__68012),
            .I(N__67916));
    LocalMux I__16743 (
            .O(N__68009),
            .I(N__67913));
    InMux I__16742 (
            .O(N__68008),
            .I(N__67904));
    InMux I__16741 (
            .O(N__68007),
            .I(N__67904));
    InMux I__16740 (
            .O(N__68006),
            .I(N__67904));
    LocalMux I__16739 (
            .O(N__68003),
            .I(N__67901));
    LocalMux I__16738 (
            .O(N__68000),
            .I(N__67892));
    LocalMux I__16737 (
            .O(N__67995),
            .I(N__67892));
    LocalMux I__16736 (
            .O(N__67990),
            .I(N__67892));
    Span4Mux_h I__16735 (
            .O(N__67987),
            .I(N__67892));
    LocalMux I__16734 (
            .O(N__67984),
            .I(N__67885));
    LocalMux I__16733 (
            .O(N__67979),
            .I(N__67885));
    Span4Mux_v I__16732 (
            .O(N__67974),
            .I(N__67885));
    LocalMux I__16731 (
            .O(N__67971),
            .I(N__67874));
    LocalMux I__16730 (
            .O(N__67966),
            .I(N__67874));
    LocalMux I__16729 (
            .O(N__67959),
            .I(N__67874));
    Span4Mux_v I__16728 (
            .O(N__67954),
            .I(N__67874));
    Span4Mux_h I__16727 (
            .O(N__67949),
            .I(N__67874));
    InMux I__16726 (
            .O(N__67946),
            .I(N__67871));
    LocalMux I__16725 (
            .O(N__67941),
            .I(N__67866));
    Span4Mux_v I__16724 (
            .O(N__67938),
            .I(N__67866));
    Span4Mux_v I__16723 (
            .O(N__67933),
            .I(N__67861));
    Span4Mux_v I__16722 (
            .O(N__67926),
            .I(N__67861));
    LocalMux I__16721 (
            .O(N__67919),
            .I(N__67854));
    Span4Mux_v I__16720 (
            .O(N__67916),
            .I(N__67854));
    Span4Mux_h I__16719 (
            .O(N__67913),
            .I(N__67854));
    InMux I__16718 (
            .O(N__67912),
            .I(N__67849));
    InMux I__16717 (
            .O(N__67911),
            .I(N__67849));
    LocalMux I__16716 (
            .O(N__67904),
            .I(N__67838));
    Span4Mux_v I__16715 (
            .O(N__67901),
            .I(N__67838));
    Span4Mux_v I__16714 (
            .O(N__67892),
            .I(N__67838));
    Span4Mux_h I__16713 (
            .O(N__67885),
            .I(N__67838));
    Span4Mux_v I__16712 (
            .O(N__67874),
            .I(N__67838));
    LocalMux I__16711 (
            .O(N__67871),
            .I(N__67831));
    Span4Mux_h I__16710 (
            .O(N__67866),
            .I(N__67831));
    Span4Mux_h I__16709 (
            .O(N__67861),
            .I(N__67831));
    Span4Mux_v I__16708 (
            .O(N__67854),
            .I(N__67828));
    LocalMux I__16707 (
            .O(N__67849),
            .I(\c0.n21758 ));
    Odrv4 I__16706 (
            .O(N__67838),
            .I(\c0.n21758 ));
    Odrv4 I__16705 (
            .O(N__67831),
            .I(\c0.n21758 ));
    Odrv4 I__16704 (
            .O(N__67828),
            .I(\c0.n21758 ));
    CascadeMux I__16703 (
            .O(N__67819),
            .I(N__67815));
    InMux I__16702 (
            .O(N__67818),
            .I(N__67812));
    InMux I__16701 (
            .O(N__67815),
            .I(N__67808));
    LocalMux I__16700 (
            .O(N__67812),
            .I(N__67805));
    InMux I__16699 (
            .O(N__67811),
            .I(N__67802));
    LocalMux I__16698 (
            .O(N__67808),
            .I(\c0.data_in_frame_23_2 ));
    Odrv12 I__16697 (
            .O(N__67805),
            .I(\c0.data_in_frame_23_2 ));
    LocalMux I__16696 (
            .O(N__67802),
            .I(\c0.data_in_frame_23_2 ));
    InMux I__16695 (
            .O(N__67795),
            .I(N__67784));
    InMux I__16694 (
            .O(N__67794),
            .I(N__67784));
    InMux I__16693 (
            .O(N__67793),
            .I(N__67784));
    InMux I__16692 (
            .O(N__67792),
            .I(N__67779));
    InMux I__16691 (
            .O(N__67791),
            .I(N__67779));
    LocalMux I__16690 (
            .O(N__67784),
            .I(N__67770));
    LocalMux I__16689 (
            .O(N__67779),
            .I(N__67770));
    InMux I__16688 (
            .O(N__67778),
            .I(N__67765));
    InMux I__16687 (
            .O(N__67777),
            .I(N__67765));
    InMux I__16686 (
            .O(N__67776),
            .I(N__67753));
    InMux I__16685 (
            .O(N__67775),
            .I(N__67745));
    Span4Mux_v I__16684 (
            .O(N__67770),
            .I(N__67739));
    LocalMux I__16683 (
            .O(N__67765),
            .I(N__67739));
    InMux I__16682 (
            .O(N__67764),
            .I(N__67734));
    InMux I__16681 (
            .O(N__67763),
            .I(N__67734));
    InMux I__16680 (
            .O(N__67762),
            .I(N__67724));
    InMux I__16679 (
            .O(N__67761),
            .I(N__67724));
    InMux I__16678 (
            .O(N__67760),
            .I(N__67724));
    InMux I__16677 (
            .O(N__67759),
            .I(N__67721));
    InMux I__16676 (
            .O(N__67758),
            .I(N__67718));
    InMux I__16675 (
            .O(N__67757),
            .I(N__67715));
    InMux I__16674 (
            .O(N__67756),
            .I(N__67712));
    LocalMux I__16673 (
            .O(N__67753),
            .I(N__67709));
    InMux I__16672 (
            .O(N__67752),
            .I(N__67702));
    InMux I__16671 (
            .O(N__67751),
            .I(N__67699));
    InMux I__16670 (
            .O(N__67750),
            .I(N__67692));
    InMux I__16669 (
            .O(N__67749),
            .I(N__67692));
    InMux I__16668 (
            .O(N__67748),
            .I(N__67692));
    LocalMux I__16667 (
            .O(N__67745),
            .I(N__67689));
    InMux I__16666 (
            .O(N__67744),
            .I(N__67686));
    Span4Mux_v I__16665 (
            .O(N__67739),
            .I(N__67682));
    LocalMux I__16664 (
            .O(N__67734),
            .I(N__67679));
    InMux I__16663 (
            .O(N__67733),
            .I(N__67665));
    InMux I__16662 (
            .O(N__67732),
            .I(N__67665));
    InMux I__16661 (
            .O(N__67731),
            .I(N__67665));
    LocalMux I__16660 (
            .O(N__67724),
            .I(N__67662));
    LocalMux I__16659 (
            .O(N__67721),
            .I(N__67659));
    LocalMux I__16658 (
            .O(N__67718),
            .I(N__67656));
    LocalMux I__16657 (
            .O(N__67715),
            .I(N__67649));
    LocalMux I__16656 (
            .O(N__67712),
            .I(N__67649));
    Span4Mux_v I__16655 (
            .O(N__67709),
            .I(N__67649));
    InMux I__16654 (
            .O(N__67708),
            .I(N__67646));
    InMux I__16653 (
            .O(N__67707),
            .I(N__67643));
    InMux I__16652 (
            .O(N__67706),
            .I(N__67638));
    InMux I__16651 (
            .O(N__67705),
            .I(N__67638));
    LocalMux I__16650 (
            .O(N__67702),
            .I(N__67633));
    LocalMux I__16649 (
            .O(N__67699),
            .I(N__67633));
    LocalMux I__16648 (
            .O(N__67692),
            .I(N__67630));
    Span4Mux_v I__16647 (
            .O(N__67689),
            .I(N__67625));
    LocalMux I__16646 (
            .O(N__67686),
            .I(N__67625));
    InMux I__16645 (
            .O(N__67685),
            .I(N__67617));
    Span4Mux_h I__16644 (
            .O(N__67682),
            .I(N__67612));
    Span4Mux_v I__16643 (
            .O(N__67679),
            .I(N__67612));
    InMux I__16642 (
            .O(N__67678),
            .I(N__67606));
    InMux I__16641 (
            .O(N__67677),
            .I(N__67603));
    InMux I__16640 (
            .O(N__67676),
            .I(N__67600));
    InMux I__16639 (
            .O(N__67675),
            .I(N__67597));
    InMux I__16638 (
            .O(N__67674),
            .I(N__67592));
    InMux I__16637 (
            .O(N__67673),
            .I(N__67592));
    InMux I__16636 (
            .O(N__67672),
            .I(N__67589));
    LocalMux I__16635 (
            .O(N__67665),
            .I(N__67586));
    Span4Mux_v I__16634 (
            .O(N__67662),
            .I(N__67583));
    Span4Mux_v I__16633 (
            .O(N__67659),
            .I(N__67576));
    Span4Mux_v I__16632 (
            .O(N__67656),
            .I(N__67576));
    Span4Mux_v I__16631 (
            .O(N__67649),
            .I(N__67576));
    LocalMux I__16630 (
            .O(N__67646),
            .I(N__67573));
    LocalMux I__16629 (
            .O(N__67643),
            .I(N__67564));
    LocalMux I__16628 (
            .O(N__67638),
            .I(N__67564));
    Span4Mux_v I__16627 (
            .O(N__67633),
            .I(N__67564));
    Span4Mux_h I__16626 (
            .O(N__67630),
            .I(N__67564));
    Span4Mux_v I__16625 (
            .O(N__67625),
            .I(N__67561));
    InMux I__16624 (
            .O(N__67624),
            .I(N__67556));
    InMux I__16623 (
            .O(N__67623),
            .I(N__67556));
    InMux I__16622 (
            .O(N__67622),
            .I(N__67553));
    InMux I__16621 (
            .O(N__67621),
            .I(N__67548));
    InMux I__16620 (
            .O(N__67620),
            .I(N__67548));
    LocalMux I__16619 (
            .O(N__67617),
            .I(N__67545));
    Span4Mux_h I__16618 (
            .O(N__67612),
            .I(N__67542));
    InMux I__16617 (
            .O(N__67611),
            .I(N__67539));
    InMux I__16616 (
            .O(N__67610),
            .I(N__67536));
    InMux I__16615 (
            .O(N__67609),
            .I(N__67533));
    LocalMux I__16614 (
            .O(N__67606),
            .I(N__67522));
    LocalMux I__16613 (
            .O(N__67603),
            .I(N__67522));
    LocalMux I__16612 (
            .O(N__67600),
            .I(N__67522));
    LocalMux I__16611 (
            .O(N__67597),
            .I(N__67522));
    LocalMux I__16610 (
            .O(N__67592),
            .I(N__67522));
    LocalMux I__16609 (
            .O(N__67589),
            .I(N__67513));
    Span4Mux_v I__16608 (
            .O(N__67586),
            .I(N__67513));
    Span4Mux_v I__16607 (
            .O(N__67583),
            .I(N__67513));
    Span4Mux_h I__16606 (
            .O(N__67576),
            .I(N__67513));
    Span4Mux_v I__16605 (
            .O(N__67573),
            .I(N__67506));
    Span4Mux_v I__16604 (
            .O(N__67564),
            .I(N__67506));
    Span4Mux_h I__16603 (
            .O(N__67561),
            .I(N__67506));
    LocalMux I__16602 (
            .O(N__67556),
            .I(N__67495));
    LocalMux I__16601 (
            .O(N__67553),
            .I(N__67495));
    LocalMux I__16600 (
            .O(N__67548),
            .I(N__67495));
    Span4Mux_v I__16599 (
            .O(N__67545),
            .I(N__67495));
    Span4Mux_h I__16598 (
            .O(N__67542),
            .I(N__67495));
    LocalMux I__16597 (
            .O(N__67539),
            .I(\c0.n21775 ));
    LocalMux I__16596 (
            .O(N__67536),
            .I(\c0.n21775 ));
    LocalMux I__16595 (
            .O(N__67533),
            .I(\c0.n21775 ));
    Odrv12 I__16594 (
            .O(N__67522),
            .I(\c0.n21775 ));
    Odrv4 I__16593 (
            .O(N__67513),
            .I(\c0.n21775 ));
    Odrv4 I__16592 (
            .O(N__67506),
            .I(\c0.n21775 ));
    Odrv4 I__16591 (
            .O(N__67495),
            .I(\c0.n21775 ));
    CascadeMux I__16590 (
            .O(N__67480),
            .I(N__67472));
    CascadeMux I__16589 (
            .O(N__67479),
            .I(N__67466));
    CascadeMux I__16588 (
            .O(N__67478),
            .I(N__67463));
    InMux I__16587 (
            .O(N__67477),
            .I(N__67454));
    InMux I__16586 (
            .O(N__67476),
            .I(N__67446));
    InMux I__16585 (
            .O(N__67475),
            .I(N__67446));
    InMux I__16584 (
            .O(N__67472),
            .I(N__67440));
    InMux I__16583 (
            .O(N__67471),
            .I(N__67440));
    InMux I__16582 (
            .O(N__67470),
            .I(N__67437));
    InMux I__16581 (
            .O(N__67469),
            .I(N__67434));
    InMux I__16580 (
            .O(N__67466),
            .I(N__67425));
    InMux I__16579 (
            .O(N__67463),
            .I(N__67425));
    InMux I__16578 (
            .O(N__67462),
            .I(N__67425));
    InMux I__16577 (
            .O(N__67461),
            .I(N__67425));
    InMux I__16576 (
            .O(N__67460),
            .I(N__67418));
    InMux I__16575 (
            .O(N__67459),
            .I(N__67418));
    InMux I__16574 (
            .O(N__67458),
            .I(N__67418));
    InMux I__16573 (
            .O(N__67457),
            .I(N__67415));
    LocalMux I__16572 (
            .O(N__67454),
            .I(N__67412));
    InMux I__16571 (
            .O(N__67453),
            .I(N__67409));
    InMux I__16570 (
            .O(N__67452),
            .I(N__67404));
    InMux I__16569 (
            .O(N__67451),
            .I(N__67399));
    LocalMux I__16568 (
            .O(N__67446),
            .I(N__67396));
    InMux I__16567 (
            .O(N__67445),
            .I(N__67393));
    LocalMux I__16566 (
            .O(N__67440),
            .I(N__67386));
    LocalMux I__16565 (
            .O(N__67437),
            .I(N__67386));
    LocalMux I__16564 (
            .O(N__67434),
            .I(N__67383));
    LocalMux I__16563 (
            .O(N__67425),
            .I(N__67380));
    LocalMux I__16562 (
            .O(N__67418),
            .I(N__67376));
    LocalMux I__16561 (
            .O(N__67415),
            .I(N__67373));
    Span4Mux_h I__16560 (
            .O(N__67412),
            .I(N__67368));
    LocalMux I__16559 (
            .O(N__67409),
            .I(N__67368));
    InMux I__16558 (
            .O(N__67408),
            .I(N__67365));
    InMux I__16557 (
            .O(N__67407),
            .I(N__67358));
    LocalMux I__16556 (
            .O(N__67404),
            .I(N__67355));
    InMux I__16555 (
            .O(N__67403),
            .I(N__67352));
    CascadeMux I__16554 (
            .O(N__67402),
            .I(N__67349));
    LocalMux I__16553 (
            .O(N__67399),
            .I(N__67345));
    Span4Mux_h I__16552 (
            .O(N__67396),
            .I(N__67340));
    LocalMux I__16551 (
            .O(N__67393),
            .I(N__67340));
    InMux I__16550 (
            .O(N__67392),
            .I(N__67334));
    InMux I__16549 (
            .O(N__67391),
            .I(N__67334));
    Span4Mux_v I__16548 (
            .O(N__67386),
            .I(N__67331));
    Span4Mux_v I__16547 (
            .O(N__67383),
            .I(N__67326));
    Span4Mux_v I__16546 (
            .O(N__67380),
            .I(N__67326));
    InMux I__16545 (
            .O(N__67379),
            .I(N__67323));
    Span4Mux_v I__16544 (
            .O(N__67376),
            .I(N__67320));
    Span4Mux_v I__16543 (
            .O(N__67373),
            .I(N__67317));
    Span4Mux_v I__16542 (
            .O(N__67368),
            .I(N__67312));
    LocalMux I__16541 (
            .O(N__67365),
            .I(N__67312));
    InMux I__16540 (
            .O(N__67364),
            .I(N__67307));
    InMux I__16539 (
            .O(N__67363),
            .I(N__67307));
    InMux I__16538 (
            .O(N__67362),
            .I(N__67304));
    InMux I__16537 (
            .O(N__67361),
            .I(N__67301));
    LocalMux I__16536 (
            .O(N__67358),
            .I(N__67296));
    Span4Mux_v I__16535 (
            .O(N__67355),
            .I(N__67296));
    LocalMux I__16534 (
            .O(N__67352),
            .I(N__67293));
    InMux I__16533 (
            .O(N__67349),
            .I(N__67290));
    InMux I__16532 (
            .O(N__67348),
            .I(N__67287));
    Sp12to4 I__16531 (
            .O(N__67345),
            .I(N__67282));
    Sp12to4 I__16530 (
            .O(N__67340),
            .I(N__67282));
    InMux I__16529 (
            .O(N__67339),
            .I(N__67279));
    LocalMux I__16528 (
            .O(N__67334),
            .I(N__67272));
    Span4Mux_h I__16527 (
            .O(N__67331),
            .I(N__67272));
    Span4Mux_h I__16526 (
            .O(N__67326),
            .I(N__67272));
    LocalMux I__16525 (
            .O(N__67323),
            .I(N__67269));
    Span4Mux_h I__16524 (
            .O(N__67320),
            .I(N__67262));
    Span4Mux_h I__16523 (
            .O(N__67317),
            .I(N__67262));
    Span4Mux_v I__16522 (
            .O(N__67312),
            .I(N__67262));
    LocalMux I__16521 (
            .O(N__67307),
            .I(N__67251));
    LocalMux I__16520 (
            .O(N__67304),
            .I(N__67251));
    LocalMux I__16519 (
            .O(N__67301),
            .I(N__67251));
    Sp12to4 I__16518 (
            .O(N__67296),
            .I(N__67251));
    Span12Mux_v I__16517 (
            .O(N__67293),
            .I(N__67251));
    LocalMux I__16516 (
            .O(N__67290),
            .I(N__67240));
    LocalMux I__16515 (
            .O(N__67287),
            .I(N__67240));
    Span12Mux_h I__16514 (
            .O(N__67282),
            .I(N__67240));
    LocalMux I__16513 (
            .O(N__67279),
            .I(N__67240));
    Sp12to4 I__16512 (
            .O(N__67272),
            .I(N__67240));
    Span4Mux_h I__16511 (
            .O(N__67269),
            .I(N__67237));
    Span4Mux_h I__16510 (
            .O(N__67262),
            .I(N__67234));
    Span12Mux_v I__16509 (
            .O(N__67251),
            .I(N__67231));
    Span12Mux_v I__16508 (
            .O(N__67240),
            .I(N__67228));
    Odrv4 I__16507 (
            .O(N__67237),
            .I(\c0.n9 ));
    Odrv4 I__16506 (
            .O(N__67234),
            .I(\c0.n9 ));
    Odrv12 I__16505 (
            .O(N__67231),
            .I(\c0.n9 ));
    Odrv12 I__16504 (
            .O(N__67228),
            .I(\c0.n9 ));
    InMux I__16503 (
            .O(N__67219),
            .I(N__67211));
    InMux I__16502 (
            .O(N__67218),
            .I(N__67203));
    InMux I__16501 (
            .O(N__67217),
            .I(N__67196));
    InMux I__16500 (
            .O(N__67216),
            .I(N__67196));
    InMux I__16499 (
            .O(N__67215),
            .I(N__67193));
    InMux I__16498 (
            .O(N__67214),
            .I(N__67190));
    LocalMux I__16497 (
            .O(N__67211),
            .I(N__67187));
    CascadeMux I__16496 (
            .O(N__67210),
            .I(N__67183));
    CascadeMux I__16495 (
            .O(N__67209),
            .I(N__67180));
    CascadeMux I__16494 (
            .O(N__67208),
            .I(N__67177));
    InMux I__16493 (
            .O(N__67207),
            .I(N__67172));
    InMux I__16492 (
            .O(N__67206),
            .I(N__67172));
    LocalMux I__16491 (
            .O(N__67203),
            .I(N__67167));
    InMux I__16490 (
            .O(N__67202),
            .I(N__67164));
    InMux I__16489 (
            .O(N__67201),
            .I(N__67158));
    LocalMux I__16488 (
            .O(N__67196),
            .I(N__67154));
    LocalMux I__16487 (
            .O(N__67193),
            .I(N__67149));
    LocalMux I__16486 (
            .O(N__67190),
            .I(N__67149));
    Span4Mux_v I__16485 (
            .O(N__67187),
            .I(N__67146));
    InMux I__16484 (
            .O(N__67186),
            .I(N__67143));
    InMux I__16483 (
            .O(N__67183),
            .I(N__67139));
    InMux I__16482 (
            .O(N__67180),
            .I(N__67134));
    InMux I__16481 (
            .O(N__67177),
            .I(N__67134));
    LocalMux I__16480 (
            .O(N__67172),
            .I(N__67131));
    InMux I__16479 (
            .O(N__67171),
            .I(N__67128));
    InMux I__16478 (
            .O(N__67170),
            .I(N__67125));
    Span4Mux_v I__16477 (
            .O(N__67167),
            .I(N__67117));
    LocalMux I__16476 (
            .O(N__67164),
            .I(N__67117));
    InMux I__16475 (
            .O(N__67163),
            .I(N__67114));
    InMux I__16474 (
            .O(N__67162),
            .I(N__67111));
    InMux I__16473 (
            .O(N__67161),
            .I(N__67108));
    LocalMux I__16472 (
            .O(N__67158),
            .I(N__67105));
    InMux I__16471 (
            .O(N__67157),
            .I(N__67100));
    Span4Mux_v I__16470 (
            .O(N__67154),
            .I(N__67097));
    Span4Mux_v I__16469 (
            .O(N__67149),
            .I(N__67094));
    Span4Mux_h I__16468 (
            .O(N__67146),
            .I(N__67089));
    LocalMux I__16467 (
            .O(N__67143),
            .I(N__67089));
    InMux I__16466 (
            .O(N__67142),
            .I(N__67086));
    LocalMux I__16465 (
            .O(N__67139),
            .I(N__67083));
    LocalMux I__16464 (
            .O(N__67134),
            .I(N__67080));
    Span4Mux_v I__16463 (
            .O(N__67131),
            .I(N__67076));
    LocalMux I__16462 (
            .O(N__67128),
            .I(N__67071));
    LocalMux I__16461 (
            .O(N__67125),
            .I(N__67071));
    InMux I__16460 (
            .O(N__67124),
            .I(N__67067));
    InMux I__16459 (
            .O(N__67123),
            .I(N__67064));
    InMux I__16458 (
            .O(N__67122),
            .I(N__67060));
    Span4Mux_h I__16457 (
            .O(N__67117),
            .I(N__67057));
    LocalMux I__16456 (
            .O(N__67114),
            .I(N__67054));
    LocalMux I__16455 (
            .O(N__67111),
            .I(N__67051));
    LocalMux I__16454 (
            .O(N__67108),
            .I(N__67046));
    Span4Mux_h I__16453 (
            .O(N__67105),
            .I(N__67046));
    InMux I__16452 (
            .O(N__67104),
            .I(N__67043));
    InMux I__16451 (
            .O(N__67103),
            .I(N__67040));
    LocalMux I__16450 (
            .O(N__67100),
            .I(N__67033));
    Span4Mux_h I__16449 (
            .O(N__67097),
            .I(N__67033));
    Span4Mux_h I__16448 (
            .O(N__67094),
            .I(N__67033));
    Span4Mux_h I__16447 (
            .O(N__67089),
            .I(N__67030));
    LocalMux I__16446 (
            .O(N__67086),
            .I(N__67027));
    Span4Mux_v I__16445 (
            .O(N__67083),
            .I(N__67022));
    Span4Mux_v I__16444 (
            .O(N__67080),
            .I(N__67022));
    InMux I__16443 (
            .O(N__67079),
            .I(N__67019));
    Span4Mux_h I__16442 (
            .O(N__67076),
            .I(N__67014));
    Span4Mux_v I__16441 (
            .O(N__67071),
            .I(N__67014));
    InMux I__16440 (
            .O(N__67070),
            .I(N__67011));
    LocalMux I__16439 (
            .O(N__67067),
            .I(N__67006));
    LocalMux I__16438 (
            .O(N__67064),
            .I(N__67006));
    InMux I__16437 (
            .O(N__67063),
            .I(N__67002));
    LocalMux I__16436 (
            .O(N__67060),
            .I(N__66991));
    Span4Mux_v I__16435 (
            .O(N__67057),
            .I(N__66991));
    Span4Mux_v I__16434 (
            .O(N__67054),
            .I(N__66991));
    Span4Mux_v I__16433 (
            .O(N__67051),
            .I(N__66991));
    Span4Mux_h I__16432 (
            .O(N__67046),
            .I(N__66991));
    LocalMux I__16431 (
            .O(N__67043),
            .I(N__66982));
    LocalMux I__16430 (
            .O(N__67040),
            .I(N__66982));
    Span4Mux_h I__16429 (
            .O(N__67033),
            .I(N__66982));
    Span4Mux_v I__16428 (
            .O(N__67030),
            .I(N__66982));
    Sp12to4 I__16427 (
            .O(N__67027),
            .I(N__66979));
    Sp12to4 I__16426 (
            .O(N__67022),
            .I(N__66976));
    LocalMux I__16425 (
            .O(N__67019),
            .I(N__66971));
    Sp12to4 I__16424 (
            .O(N__67014),
            .I(N__66968));
    LocalMux I__16423 (
            .O(N__67011),
            .I(N__66963));
    Sp12to4 I__16422 (
            .O(N__67006),
            .I(N__66963));
    InMux I__16421 (
            .O(N__67005),
            .I(N__66960));
    LocalMux I__16420 (
            .O(N__67002),
            .I(N__66953));
    Span4Mux_h I__16419 (
            .O(N__66991),
            .I(N__66953));
    Span4Mux_v I__16418 (
            .O(N__66982),
            .I(N__66953));
    Span12Mux_s10_v I__16417 (
            .O(N__66979),
            .I(N__66948));
    Span12Mux_h I__16416 (
            .O(N__66976),
            .I(N__66948));
    InMux I__16415 (
            .O(N__66975),
            .I(N__66945));
    InMux I__16414 (
            .O(N__66974),
            .I(N__66942));
    Span4Mux_v I__16413 (
            .O(N__66971),
            .I(N__66939));
    Span12Mux_s9_h I__16412 (
            .O(N__66968),
            .I(N__66934));
    Span12Mux_v I__16411 (
            .O(N__66963),
            .I(N__66934));
    LocalMux I__16410 (
            .O(N__66960),
            .I(N__66929));
    Span4Mux_v I__16409 (
            .O(N__66953),
            .I(N__66929));
    Span12Mux_v I__16408 (
            .O(N__66948),
            .I(N__66926));
    LocalMux I__16407 (
            .O(N__66945),
            .I(rx_data_5));
    LocalMux I__16406 (
            .O(N__66942),
            .I(rx_data_5));
    Odrv4 I__16405 (
            .O(N__66939),
            .I(rx_data_5));
    Odrv12 I__16404 (
            .O(N__66934),
            .I(rx_data_5));
    Odrv4 I__16403 (
            .O(N__66929),
            .I(rx_data_5));
    Odrv12 I__16402 (
            .O(N__66926),
            .I(rx_data_5));
    CascadeMux I__16401 (
            .O(N__66913),
            .I(N__66909));
    CascadeMux I__16400 (
            .O(N__66912),
            .I(N__66905));
    InMux I__16399 (
            .O(N__66909),
            .I(N__66902));
    InMux I__16398 (
            .O(N__66908),
            .I(N__66899));
    InMux I__16397 (
            .O(N__66905),
            .I(N__66896));
    LocalMux I__16396 (
            .O(N__66902),
            .I(N__66893));
    LocalMux I__16395 (
            .O(N__66899),
            .I(N__66890));
    LocalMux I__16394 (
            .O(N__66896),
            .I(N__66883));
    Span4Mux_h I__16393 (
            .O(N__66893),
            .I(N__66883));
    Span4Mux_h I__16392 (
            .O(N__66890),
            .I(N__66883));
    Odrv4 I__16391 (
            .O(N__66883),
            .I(\c0.data_in_frame_27_5 ));
    InMux I__16390 (
            .O(N__66880),
            .I(N__66877));
    LocalMux I__16389 (
            .O(N__66877),
            .I(N__66872));
    ClkMux I__16388 (
            .O(N__66876),
            .I(N__66139));
    ClkMux I__16387 (
            .O(N__66875),
            .I(N__66139));
    Glb2LocalMux I__16386 (
            .O(N__66872),
            .I(N__66139));
    ClkMux I__16385 (
            .O(N__66871),
            .I(N__66139));
    ClkMux I__16384 (
            .O(N__66870),
            .I(N__66139));
    ClkMux I__16383 (
            .O(N__66869),
            .I(N__66139));
    ClkMux I__16382 (
            .O(N__66868),
            .I(N__66139));
    ClkMux I__16381 (
            .O(N__66867),
            .I(N__66139));
    ClkMux I__16380 (
            .O(N__66866),
            .I(N__66139));
    ClkMux I__16379 (
            .O(N__66865),
            .I(N__66139));
    ClkMux I__16378 (
            .O(N__66864),
            .I(N__66139));
    ClkMux I__16377 (
            .O(N__66863),
            .I(N__66139));
    ClkMux I__16376 (
            .O(N__66862),
            .I(N__66139));
    ClkMux I__16375 (
            .O(N__66861),
            .I(N__66139));
    ClkMux I__16374 (
            .O(N__66860),
            .I(N__66139));
    ClkMux I__16373 (
            .O(N__66859),
            .I(N__66139));
    ClkMux I__16372 (
            .O(N__66858),
            .I(N__66139));
    ClkMux I__16371 (
            .O(N__66857),
            .I(N__66139));
    ClkMux I__16370 (
            .O(N__66856),
            .I(N__66139));
    ClkMux I__16369 (
            .O(N__66855),
            .I(N__66139));
    ClkMux I__16368 (
            .O(N__66854),
            .I(N__66139));
    ClkMux I__16367 (
            .O(N__66853),
            .I(N__66139));
    ClkMux I__16366 (
            .O(N__66852),
            .I(N__66139));
    ClkMux I__16365 (
            .O(N__66851),
            .I(N__66139));
    ClkMux I__16364 (
            .O(N__66850),
            .I(N__66139));
    ClkMux I__16363 (
            .O(N__66849),
            .I(N__66139));
    ClkMux I__16362 (
            .O(N__66848),
            .I(N__66139));
    ClkMux I__16361 (
            .O(N__66847),
            .I(N__66139));
    ClkMux I__16360 (
            .O(N__66846),
            .I(N__66139));
    ClkMux I__16359 (
            .O(N__66845),
            .I(N__66139));
    ClkMux I__16358 (
            .O(N__66844),
            .I(N__66139));
    ClkMux I__16357 (
            .O(N__66843),
            .I(N__66139));
    ClkMux I__16356 (
            .O(N__66842),
            .I(N__66139));
    ClkMux I__16355 (
            .O(N__66841),
            .I(N__66139));
    ClkMux I__16354 (
            .O(N__66840),
            .I(N__66139));
    ClkMux I__16353 (
            .O(N__66839),
            .I(N__66139));
    ClkMux I__16352 (
            .O(N__66838),
            .I(N__66139));
    ClkMux I__16351 (
            .O(N__66837),
            .I(N__66139));
    ClkMux I__16350 (
            .O(N__66836),
            .I(N__66139));
    ClkMux I__16349 (
            .O(N__66835),
            .I(N__66139));
    ClkMux I__16348 (
            .O(N__66834),
            .I(N__66139));
    ClkMux I__16347 (
            .O(N__66833),
            .I(N__66139));
    ClkMux I__16346 (
            .O(N__66832),
            .I(N__66139));
    ClkMux I__16345 (
            .O(N__66831),
            .I(N__66139));
    ClkMux I__16344 (
            .O(N__66830),
            .I(N__66139));
    ClkMux I__16343 (
            .O(N__66829),
            .I(N__66139));
    ClkMux I__16342 (
            .O(N__66828),
            .I(N__66139));
    ClkMux I__16341 (
            .O(N__66827),
            .I(N__66139));
    ClkMux I__16340 (
            .O(N__66826),
            .I(N__66139));
    ClkMux I__16339 (
            .O(N__66825),
            .I(N__66139));
    ClkMux I__16338 (
            .O(N__66824),
            .I(N__66139));
    ClkMux I__16337 (
            .O(N__66823),
            .I(N__66139));
    ClkMux I__16336 (
            .O(N__66822),
            .I(N__66139));
    ClkMux I__16335 (
            .O(N__66821),
            .I(N__66139));
    ClkMux I__16334 (
            .O(N__66820),
            .I(N__66139));
    ClkMux I__16333 (
            .O(N__66819),
            .I(N__66139));
    ClkMux I__16332 (
            .O(N__66818),
            .I(N__66139));
    ClkMux I__16331 (
            .O(N__66817),
            .I(N__66139));
    ClkMux I__16330 (
            .O(N__66816),
            .I(N__66139));
    ClkMux I__16329 (
            .O(N__66815),
            .I(N__66139));
    ClkMux I__16328 (
            .O(N__66814),
            .I(N__66139));
    ClkMux I__16327 (
            .O(N__66813),
            .I(N__66139));
    ClkMux I__16326 (
            .O(N__66812),
            .I(N__66139));
    ClkMux I__16325 (
            .O(N__66811),
            .I(N__66139));
    ClkMux I__16324 (
            .O(N__66810),
            .I(N__66139));
    ClkMux I__16323 (
            .O(N__66809),
            .I(N__66139));
    ClkMux I__16322 (
            .O(N__66808),
            .I(N__66139));
    ClkMux I__16321 (
            .O(N__66807),
            .I(N__66139));
    ClkMux I__16320 (
            .O(N__66806),
            .I(N__66139));
    ClkMux I__16319 (
            .O(N__66805),
            .I(N__66139));
    ClkMux I__16318 (
            .O(N__66804),
            .I(N__66139));
    ClkMux I__16317 (
            .O(N__66803),
            .I(N__66139));
    ClkMux I__16316 (
            .O(N__66802),
            .I(N__66139));
    ClkMux I__16315 (
            .O(N__66801),
            .I(N__66139));
    ClkMux I__16314 (
            .O(N__66800),
            .I(N__66139));
    ClkMux I__16313 (
            .O(N__66799),
            .I(N__66139));
    ClkMux I__16312 (
            .O(N__66798),
            .I(N__66139));
    ClkMux I__16311 (
            .O(N__66797),
            .I(N__66139));
    ClkMux I__16310 (
            .O(N__66796),
            .I(N__66139));
    ClkMux I__16309 (
            .O(N__66795),
            .I(N__66139));
    ClkMux I__16308 (
            .O(N__66794),
            .I(N__66139));
    ClkMux I__16307 (
            .O(N__66793),
            .I(N__66139));
    ClkMux I__16306 (
            .O(N__66792),
            .I(N__66139));
    ClkMux I__16305 (
            .O(N__66791),
            .I(N__66139));
    ClkMux I__16304 (
            .O(N__66790),
            .I(N__66139));
    ClkMux I__16303 (
            .O(N__66789),
            .I(N__66139));
    ClkMux I__16302 (
            .O(N__66788),
            .I(N__66139));
    ClkMux I__16301 (
            .O(N__66787),
            .I(N__66139));
    ClkMux I__16300 (
            .O(N__66786),
            .I(N__66139));
    ClkMux I__16299 (
            .O(N__66785),
            .I(N__66139));
    ClkMux I__16298 (
            .O(N__66784),
            .I(N__66139));
    ClkMux I__16297 (
            .O(N__66783),
            .I(N__66139));
    ClkMux I__16296 (
            .O(N__66782),
            .I(N__66139));
    ClkMux I__16295 (
            .O(N__66781),
            .I(N__66139));
    ClkMux I__16294 (
            .O(N__66780),
            .I(N__66139));
    ClkMux I__16293 (
            .O(N__66779),
            .I(N__66139));
    ClkMux I__16292 (
            .O(N__66778),
            .I(N__66139));
    ClkMux I__16291 (
            .O(N__66777),
            .I(N__66139));
    ClkMux I__16290 (
            .O(N__66776),
            .I(N__66139));
    ClkMux I__16289 (
            .O(N__66775),
            .I(N__66139));
    ClkMux I__16288 (
            .O(N__66774),
            .I(N__66139));
    ClkMux I__16287 (
            .O(N__66773),
            .I(N__66139));
    ClkMux I__16286 (
            .O(N__66772),
            .I(N__66139));
    ClkMux I__16285 (
            .O(N__66771),
            .I(N__66139));
    ClkMux I__16284 (
            .O(N__66770),
            .I(N__66139));
    ClkMux I__16283 (
            .O(N__66769),
            .I(N__66139));
    ClkMux I__16282 (
            .O(N__66768),
            .I(N__66139));
    ClkMux I__16281 (
            .O(N__66767),
            .I(N__66139));
    ClkMux I__16280 (
            .O(N__66766),
            .I(N__66139));
    ClkMux I__16279 (
            .O(N__66765),
            .I(N__66139));
    ClkMux I__16278 (
            .O(N__66764),
            .I(N__66139));
    ClkMux I__16277 (
            .O(N__66763),
            .I(N__66139));
    ClkMux I__16276 (
            .O(N__66762),
            .I(N__66139));
    ClkMux I__16275 (
            .O(N__66761),
            .I(N__66139));
    ClkMux I__16274 (
            .O(N__66760),
            .I(N__66139));
    ClkMux I__16273 (
            .O(N__66759),
            .I(N__66139));
    ClkMux I__16272 (
            .O(N__66758),
            .I(N__66139));
    ClkMux I__16271 (
            .O(N__66757),
            .I(N__66139));
    ClkMux I__16270 (
            .O(N__66756),
            .I(N__66139));
    ClkMux I__16269 (
            .O(N__66755),
            .I(N__66139));
    ClkMux I__16268 (
            .O(N__66754),
            .I(N__66139));
    ClkMux I__16267 (
            .O(N__66753),
            .I(N__66139));
    ClkMux I__16266 (
            .O(N__66752),
            .I(N__66139));
    ClkMux I__16265 (
            .O(N__66751),
            .I(N__66139));
    ClkMux I__16264 (
            .O(N__66750),
            .I(N__66139));
    ClkMux I__16263 (
            .O(N__66749),
            .I(N__66139));
    ClkMux I__16262 (
            .O(N__66748),
            .I(N__66139));
    ClkMux I__16261 (
            .O(N__66747),
            .I(N__66139));
    ClkMux I__16260 (
            .O(N__66746),
            .I(N__66139));
    ClkMux I__16259 (
            .O(N__66745),
            .I(N__66139));
    ClkMux I__16258 (
            .O(N__66744),
            .I(N__66139));
    ClkMux I__16257 (
            .O(N__66743),
            .I(N__66139));
    ClkMux I__16256 (
            .O(N__66742),
            .I(N__66139));
    ClkMux I__16255 (
            .O(N__66741),
            .I(N__66139));
    ClkMux I__16254 (
            .O(N__66740),
            .I(N__66139));
    ClkMux I__16253 (
            .O(N__66739),
            .I(N__66139));
    ClkMux I__16252 (
            .O(N__66738),
            .I(N__66139));
    ClkMux I__16251 (
            .O(N__66737),
            .I(N__66139));
    ClkMux I__16250 (
            .O(N__66736),
            .I(N__66139));
    ClkMux I__16249 (
            .O(N__66735),
            .I(N__66139));
    ClkMux I__16248 (
            .O(N__66734),
            .I(N__66139));
    ClkMux I__16247 (
            .O(N__66733),
            .I(N__66139));
    ClkMux I__16246 (
            .O(N__66732),
            .I(N__66139));
    ClkMux I__16245 (
            .O(N__66731),
            .I(N__66139));
    ClkMux I__16244 (
            .O(N__66730),
            .I(N__66139));
    ClkMux I__16243 (
            .O(N__66729),
            .I(N__66139));
    ClkMux I__16242 (
            .O(N__66728),
            .I(N__66139));
    ClkMux I__16241 (
            .O(N__66727),
            .I(N__66139));
    ClkMux I__16240 (
            .O(N__66726),
            .I(N__66139));
    ClkMux I__16239 (
            .O(N__66725),
            .I(N__66139));
    ClkMux I__16238 (
            .O(N__66724),
            .I(N__66139));
    ClkMux I__16237 (
            .O(N__66723),
            .I(N__66139));
    ClkMux I__16236 (
            .O(N__66722),
            .I(N__66139));
    ClkMux I__16235 (
            .O(N__66721),
            .I(N__66139));
    ClkMux I__16234 (
            .O(N__66720),
            .I(N__66139));
    ClkMux I__16233 (
            .O(N__66719),
            .I(N__66139));
    ClkMux I__16232 (
            .O(N__66718),
            .I(N__66139));
    ClkMux I__16231 (
            .O(N__66717),
            .I(N__66139));
    ClkMux I__16230 (
            .O(N__66716),
            .I(N__66139));
    ClkMux I__16229 (
            .O(N__66715),
            .I(N__66139));
    ClkMux I__16228 (
            .O(N__66714),
            .I(N__66139));
    ClkMux I__16227 (
            .O(N__66713),
            .I(N__66139));
    ClkMux I__16226 (
            .O(N__66712),
            .I(N__66139));
    ClkMux I__16225 (
            .O(N__66711),
            .I(N__66139));
    ClkMux I__16224 (
            .O(N__66710),
            .I(N__66139));
    ClkMux I__16223 (
            .O(N__66709),
            .I(N__66139));
    ClkMux I__16222 (
            .O(N__66708),
            .I(N__66139));
    ClkMux I__16221 (
            .O(N__66707),
            .I(N__66139));
    ClkMux I__16220 (
            .O(N__66706),
            .I(N__66139));
    ClkMux I__16219 (
            .O(N__66705),
            .I(N__66139));
    ClkMux I__16218 (
            .O(N__66704),
            .I(N__66139));
    ClkMux I__16217 (
            .O(N__66703),
            .I(N__66139));
    ClkMux I__16216 (
            .O(N__66702),
            .I(N__66139));
    ClkMux I__16215 (
            .O(N__66701),
            .I(N__66139));
    ClkMux I__16214 (
            .O(N__66700),
            .I(N__66139));
    ClkMux I__16213 (
            .O(N__66699),
            .I(N__66139));
    ClkMux I__16212 (
            .O(N__66698),
            .I(N__66139));
    ClkMux I__16211 (
            .O(N__66697),
            .I(N__66139));
    ClkMux I__16210 (
            .O(N__66696),
            .I(N__66139));
    ClkMux I__16209 (
            .O(N__66695),
            .I(N__66139));
    ClkMux I__16208 (
            .O(N__66694),
            .I(N__66139));
    ClkMux I__16207 (
            .O(N__66693),
            .I(N__66139));
    ClkMux I__16206 (
            .O(N__66692),
            .I(N__66139));
    ClkMux I__16205 (
            .O(N__66691),
            .I(N__66139));
    ClkMux I__16204 (
            .O(N__66690),
            .I(N__66139));
    ClkMux I__16203 (
            .O(N__66689),
            .I(N__66139));
    ClkMux I__16202 (
            .O(N__66688),
            .I(N__66139));
    ClkMux I__16201 (
            .O(N__66687),
            .I(N__66139));
    ClkMux I__16200 (
            .O(N__66686),
            .I(N__66139));
    ClkMux I__16199 (
            .O(N__66685),
            .I(N__66139));
    ClkMux I__16198 (
            .O(N__66684),
            .I(N__66139));
    ClkMux I__16197 (
            .O(N__66683),
            .I(N__66139));
    ClkMux I__16196 (
            .O(N__66682),
            .I(N__66139));
    ClkMux I__16195 (
            .O(N__66681),
            .I(N__66139));
    ClkMux I__16194 (
            .O(N__66680),
            .I(N__66139));
    ClkMux I__16193 (
            .O(N__66679),
            .I(N__66139));
    ClkMux I__16192 (
            .O(N__66678),
            .I(N__66139));
    ClkMux I__16191 (
            .O(N__66677),
            .I(N__66139));
    ClkMux I__16190 (
            .O(N__66676),
            .I(N__66139));
    ClkMux I__16189 (
            .O(N__66675),
            .I(N__66139));
    ClkMux I__16188 (
            .O(N__66674),
            .I(N__66139));
    ClkMux I__16187 (
            .O(N__66673),
            .I(N__66139));
    ClkMux I__16186 (
            .O(N__66672),
            .I(N__66139));
    ClkMux I__16185 (
            .O(N__66671),
            .I(N__66139));
    ClkMux I__16184 (
            .O(N__66670),
            .I(N__66139));
    ClkMux I__16183 (
            .O(N__66669),
            .I(N__66139));
    ClkMux I__16182 (
            .O(N__66668),
            .I(N__66139));
    ClkMux I__16181 (
            .O(N__66667),
            .I(N__66139));
    ClkMux I__16180 (
            .O(N__66666),
            .I(N__66139));
    ClkMux I__16179 (
            .O(N__66665),
            .I(N__66139));
    ClkMux I__16178 (
            .O(N__66664),
            .I(N__66139));
    ClkMux I__16177 (
            .O(N__66663),
            .I(N__66139));
    ClkMux I__16176 (
            .O(N__66662),
            .I(N__66139));
    ClkMux I__16175 (
            .O(N__66661),
            .I(N__66139));
    ClkMux I__16174 (
            .O(N__66660),
            .I(N__66139));
    ClkMux I__16173 (
            .O(N__66659),
            .I(N__66139));
    ClkMux I__16172 (
            .O(N__66658),
            .I(N__66139));
    ClkMux I__16171 (
            .O(N__66657),
            .I(N__66139));
    ClkMux I__16170 (
            .O(N__66656),
            .I(N__66139));
    ClkMux I__16169 (
            .O(N__66655),
            .I(N__66139));
    ClkMux I__16168 (
            .O(N__66654),
            .I(N__66139));
    ClkMux I__16167 (
            .O(N__66653),
            .I(N__66139));
    ClkMux I__16166 (
            .O(N__66652),
            .I(N__66139));
    ClkMux I__16165 (
            .O(N__66651),
            .I(N__66139));
    ClkMux I__16164 (
            .O(N__66650),
            .I(N__66139));
    ClkMux I__16163 (
            .O(N__66649),
            .I(N__66139));
    ClkMux I__16162 (
            .O(N__66648),
            .I(N__66139));
    ClkMux I__16161 (
            .O(N__66647),
            .I(N__66139));
    ClkMux I__16160 (
            .O(N__66646),
            .I(N__66139));
    ClkMux I__16159 (
            .O(N__66645),
            .I(N__66139));
    ClkMux I__16158 (
            .O(N__66644),
            .I(N__66139));
    ClkMux I__16157 (
            .O(N__66643),
            .I(N__66139));
    ClkMux I__16156 (
            .O(N__66642),
            .I(N__66139));
    ClkMux I__16155 (
            .O(N__66641),
            .I(N__66139));
    ClkMux I__16154 (
            .O(N__66640),
            .I(N__66139));
    ClkMux I__16153 (
            .O(N__66639),
            .I(N__66139));
    ClkMux I__16152 (
            .O(N__66638),
            .I(N__66139));
    ClkMux I__16151 (
            .O(N__66637),
            .I(N__66139));
    ClkMux I__16150 (
            .O(N__66636),
            .I(N__66139));
    ClkMux I__16149 (
            .O(N__66635),
            .I(N__66139));
    ClkMux I__16148 (
            .O(N__66634),
            .I(N__66139));
    ClkMux I__16147 (
            .O(N__66633),
            .I(N__66139));
    ClkMux I__16146 (
            .O(N__66632),
            .I(N__66139));
    ClkMux I__16145 (
            .O(N__66631),
            .I(N__66139));
    ClkMux I__16144 (
            .O(N__66630),
            .I(N__66139));
    GlobalMux I__16143 (
            .O(N__66139),
            .I(PIN_9_c));
    InMux I__16142 (
            .O(N__66136),
            .I(N__66132));
    InMux I__16141 (
            .O(N__66135),
            .I(N__66129));
    LocalMux I__16140 (
            .O(N__66132),
            .I(N__66125));
    LocalMux I__16139 (
            .O(N__66129),
            .I(N__66121));
    InMux I__16138 (
            .O(N__66128),
            .I(N__66118));
    Span4Mux_h I__16137 (
            .O(N__66125),
            .I(N__66115));
    InMux I__16136 (
            .O(N__66124),
            .I(N__66112));
    Span4Mux_h I__16135 (
            .O(N__66121),
            .I(N__66107));
    LocalMux I__16134 (
            .O(N__66118),
            .I(N__66107));
    Span4Mux_h I__16133 (
            .O(N__66115),
            .I(N__66104));
    LocalMux I__16132 (
            .O(N__66112),
            .I(\c0.data_in_frame_27_7 ));
    Odrv4 I__16131 (
            .O(N__66107),
            .I(\c0.data_in_frame_27_7 ));
    Odrv4 I__16130 (
            .O(N__66104),
            .I(\c0.data_in_frame_27_7 ));
    InMux I__16129 (
            .O(N__66097),
            .I(N__66092));
    CascadeMux I__16128 (
            .O(N__66096),
            .I(N__66089));
    CascadeMux I__16127 (
            .O(N__66095),
            .I(N__66086));
    LocalMux I__16126 (
            .O(N__66092),
            .I(N__66083));
    InMux I__16125 (
            .O(N__66089),
            .I(N__66080));
    InMux I__16124 (
            .O(N__66086),
            .I(N__66077));
    Span4Mux_h I__16123 (
            .O(N__66083),
            .I(N__66072));
    LocalMux I__16122 (
            .O(N__66080),
            .I(N__66072));
    LocalMux I__16121 (
            .O(N__66077),
            .I(\c0.data_in_frame_27_6 ));
    Odrv4 I__16120 (
            .O(N__66072),
            .I(\c0.data_in_frame_27_6 ));
    InMux I__16119 (
            .O(N__66067),
            .I(N__66060));
    InMux I__16118 (
            .O(N__66066),
            .I(N__66060));
    InMux I__16117 (
            .O(N__66065),
            .I(N__66057));
    LocalMux I__16116 (
            .O(N__66060),
            .I(N__66054));
    LocalMux I__16115 (
            .O(N__66057),
            .I(\c0.data_in_frame_27_0 ));
    Odrv4 I__16114 (
            .O(N__66054),
            .I(\c0.data_in_frame_27_0 ));
    InMux I__16113 (
            .O(N__66049),
            .I(N__66045));
    InMux I__16112 (
            .O(N__66048),
            .I(N__66042));
    LocalMux I__16111 (
            .O(N__66045),
            .I(N__66039));
    LocalMux I__16110 (
            .O(N__66042),
            .I(N__66034));
    Span4Mux_h I__16109 (
            .O(N__66039),
            .I(N__66034));
    Odrv4 I__16108 (
            .O(N__66034),
            .I(\c0.n6268 ));
    InMux I__16107 (
            .O(N__66031),
            .I(N__66025));
    InMux I__16106 (
            .O(N__66030),
            .I(N__66022));
    CascadeMux I__16105 (
            .O(N__66029),
            .I(N__66016));
    CascadeMux I__16104 (
            .O(N__66028),
            .I(N__66009));
    LocalMux I__16103 (
            .O(N__66025),
            .I(N__66004));
    LocalMux I__16102 (
            .O(N__66022),
            .I(N__65998));
    InMux I__16101 (
            .O(N__66021),
            .I(N__65993));
    InMux I__16100 (
            .O(N__66020),
            .I(N__65993));
    CascadeMux I__16099 (
            .O(N__66019),
            .I(N__65988));
    InMux I__16098 (
            .O(N__66016),
            .I(N__65985));
    CascadeMux I__16097 (
            .O(N__66015),
            .I(N__65982));
    InMux I__16096 (
            .O(N__66014),
            .I(N__65977));
    InMux I__16095 (
            .O(N__66013),
            .I(N__65977));
    CascadeMux I__16094 (
            .O(N__66012),
            .I(N__65974));
    InMux I__16093 (
            .O(N__66009),
            .I(N__65964));
    InMux I__16092 (
            .O(N__66008),
            .I(N__65964));
    InMux I__16091 (
            .O(N__66007),
            .I(N__65961));
    Span4Mux_v I__16090 (
            .O(N__66004),
            .I(N__65958));
    InMux I__16089 (
            .O(N__66003),
            .I(N__65953));
    InMux I__16088 (
            .O(N__66002),
            .I(N__65953));
    InMux I__16087 (
            .O(N__66001),
            .I(N__65950));
    Span4Mux_h I__16086 (
            .O(N__65998),
            .I(N__65944));
    LocalMux I__16085 (
            .O(N__65993),
            .I(N__65944));
    InMux I__16084 (
            .O(N__65992),
            .I(N__65941));
    CascadeMux I__16083 (
            .O(N__65991),
            .I(N__65933));
    InMux I__16082 (
            .O(N__65988),
            .I(N__65929));
    LocalMux I__16081 (
            .O(N__65985),
            .I(N__65926));
    InMux I__16080 (
            .O(N__65982),
            .I(N__65923));
    LocalMux I__16079 (
            .O(N__65977),
            .I(N__65920));
    InMux I__16078 (
            .O(N__65974),
            .I(N__65917));
    InMux I__16077 (
            .O(N__65973),
            .I(N__65908));
    InMux I__16076 (
            .O(N__65972),
            .I(N__65908));
    InMux I__16075 (
            .O(N__65971),
            .I(N__65908));
    InMux I__16074 (
            .O(N__65970),
            .I(N__65908));
    InMux I__16073 (
            .O(N__65969),
            .I(N__65905));
    LocalMux I__16072 (
            .O(N__65964),
            .I(N__65900));
    LocalMux I__16071 (
            .O(N__65961),
            .I(N__65900));
    Span4Mux_h I__16070 (
            .O(N__65958),
            .I(N__65894));
    LocalMux I__16069 (
            .O(N__65953),
            .I(N__65894));
    LocalMux I__16068 (
            .O(N__65950),
            .I(N__65891));
    InMux I__16067 (
            .O(N__65949),
            .I(N__65888));
    Span4Mux_h I__16066 (
            .O(N__65944),
            .I(N__65885));
    LocalMux I__16065 (
            .O(N__65941),
            .I(N__65882));
    InMux I__16064 (
            .O(N__65940),
            .I(N__65879));
    InMux I__16063 (
            .O(N__65939),
            .I(N__65876));
    InMux I__16062 (
            .O(N__65938),
            .I(N__65869));
    InMux I__16061 (
            .O(N__65937),
            .I(N__65869));
    InMux I__16060 (
            .O(N__65936),
            .I(N__65869));
    InMux I__16059 (
            .O(N__65933),
            .I(N__65866));
    InMux I__16058 (
            .O(N__65932),
            .I(N__65862));
    LocalMux I__16057 (
            .O(N__65929),
            .I(N__65859));
    Span4Mux_h I__16056 (
            .O(N__65926),
            .I(N__65850));
    LocalMux I__16055 (
            .O(N__65923),
            .I(N__65850));
    Span4Mux_v I__16054 (
            .O(N__65920),
            .I(N__65850));
    LocalMux I__16053 (
            .O(N__65917),
            .I(N__65850));
    LocalMux I__16052 (
            .O(N__65908),
            .I(N__65847));
    LocalMux I__16051 (
            .O(N__65905),
            .I(N__65842));
    Span4Mux_h I__16050 (
            .O(N__65900),
            .I(N__65842));
    InMux I__16049 (
            .O(N__65899),
            .I(N__65839));
    Span4Mux_v I__16048 (
            .O(N__65894),
            .I(N__65834));
    Span4Mux_v I__16047 (
            .O(N__65891),
            .I(N__65834));
    LocalMux I__16046 (
            .O(N__65888),
            .I(N__65825));
    Span4Mux_v I__16045 (
            .O(N__65885),
            .I(N__65825));
    Span4Mux_h I__16044 (
            .O(N__65882),
            .I(N__65825));
    LocalMux I__16043 (
            .O(N__65879),
            .I(N__65825));
    LocalMux I__16042 (
            .O(N__65876),
            .I(N__65822));
    LocalMux I__16041 (
            .O(N__65869),
            .I(N__65819));
    LocalMux I__16040 (
            .O(N__65866),
            .I(N__65816));
    InMux I__16039 (
            .O(N__65865),
            .I(N__65813));
    LocalMux I__16038 (
            .O(N__65862),
            .I(N__65806));
    Span4Mux_h I__16037 (
            .O(N__65859),
            .I(N__65806));
    Span4Mux_v I__16036 (
            .O(N__65850),
            .I(N__65806));
    Span4Mux_h I__16035 (
            .O(N__65847),
            .I(N__65801));
    Span4Mux_v I__16034 (
            .O(N__65842),
            .I(N__65801));
    LocalMux I__16033 (
            .O(N__65839),
            .I(N__65798));
    Span4Mux_h I__16032 (
            .O(N__65834),
            .I(N__65793));
    Span4Mux_v I__16031 (
            .O(N__65825),
            .I(N__65793));
    Span4Mux_v I__16030 (
            .O(N__65822),
            .I(N__65788));
    Span4Mux_v I__16029 (
            .O(N__65819),
            .I(N__65788));
    Span12Mux_v I__16028 (
            .O(N__65816),
            .I(N__65785));
    LocalMux I__16027 (
            .O(N__65813),
            .I(N__65780));
    Sp12to4 I__16026 (
            .O(N__65806),
            .I(N__65780));
    Span4Mux_v I__16025 (
            .O(N__65801),
            .I(N__65777));
    Span4Mux_v I__16024 (
            .O(N__65798),
            .I(N__65772));
    Span4Mux_h I__16023 (
            .O(N__65793),
            .I(N__65772));
    Odrv4 I__16022 (
            .O(N__65788),
            .I(\c0.n9_adj_4278 ));
    Odrv12 I__16021 (
            .O(N__65785),
            .I(\c0.n9_adj_4278 ));
    Odrv12 I__16020 (
            .O(N__65780),
            .I(\c0.n9_adj_4278 ));
    Odrv4 I__16019 (
            .O(N__65777),
            .I(\c0.n9_adj_4278 ));
    Odrv4 I__16018 (
            .O(N__65772),
            .I(\c0.n9_adj_4278 ));
    InMux I__16017 (
            .O(N__65761),
            .I(N__65756));
    InMux I__16016 (
            .O(N__65760),
            .I(N__65751));
    InMux I__16015 (
            .O(N__65759),
            .I(N__65751));
    LocalMux I__16014 (
            .O(N__65756),
            .I(N__65747));
    LocalMux I__16013 (
            .O(N__65751),
            .I(N__65744));
    CascadeMux I__16012 (
            .O(N__65750),
            .I(N__65741));
    Span4Mux_h I__16011 (
            .O(N__65747),
            .I(N__65738));
    Span4Mux_h I__16010 (
            .O(N__65744),
            .I(N__65735));
    InMux I__16009 (
            .O(N__65741),
            .I(N__65732));
    Span4Mux_v I__16008 (
            .O(N__65738),
            .I(N__65729));
    Span4Mux_v I__16007 (
            .O(N__65735),
            .I(N__65726));
    LocalMux I__16006 (
            .O(N__65732),
            .I(\c0.data_in_frame_16_7 ));
    Odrv4 I__16005 (
            .O(N__65729),
            .I(\c0.data_in_frame_16_7 ));
    Odrv4 I__16004 (
            .O(N__65726),
            .I(\c0.data_in_frame_16_7 ));
    InMux I__16003 (
            .O(N__65719),
            .I(N__65715));
    CascadeMux I__16002 (
            .O(N__65718),
            .I(N__65712));
    LocalMux I__16001 (
            .O(N__65715),
            .I(N__65709));
    InMux I__16000 (
            .O(N__65712),
            .I(N__65706));
    Span4Mux_h I__15999 (
            .O(N__65709),
            .I(N__65703));
    LocalMux I__15998 (
            .O(N__65706),
            .I(\c0.data_in_frame_19_0 ));
    Odrv4 I__15997 (
            .O(N__65703),
            .I(\c0.data_in_frame_19_0 ));
    InMux I__15996 (
            .O(N__65698),
            .I(N__65693));
    InMux I__15995 (
            .O(N__65697),
            .I(N__65690));
    CascadeMux I__15994 (
            .O(N__65696),
            .I(N__65686));
    LocalMux I__15993 (
            .O(N__65693),
            .I(N__65681));
    LocalMux I__15992 (
            .O(N__65690),
            .I(N__65681));
    InMux I__15991 (
            .O(N__65689),
            .I(N__65678));
    InMux I__15990 (
            .O(N__65686),
            .I(N__65675));
    Span4Mux_v I__15989 (
            .O(N__65681),
            .I(N__65667));
    LocalMux I__15988 (
            .O(N__65678),
            .I(N__65662));
    LocalMux I__15987 (
            .O(N__65675),
            .I(N__65662));
    InMux I__15986 (
            .O(N__65674),
            .I(N__65658));
    InMux I__15985 (
            .O(N__65673),
            .I(N__65655));
    InMux I__15984 (
            .O(N__65672),
            .I(N__65650));
    InMux I__15983 (
            .O(N__65671),
            .I(N__65650));
    InMux I__15982 (
            .O(N__65670),
            .I(N__65644));
    Span4Mux_h I__15981 (
            .O(N__65667),
            .I(N__65639));
    Span4Mux_v I__15980 (
            .O(N__65662),
            .I(N__65639));
    InMux I__15979 (
            .O(N__65661),
            .I(N__65636));
    LocalMux I__15978 (
            .O(N__65658),
            .I(N__65631));
    LocalMux I__15977 (
            .O(N__65655),
            .I(N__65631));
    LocalMux I__15976 (
            .O(N__65650),
            .I(N__65628));
    InMux I__15975 (
            .O(N__65649),
            .I(N__65625));
    InMux I__15974 (
            .O(N__65648),
            .I(N__65620));
    CascadeMux I__15973 (
            .O(N__65647),
            .I(N__65617));
    LocalMux I__15972 (
            .O(N__65644),
            .I(N__65604));
    Span4Mux_h I__15971 (
            .O(N__65639),
            .I(N__65604));
    LocalMux I__15970 (
            .O(N__65636),
            .I(N__65604));
    Span4Mux_v I__15969 (
            .O(N__65631),
            .I(N__65604));
    Span4Mux_h I__15968 (
            .O(N__65628),
            .I(N__65604));
    LocalMux I__15967 (
            .O(N__65625),
            .I(N__65604));
    InMux I__15966 (
            .O(N__65624),
            .I(N__65601));
    InMux I__15965 (
            .O(N__65623),
            .I(N__65598));
    LocalMux I__15964 (
            .O(N__65620),
            .I(N__65595));
    InMux I__15963 (
            .O(N__65617),
            .I(N__65592));
    Span4Mux_h I__15962 (
            .O(N__65604),
            .I(N__65588));
    LocalMux I__15961 (
            .O(N__65601),
            .I(N__65583));
    LocalMux I__15960 (
            .O(N__65598),
            .I(N__65583));
    Span4Mux_v I__15959 (
            .O(N__65595),
            .I(N__65577));
    LocalMux I__15958 (
            .O(N__65592),
            .I(N__65577));
    CascadeMux I__15957 (
            .O(N__65591),
            .I(N__65564));
    Span4Mux_v I__15956 (
            .O(N__65588),
            .I(N__65557));
    Span4Mux_v I__15955 (
            .O(N__65583),
            .I(N__65557));
    InMux I__15954 (
            .O(N__65582),
            .I(N__65554));
    Span4Mux_h I__15953 (
            .O(N__65577),
            .I(N__65551));
    InMux I__15952 (
            .O(N__65576),
            .I(N__65548));
    InMux I__15951 (
            .O(N__65575),
            .I(N__65545));
    InMux I__15950 (
            .O(N__65574),
            .I(N__65542));
    InMux I__15949 (
            .O(N__65573),
            .I(N__65537));
    InMux I__15948 (
            .O(N__65572),
            .I(N__65537));
    InMux I__15947 (
            .O(N__65571),
            .I(N__65532));
    InMux I__15946 (
            .O(N__65570),
            .I(N__65532));
    InMux I__15945 (
            .O(N__65569),
            .I(N__65529));
    InMux I__15944 (
            .O(N__65568),
            .I(N__65524));
    InMux I__15943 (
            .O(N__65567),
            .I(N__65524));
    InMux I__15942 (
            .O(N__65564),
            .I(N__65521));
    InMux I__15941 (
            .O(N__65563),
            .I(N__65518));
    InMux I__15940 (
            .O(N__65562),
            .I(N__65515));
    Sp12to4 I__15939 (
            .O(N__65557),
            .I(N__65512));
    LocalMux I__15938 (
            .O(N__65554),
            .I(N__65509));
    Sp12to4 I__15937 (
            .O(N__65551),
            .I(N__65504));
    LocalMux I__15936 (
            .O(N__65548),
            .I(N__65504));
    LocalMux I__15935 (
            .O(N__65545),
            .I(N__65498));
    LocalMux I__15934 (
            .O(N__65542),
            .I(N__65495));
    LocalMux I__15933 (
            .O(N__65537),
            .I(N__65492));
    LocalMux I__15932 (
            .O(N__65532),
            .I(N__65489));
    LocalMux I__15931 (
            .O(N__65529),
            .I(N__65486));
    LocalMux I__15930 (
            .O(N__65524),
            .I(N__65481));
    LocalMux I__15929 (
            .O(N__65521),
            .I(N__65481));
    LocalMux I__15928 (
            .O(N__65518),
            .I(N__65470));
    LocalMux I__15927 (
            .O(N__65515),
            .I(N__65470));
    Span12Mux_h I__15926 (
            .O(N__65512),
            .I(N__65470));
    Span12Mux_h I__15925 (
            .O(N__65509),
            .I(N__65470));
    Span12Mux_s9_v I__15924 (
            .O(N__65504),
            .I(N__65470));
    InMux I__15923 (
            .O(N__65503),
            .I(N__65465));
    InMux I__15922 (
            .O(N__65502),
            .I(N__65465));
    InMux I__15921 (
            .O(N__65501),
            .I(N__65462));
    Span4Mux_h I__15920 (
            .O(N__65498),
            .I(N__65459));
    Span4Mux_v I__15919 (
            .O(N__65495),
            .I(N__65454));
    Span4Mux_v I__15918 (
            .O(N__65492),
            .I(N__65454));
    Span12Mux_v I__15917 (
            .O(N__65489),
            .I(N__65451));
    Span12Mux_v I__15916 (
            .O(N__65486),
            .I(N__65446));
    Span12Mux_h I__15915 (
            .O(N__65481),
            .I(N__65446));
    Span12Mux_v I__15914 (
            .O(N__65470),
            .I(N__65443));
    LocalMux I__15913 (
            .O(N__65465),
            .I(rx_data_6));
    LocalMux I__15912 (
            .O(N__65462),
            .I(rx_data_6));
    Odrv4 I__15911 (
            .O(N__65459),
            .I(rx_data_6));
    Odrv4 I__15910 (
            .O(N__65454),
            .I(rx_data_6));
    Odrv12 I__15909 (
            .O(N__65451),
            .I(rx_data_6));
    Odrv12 I__15908 (
            .O(N__65446),
            .I(rx_data_6));
    Odrv12 I__15907 (
            .O(N__65443),
            .I(rx_data_6));
    InMux I__15906 (
            .O(N__65428),
            .I(N__65425));
    LocalMux I__15905 (
            .O(N__65425),
            .I(N__65421));
    CascadeMux I__15904 (
            .O(N__65424),
            .I(N__65418));
    Span4Mux_h I__15903 (
            .O(N__65421),
            .I(N__65414));
    InMux I__15902 (
            .O(N__65418),
            .I(N__65409));
    InMux I__15901 (
            .O(N__65417),
            .I(N__65409));
    Odrv4 I__15900 (
            .O(N__65414),
            .I(\c0.data_in_frame_18_6 ));
    LocalMux I__15899 (
            .O(N__65409),
            .I(\c0.data_in_frame_18_6 ));
    CascadeMux I__15898 (
            .O(N__65404),
            .I(N__65401));
    InMux I__15897 (
            .O(N__65401),
            .I(N__65397));
    CascadeMux I__15896 (
            .O(N__65400),
            .I(N__65394));
    LocalMux I__15895 (
            .O(N__65397),
            .I(N__65391));
    InMux I__15894 (
            .O(N__65394),
            .I(N__65388));
    Span4Mux_h I__15893 (
            .O(N__65391),
            .I(N__65385));
    LocalMux I__15892 (
            .O(N__65388),
            .I(N__65380));
    Span4Mux_v I__15891 (
            .O(N__65385),
            .I(N__65380));
    Span4Mux_v I__15890 (
            .O(N__65380),
            .I(N__65375));
    InMux I__15889 (
            .O(N__65379),
            .I(N__65370));
    InMux I__15888 (
            .O(N__65378),
            .I(N__65370));
    Odrv4 I__15887 (
            .O(N__65375),
            .I(\c0.data_in_frame_18_7 ));
    LocalMux I__15886 (
            .O(N__65370),
            .I(\c0.data_in_frame_18_7 ));
    InMux I__15885 (
            .O(N__65365),
            .I(N__65361));
    InMux I__15884 (
            .O(N__65364),
            .I(N__65358));
    LocalMux I__15883 (
            .O(N__65361),
            .I(N__65352));
    LocalMux I__15882 (
            .O(N__65358),
            .I(N__65349));
    InMux I__15881 (
            .O(N__65357),
            .I(N__65344));
    InMux I__15880 (
            .O(N__65356),
            .I(N__65344));
    InMux I__15879 (
            .O(N__65355),
            .I(N__65341));
    Span4Mux_v I__15878 (
            .O(N__65352),
            .I(N__65338));
    Span4Mux_h I__15877 (
            .O(N__65349),
            .I(N__65335));
    LocalMux I__15876 (
            .O(N__65344),
            .I(\c0.data_in_frame_21_5 ));
    LocalMux I__15875 (
            .O(N__65341),
            .I(\c0.data_in_frame_21_5 ));
    Odrv4 I__15874 (
            .O(N__65338),
            .I(\c0.data_in_frame_21_5 ));
    Odrv4 I__15873 (
            .O(N__65335),
            .I(\c0.data_in_frame_21_5 ));
    InMux I__15872 (
            .O(N__65326),
            .I(N__65323));
    LocalMux I__15871 (
            .O(N__65323),
            .I(N__65319));
    InMux I__15870 (
            .O(N__65322),
            .I(N__65316));
    Span4Mux_h I__15869 (
            .O(N__65319),
            .I(N__65311));
    LocalMux I__15868 (
            .O(N__65316),
            .I(N__65311));
    Span4Mux_h I__15867 (
            .O(N__65311),
            .I(N__65308));
    Odrv4 I__15866 (
            .O(N__65308),
            .I(\c0.n22123 ));
    InMux I__15865 (
            .O(N__65305),
            .I(N__65301));
    InMux I__15864 (
            .O(N__65304),
            .I(N__65298));
    LocalMux I__15863 (
            .O(N__65301),
            .I(N__65292));
    LocalMux I__15862 (
            .O(N__65298),
            .I(N__65292));
    CascadeMux I__15861 (
            .O(N__65297),
            .I(N__65289));
    Span4Mux_v I__15860 (
            .O(N__65292),
            .I(N__65286));
    InMux I__15859 (
            .O(N__65289),
            .I(N__65283));
    Span4Mux_v I__15858 (
            .O(N__65286),
            .I(N__65280));
    LocalMux I__15857 (
            .O(N__65283),
            .I(\c0.data_in_frame_23_7 ));
    Odrv4 I__15856 (
            .O(N__65280),
            .I(\c0.data_in_frame_23_7 ));
    CascadeMux I__15855 (
            .O(N__65275),
            .I(N__65272));
    InMux I__15854 (
            .O(N__65272),
            .I(N__65269));
    LocalMux I__15853 (
            .O(N__65269),
            .I(N__65266));
    Span4Mux_h I__15852 (
            .O(N__65266),
            .I(N__65262));
    InMux I__15851 (
            .O(N__65265),
            .I(N__65259));
    Sp12to4 I__15850 (
            .O(N__65262),
            .I(N__65256));
    LocalMux I__15849 (
            .O(N__65259),
            .I(N__65253));
    Odrv12 I__15848 (
            .O(N__65256),
            .I(\c0.n22396 ));
    Odrv12 I__15847 (
            .O(N__65253),
            .I(\c0.n22396 ));
    InMux I__15846 (
            .O(N__65248),
            .I(N__65242));
    InMux I__15845 (
            .O(N__65247),
            .I(N__65239));
    InMux I__15844 (
            .O(N__65246),
            .I(N__65234));
    InMux I__15843 (
            .O(N__65245),
            .I(N__65234));
    LocalMux I__15842 (
            .O(N__65242),
            .I(N__65231));
    LocalMux I__15841 (
            .O(N__65239),
            .I(N__65227));
    LocalMux I__15840 (
            .O(N__65234),
            .I(N__65224));
    Span4Mux_h I__15839 (
            .O(N__65231),
            .I(N__65221));
    InMux I__15838 (
            .O(N__65230),
            .I(N__65218));
    Span4Mux_v I__15837 (
            .O(N__65227),
            .I(N__65213));
    Span4Mux_h I__15836 (
            .O(N__65224),
            .I(N__65213));
    Odrv4 I__15835 (
            .O(N__65221),
            .I(\c0.n20288 ));
    LocalMux I__15834 (
            .O(N__65218),
            .I(\c0.n20288 ));
    Odrv4 I__15833 (
            .O(N__65213),
            .I(\c0.n20288 ));
    InMux I__15832 (
            .O(N__65206),
            .I(N__65203));
    LocalMux I__15831 (
            .O(N__65203),
            .I(\c0.n23 ));
    InMux I__15830 (
            .O(N__65200),
            .I(N__65197));
    LocalMux I__15829 (
            .O(N__65197),
            .I(N__65194));
    Span4Mux_v I__15828 (
            .O(N__65194),
            .I(N__65189));
    InMux I__15827 (
            .O(N__65193),
            .I(N__65186));
    CascadeMux I__15826 (
            .O(N__65192),
            .I(N__65183));
    Span4Mux_v I__15825 (
            .O(N__65189),
            .I(N__65180));
    LocalMux I__15824 (
            .O(N__65186),
            .I(N__65176));
    InMux I__15823 (
            .O(N__65183),
            .I(N__65173));
    Span4Mux_h I__15822 (
            .O(N__65180),
            .I(N__65170));
    InMux I__15821 (
            .O(N__65179),
            .I(N__65167));
    Span4Mux_v I__15820 (
            .O(N__65176),
            .I(N__65164));
    LocalMux I__15819 (
            .O(N__65173),
            .I(\c0.data_in_frame_24_2 ));
    Odrv4 I__15818 (
            .O(N__65170),
            .I(\c0.data_in_frame_24_2 ));
    LocalMux I__15817 (
            .O(N__65167),
            .I(\c0.data_in_frame_24_2 ));
    Odrv4 I__15816 (
            .O(N__65164),
            .I(\c0.data_in_frame_24_2 ));
    InMux I__15815 (
            .O(N__65155),
            .I(N__65150));
    InMux I__15814 (
            .O(N__65154),
            .I(N__65147));
    InMux I__15813 (
            .O(N__65153),
            .I(N__65143));
    LocalMux I__15812 (
            .O(N__65150),
            .I(N__65140));
    LocalMux I__15811 (
            .O(N__65147),
            .I(N__65137));
    InMux I__15810 (
            .O(N__65146),
            .I(N__65134));
    LocalMux I__15809 (
            .O(N__65143),
            .I(N__65131));
    Span4Mux_h I__15808 (
            .O(N__65140),
            .I(N__65128));
    Span4Mux_v I__15807 (
            .O(N__65137),
            .I(N__65123));
    LocalMux I__15806 (
            .O(N__65134),
            .I(N__65123));
    Span4Mux_v I__15805 (
            .O(N__65131),
            .I(N__65120));
    Odrv4 I__15804 (
            .O(N__65128),
            .I(\c0.n13443 ));
    Odrv4 I__15803 (
            .O(N__65123),
            .I(\c0.n13443 ));
    Odrv4 I__15802 (
            .O(N__65120),
            .I(\c0.n13443 ));
    CascadeMux I__15801 (
            .O(N__65113),
            .I(N__65110));
    InMux I__15800 (
            .O(N__65110),
            .I(N__65107));
    LocalMux I__15799 (
            .O(N__65107),
            .I(N__65104));
    Span4Mux_v I__15798 (
            .O(N__65104),
            .I(N__65100));
    CascadeMux I__15797 (
            .O(N__65103),
            .I(N__65097));
    Span4Mux_h I__15796 (
            .O(N__65100),
            .I(N__65094));
    InMux I__15795 (
            .O(N__65097),
            .I(N__65091));
    Sp12to4 I__15794 (
            .O(N__65094),
            .I(N__65086));
    LocalMux I__15793 (
            .O(N__65091),
            .I(N__65086));
    Span12Mux_v I__15792 (
            .O(N__65086),
            .I(N__65083));
    Odrv12 I__15791 (
            .O(N__65083),
            .I(\c0.n22358 ));
    InMux I__15790 (
            .O(N__65080),
            .I(N__65077));
    LocalMux I__15789 (
            .O(N__65077),
            .I(N__65074));
    Span4Mux_v I__15788 (
            .O(N__65074),
            .I(N__65070));
    InMux I__15787 (
            .O(N__65073),
            .I(N__65067));
    Odrv4 I__15786 (
            .O(N__65070),
            .I(\c0.n22099 ));
    LocalMux I__15785 (
            .O(N__65067),
            .I(\c0.n22099 ));
    InMux I__15784 (
            .O(N__65062),
            .I(N__65054));
    InMux I__15783 (
            .O(N__65061),
            .I(N__65054));
    CascadeMux I__15782 (
            .O(N__65060),
            .I(N__65050));
    InMux I__15781 (
            .O(N__65059),
            .I(N__65047));
    LocalMux I__15780 (
            .O(N__65054),
            .I(N__65044));
    CascadeMux I__15779 (
            .O(N__65053),
            .I(N__65041));
    InMux I__15778 (
            .O(N__65050),
            .I(N__65038));
    LocalMux I__15777 (
            .O(N__65047),
            .I(N__65035));
    Span4Mux_h I__15776 (
            .O(N__65044),
            .I(N__65032));
    InMux I__15775 (
            .O(N__65041),
            .I(N__65029));
    LocalMux I__15774 (
            .O(N__65038),
            .I(\c0.data_in_frame_24_1 ));
    Odrv12 I__15773 (
            .O(N__65035),
            .I(\c0.data_in_frame_24_1 ));
    Odrv4 I__15772 (
            .O(N__65032),
            .I(\c0.data_in_frame_24_1 ));
    LocalMux I__15771 (
            .O(N__65029),
            .I(\c0.data_in_frame_24_1 ));
    InMux I__15770 (
            .O(N__65020),
            .I(N__65017));
    LocalMux I__15769 (
            .O(N__65017),
            .I(N__65013));
    InMux I__15768 (
            .O(N__65016),
            .I(N__65010));
    Span4Mux_h I__15767 (
            .O(N__65013),
            .I(N__65007));
    LocalMux I__15766 (
            .O(N__65010),
            .I(N__65004));
    Span4Mux_h I__15765 (
            .O(N__65007),
            .I(N__65001));
    Span12Mux_v I__15764 (
            .O(N__65004),
            .I(N__64998));
    Span4Mux_v I__15763 (
            .O(N__65001),
            .I(N__64995));
    Odrv12 I__15762 (
            .O(N__64998),
            .I(\c0.n22057 ));
    Odrv4 I__15761 (
            .O(N__64995),
            .I(\c0.n22057 ));
    InMux I__15760 (
            .O(N__64990),
            .I(N__64986));
    InMux I__15759 (
            .O(N__64989),
            .I(N__64983));
    LocalMux I__15758 (
            .O(N__64986),
            .I(N__64980));
    LocalMux I__15757 (
            .O(N__64983),
            .I(\c0.n22373 ));
    Odrv12 I__15756 (
            .O(N__64980),
            .I(\c0.n22373 ));
    CascadeMux I__15755 (
            .O(N__64975),
            .I(\c0.n8_adj_4288_cascade_ ));
    InMux I__15754 (
            .O(N__64972),
            .I(N__64969));
    LocalMux I__15753 (
            .O(N__64969),
            .I(N__64966));
    Odrv12 I__15752 (
            .O(N__64966),
            .I(\c0.n24_adj_4289 ));
    InMux I__15751 (
            .O(N__64963),
            .I(N__64957));
    InMux I__15750 (
            .O(N__64962),
            .I(N__64957));
    LocalMux I__15749 (
            .O(N__64957),
            .I(N__64954));
    Odrv4 I__15748 (
            .O(N__64954),
            .I(\c0.n22215 ));
    InMux I__15747 (
            .O(N__64951),
            .I(N__64948));
    LocalMux I__15746 (
            .O(N__64948),
            .I(N__64944));
    InMux I__15745 (
            .O(N__64947),
            .I(N__64941));
    Span4Mux_v I__15744 (
            .O(N__64944),
            .I(N__64938));
    LocalMux I__15743 (
            .O(N__64941),
            .I(\c0.n22402 ));
    Odrv4 I__15742 (
            .O(N__64938),
            .I(\c0.n22402 ));
    CascadeMux I__15741 (
            .O(N__64933),
            .I(N__64929));
    CascadeMux I__15740 (
            .O(N__64932),
            .I(N__64926));
    InMux I__15739 (
            .O(N__64929),
            .I(N__64923));
    InMux I__15738 (
            .O(N__64926),
            .I(N__64920));
    LocalMux I__15737 (
            .O(N__64923),
            .I(N__64917));
    LocalMux I__15736 (
            .O(N__64920),
            .I(\c0.data_in_frame_28_4 ));
    Odrv12 I__15735 (
            .O(N__64917),
            .I(\c0.data_in_frame_28_4 ));
    InMux I__15734 (
            .O(N__64912),
            .I(N__64908));
    InMux I__15733 (
            .O(N__64911),
            .I(N__64905));
    LocalMux I__15732 (
            .O(N__64908),
            .I(\c0.n22455 ));
    LocalMux I__15731 (
            .O(N__64905),
            .I(\c0.n22455 ));
    InMux I__15730 (
            .O(N__64900),
            .I(N__64897));
    LocalMux I__15729 (
            .O(N__64897),
            .I(\c0.n22997 ));
    InMux I__15728 (
            .O(N__64894),
            .I(N__64889));
    CascadeMux I__15727 (
            .O(N__64893),
            .I(N__64880));
    CascadeMux I__15726 (
            .O(N__64892),
            .I(N__64876));
    LocalMux I__15725 (
            .O(N__64889),
            .I(N__64868));
    InMux I__15724 (
            .O(N__64888),
            .I(N__64865));
    InMux I__15723 (
            .O(N__64887),
            .I(N__64859));
    InMux I__15722 (
            .O(N__64886),
            .I(N__64854));
    InMux I__15721 (
            .O(N__64885),
            .I(N__64854));
    InMux I__15720 (
            .O(N__64884),
            .I(N__64846));
    InMux I__15719 (
            .O(N__64883),
            .I(N__64846));
    InMux I__15718 (
            .O(N__64880),
            .I(N__64843));
    InMux I__15717 (
            .O(N__64879),
            .I(N__64840));
    InMux I__15716 (
            .O(N__64876),
            .I(N__64837));
    InMux I__15715 (
            .O(N__64875),
            .I(N__64833));
    InMux I__15714 (
            .O(N__64874),
            .I(N__64830));
    InMux I__15713 (
            .O(N__64873),
            .I(N__64827));
    InMux I__15712 (
            .O(N__64872),
            .I(N__64820));
    InMux I__15711 (
            .O(N__64871),
            .I(N__64815));
    Span4Mux_v I__15710 (
            .O(N__64868),
            .I(N__64812));
    LocalMux I__15709 (
            .O(N__64865),
            .I(N__64809));
    InMux I__15708 (
            .O(N__64864),
            .I(N__64806));
    InMux I__15707 (
            .O(N__64863),
            .I(N__64803));
    InMux I__15706 (
            .O(N__64862),
            .I(N__64800));
    LocalMux I__15705 (
            .O(N__64859),
            .I(N__64797));
    LocalMux I__15704 (
            .O(N__64854),
            .I(N__64794));
    InMux I__15703 (
            .O(N__64853),
            .I(N__64789));
    InMux I__15702 (
            .O(N__64852),
            .I(N__64789));
    InMux I__15701 (
            .O(N__64851),
            .I(N__64786));
    LocalMux I__15700 (
            .O(N__64846),
            .I(N__64781));
    LocalMux I__15699 (
            .O(N__64843),
            .I(N__64781));
    LocalMux I__15698 (
            .O(N__64840),
            .I(N__64778));
    LocalMux I__15697 (
            .O(N__64837),
            .I(N__64775));
    InMux I__15696 (
            .O(N__64836),
            .I(N__64772));
    LocalMux I__15695 (
            .O(N__64833),
            .I(N__64767));
    LocalMux I__15694 (
            .O(N__64830),
            .I(N__64767));
    LocalMux I__15693 (
            .O(N__64827),
            .I(N__64764));
    InMux I__15692 (
            .O(N__64826),
            .I(N__64761));
    InMux I__15691 (
            .O(N__64825),
            .I(N__64758));
    InMux I__15690 (
            .O(N__64824),
            .I(N__64755));
    InMux I__15689 (
            .O(N__64823),
            .I(N__64752));
    LocalMux I__15688 (
            .O(N__64820),
            .I(N__64749));
    CascadeMux I__15687 (
            .O(N__64819),
            .I(N__64745));
    InMux I__15686 (
            .O(N__64818),
            .I(N__64742));
    LocalMux I__15685 (
            .O(N__64815),
            .I(N__64739));
    Span4Mux_h I__15684 (
            .O(N__64812),
            .I(N__64734));
    Span4Mux_v I__15683 (
            .O(N__64809),
            .I(N__64734));
    LocalMux I__15682 (
            .O(N__64806),
            .I(N__64731));
    LocalMux I__15681 (
            .O(N__64803),
            .I(N__64726));
    LocalMux I__15680 (
            .O(N__64800),
            .I(N__64726));
    Span4Mux_h I__15679 (
            .O(N__64797),
            .I(N__64721));
    Span4Mux_v I__15678 (
            .O(N__64794),
            .I(N__64721));
    LocalMux I__15677 (
            .O(N__64789),
            .I(N__64718));
    LocalMux I__15676 (
            .O(N__64786),
            .I(N__64715));
    Span4Mux_h I__15675 (
            .O(N__64781),
            .I(N__64706));
    Span4Mux_v I__15674 (
            .O(N__64778),
            .I(N__64706));
    Span4Mux_h I__15673 (
            .O(N__64775),
            .I(N__64706));
    LocalMux I__15672 (
            .O(N__64772),
            .I(N__64706));
    Span4Mux_v I__15671 (
            .O(N__64767),
            .I(N__64701));
    Span4Mux_h I__15670 (
            .O(N__64764),
            .I(N__64701));
    LocalMux I__15669 (
            .O(N__64761),
            .I(N__64695));
    LocalMux I__15668 (
            .O(N__64758),
            .I(N__64692));
    LocalMux I__15667 (
            .O(N__64755),
            .I(N__64689));
    LocalMux I__15666 (
            .O(N__64752),
            .I(N__64686));
    Span4Mux_h I__15665 (
            .O(N__64749),
            .I(N__64683));
    InMux I__15664 (
            .O(N__64748),
            .I(N__64678));
    InMux I__15663 (
            .O(N__64745),
            .I(N__64678));
    LocalMux I__15662 (
            .O(N__64742),
            .I(N__64671));
    Span4Mux_v I__15661 (
            .O(N__64739),
            .I(N__64671));
    Span4Mux_v I__15660 (
            .O(N__64734),
            .I(N__64671));
    Span4Mux_v I__15659 (
            .O(N__64731),
            .I(N__64668));
    Span4Mux_v I__15658 (
            .O(N__64726),
            .I(N__64665));
    Span4Mux_v I__15657 (
            .O(N__64721),
            .I(N__64660));
    Span4Mux_h I__15656 (
            .O(N__64718),
            .I(N__64660));
    Span4Mux_h I__15655 (
            .O(N__64715),
            .I(N__64653));
    Span4Mux_v I__15654 (
            .O(N__64706),
            .I(N__64653));
    Span4Mux_h I__15653 (
            .O(N__64701),
            .I(N__64653));
    InMux I__15652 (
            .O(N__64700),
            .I(N__64650));
    InMux I__15651 (
            .O(N__64699),
            .I(N__64645));
    InMux I__15650 (
            .O(N__64698),
            .I(N__64645));
    Span4Mux_h I__15649 (
            .O(N__64695),
            .I(N__64642));
    Span4Mux_h I__15648 (
            .O(N__64692),
            .I(N__64633));
    Span4Mux_v I__15647 (
            .O(N__64689),
            .I(N__64633));
    Span4Mux_v I__15646 (
            .O(N__64686),
            .I(N__64633));
    Span4Mux_h I__15645 (
            .O(N__64683),
            .I(N__64633));
    LocalMux I__15644 (
            .O(N__64678),
            .I(N__64626));
    Sp12to4 I__15643 (
            .O(N__64671),
            .I(N__64626));
    Sp12to4 I__15642 (
            .O(N__64668),
            .I(N__64626));
    Span4Mux_h I__15641 (
            .O(N__64665),
            .I(N__64621));
    Span4Mux_h I__15640 (
            .O(N__64660),
            .I(N__64621));
    Span4Mux_v I__15639 (
            .O(N__64653),
            .I(N__64618));
    LocalMux I__15638 (
            .O(N__64650),
            .I(rx_data_3));
    LocalMux I__15637 (
            .O(N__64645),
            .I(rx_data_3));
    Odrv4 I__15636 (
            .O(N__64642),
            .I(rx_data_3));
    Odrv4 I__15635 (
            .O(N__64633),
            .I(rx_data_3));
    Odrv12 I__15634 (
            .O(N__64626),
            .I(rx_data_3));
    Odrv4 I__15633 (
            .O(N__64621),
            .I(rx_data_3));
    Odrv4 I__15632 (
            .O(N__64618),
            .I(rx_data_3));
    CascadeMux I__15631 (
            .O(N__64603),
            .I(N__64600));
    InMux I__15630 (
            .O(N__64600),
            .I(N__64596));
    InMux I__15629 (
            .O(N__64599),
            .I(N__64593));
    LocalMux I__15628 (
            .O(N__64596),
            .I(\c0.data_in_frame_28_3 ));
    LocalMux I__15627 (
            .O(N__64593),
            .I(\c0.data_in_frame_28_3 ));
    InMux I__15626 (
            .O(N__64588),
            .I(N__64584));
    CascadeMux I__15625 (
            .O(N__64587),
            .I(N__64581));
    LocalMux I__15624 (
            .O(N__64584),
            .I(N__64578));
    InMux I__15623 (
            .O(N__64581),
            .I(N__64575));
    Span4Mux_h I__15622 (
            .O(N__64578),
            .I(N__64572));
    LocalMux I__15621 (
            .O(N__64575),
            .I(\c0.data_in_frame_28_7 ));
    Odrv4 I__15620 (
            .O(N__64572),
            .I(\c0.data_in_frame_28_7 ));
    CascadeMux I__15619 (
            .O(N__64567),
            .I(N__64562));
    InMux I__15618 (
            .O(N__64566),
            .I(N__64557));
    InMux I__15617 (
            .O(N__64565),
            .I(N__64553));
    InMux I__15616 (
            .O(N__64562),
            .I(N__64546));
    InMux I__15615 (
            .O(N__64561),
            .I(N__64543));
    InMux I__15614 (
            .O(N__64560),
            .I(N__64540));
    LocalMux I__15613 (
            .O(N__64557),
            .I(N__64537));
    CascadeMux I__15612 (
            .O(N__64556),
            .I(N__64528));
    LocalMux I__15611 (
            .O(N__64553),
            .I(N__64524));
    CascadeMux I__15610 (
            .O(N__64552),
            .I(N__64520));
    CascadeMux I__15609 (
            .O(N__64551),
            .I(N__64514));
    InMux I__15608 (
            .O(N__64550),
            .I(N__64508));
    InMux I__15607 (
            .O(N__64549),
            .I(N__64505));
    LocalMux I__15606 (
            .O(N__64546),
            .I(N__64502));
    LocalMux I__15605 (
            .O(N__64543),
            .I(N__64499));
    LocalMux I__15604 (
            .O(N__64540),
            .I(N__64495));
    Span4Mux_v I__15603 (
            .O(N__64537),
            .I(N__64492));
    InMux I__15602 (
            .O(N__64536),
            .I(N__64487));
    InMux I__15601 (
            .O(N__64535),
            .I(N__64487));
    InMux I__15600 (
            .O(N__64534),
            .I(N__64482));
    InMux I__15599 (
            .O(N__64533),
            .I(N__64482));
    InMux I__15598 (
            .O(N__64532),
            .I(N__64478));
    InMux I__15597 (
            .O(N__64531),
            .I(N__64473));
    InMux I__15596 (
            .O(N__64528),
            .I(N__64473));
    InMux I__15595 (
            .O(N__64527),
            .I(N__64470));
    Span4Mux_h I__15594 (
            .O(N__64524),
            .I(N__64467));
    InMux I__15593 (
            .O(N__64523),
            .I(N__64464));
    InMux I__15592 (
            .O(N__64520),
            .I(N__64459));
    InMux I__15591 (
            .O(N__64519),
            .I(N__64459));
    InMux I__15590 (
            .O(N__64518),
            .I(N__64455));
    InMux I__15589 (
            .O(N__64517),
            .I(N__64452));
    InMux I__15588 (
            .O(N__64514),
            .I(N__64448));
    InMux I__15587 (
            .O(N__64513),
            .I(N__64441));
    InMux I__15586 (
            .O(N__64512),
            .I(N__64441));
    InMux I__15585 (
            .O(N__64511),
            .I(N__64441));
    LocalMux I__15584 (
            .O(N__64508),
            .I(N__64438));
    LocalMux I__15583 (
            .O(N__64505),
            .I(N__64435));
    Span4Mux_v I__15582 (
            .O(N__64502),
            .I(N__64430));
    Span4Mux_h I__15581 (
            .O(N__64499),
            .I(N__64430));
    InMux I__15580 (
            .O(N__64498),
            .I(N__64427));
    Span4Mux_h I__15579 (
            .O(N__64495),
            .I(N__64420));
    Span4Mux_h I__15578 (
            .O(N__64492),
            .I(N__64420));
    LocalMux I__15577 (
            .O(N__64487),
            .I(N__64420));
    LocalMux I__15576 (
            .O(N__64482),
            .I(N__64417));
    InMux I__15575 (
            .O(N__64481),
            .I(N__64414));
    LocalMux I__15574 (
            .O(N__64478),
            .I(N__64411));
    LocalMux I__15573 (
            .O(N__64473),
            .I(N__64404));
    LocalMux I__15572 (
            .O(N__64470),
            .I(N__64404));
    Span4Mux_v I__15571 (
            .O(N__64467),
            .I(N__64404));
    LocalMux I__15570 (
            .O(N__64464),
            .I(N__64399));
    LocalMux I__15569 (
            .O(N__64459),
            .I(N__64399));
    CascadeMux I__15568 (
            .O(N__64458),
            .I(N__64396));
    LocalMux I__15567 (
            .O(N__64455),
            .I(N__64391));
    LocalMux I__15566 (
            .O(N__64452),
            .I(N__64391));
    InMux I__15565 (
            .O(N__64451),
            .I(N__64388));
    LocalMux I__15564 (
            .O(N__64448),
            .I(N__64385));
    LocalMux I__15563 (
            .O(N__64441),
            .I(N__64382));
    Span4Mux_h I__15562 (
            .O(N__64438),
            .I(N__64375));
    Span4Mux_h I__15561 (
            .O(N__64435),
            .I(N__64375));
    Span4Mux_v I__15560 (
            .O(N__64430),
            .I(N__64375));
    LocalMux I__15559 (
            .O(N__64427),
            .I(N__64372));
    Span4Mux_v I__15558 (
            .O(N__64420),
            .I(N__64365));
    Span4Mux_h I__15557 (
            .O(N__64417),
            .I(N__64365));
    LocalMux I__15556 (
            .O(N__64414),
            .I(N__64365));
    Span4Mux_h I__15555 (
            .O(N__64411),
            .I(N__64358));
    Span4Mux_v I__15554 (
            .O(N__64404),
            .I(N__64358));
    Span4Mux_h I__15553 (
            .O(N__64399),
            .I(N__64358));
    InMux I__15552 (
            .O(N__64396),
            .I(N__64353));
    Span4Mux_h I__15551 (
            .O(N__64391),
            .I(N__64350));
    LocalMux I__15550 (
            .O(N__64388),
            .I(N__64347));
    Span4Mux_v I__15549 (
            .O(N__64385),
            .I(N__64342));
    Span12Mux_h I__15548 (
            .O(N__64382),
            .I(N__64339));
    Span4Mux_v I__15547 (
            .O(N__64375),
            .I(N__64336));
    Span4Mux_v I__15546 (
            .O(N__64372),
            .I(N__64333));
    Span4Mux_v I__15545 (
            .O(N__64365),
            .I(N__64328));
    Span4Mux_v I__15544 (
            .O(N__64358),
            .I(N__64328));
    InMux I__15543 (
            .O(N__64357),
            .I(N__64323));
    InMux I__15542 (
            .O(N__64356),
            .I(N__64323));
    LocalMux I__15541 (
            .O(N__64353),
            .I(N__64316));
    Span4Mux_h I__15540 (
            .O(N__64350),
            .I(N__64316));
    Span4Mux_h I__15539 (
            .O(N__64347),
            .I(N__64316));
    InMux I__15538 (
            .O(N__64346),
            .I(N__64313));
    InMux I__15537 (
            .O(N__64345),
            .I(N__64310));
    Sp12to4 I__15536 (
            .O(N__64342),
            .I(N__64305));
    Span12Mux_v I__15535 (
            .O(N__64339),
            .I(N__64305));
    Span4Mux_h I__15534 (
            .O(N__64336),
            .I(N__64302));
    Span4Mux_v I__15533 (
            .O(N__64333),
            .I(N__64299));
    Span4Mux_h I__15532 (
            .O(N__64328),
            .I(N__64296));
    LocalMux I__15531 (
            .O(N__64323),
            .I(N__64291));
    Span4Mux_v I__15530 (
            .O(N__64316),
            .I(N__64291));
    LocalMux I__15529 (
            .O(N__64313),
            .I(\c0.n9_adj_4217 ));
    LocalMux I__15528 (
            .O(N__64310),
            .I(\c0.n9_adj_4217 ));
    Odrv12 I__15527 (
            .O(N__64305),
            .I(\c0.n9_adj_4217 ));
    Odrv4 I__15526 (
            .O(N__64302),
            .I(\c0.n9_adj_4217 ));
    Odrv4 I__15525 (
            .O(N__64299),
            .I(\c0.n9_adj_4217 ));
    Odrv4 I__15524 (
            .O(N__64296),
            .I(\c0.n9_adj_4217 ));
    Odrv4 I__15523 (
            .O(N__64291),
            .I(\c0.n9_adj_4217 ));
    CascadeMux I__15522 (
            .O(N__64276),
            .I(N__64272));
    CascadeMux I__15521 (
            .O(N__64275),
            .I(N__64269));
    InMux I__15520 (
            .O(N__64272),
            .I(N__64266));
    InMux I__15519 (
            .O(N__64269),
            .I(N__64263));
    LocalMux I__15518 (
            .O(N__64266),
            .I(\c0.data_in_frame_28_6 ));
    LocalMux I__15517 (
            .O(N__64263),
            .I(\c0.data_in_frame_28_6 ));
    InMux I__15516 (
            .O(N__64258),
            .I(N__64254));
    InMux I__15515 (
            .O(N__64257),
            .I(N__64251));
    LocalMux I__15514 (
            .O(N__64254),
            .I(N__64248));
    LocalMux I__15513 (
            .O(N__64251),
            .I(N__64245));
    Span4Mux_v I__15512 (
            .O(N__64248),
            .I(N__64239));
    Span4Mux_h I__15511 (
            .O(N__64245),
            .I(N__64239));
    InMux I__15510 (
            .O(N__64244),
            .I(N__64236));
    Sp12to4 I__15509 (
            .O(N__64239),
            .I(N__64231));
    LocalMux I__15508 (
            .O(N__64236),
            .I(N__64231));
    Odrv12 I__15507 (
            .O(N__64231),
            .I(\c0.n22105 ));
    InMux I__15506 (
            .O(N__64228),
            .I(N__64225));
    LocalMux I__15505 (
            .O(N__64225),
            .I(N__64221));
    InMux I__15504 (
            .O(N__64224),
            .I(N__64216));
    Span4Mux_h I__15503 (
            .O(N__64221),
            .I(N__64213));
    InMux I__15502 (
            .O(N__64220),
            .I(N__64208));
    InMux I__15501 (
            .O(N__64219),
            .I(N__64208));
    LocalMux I__15500 (
            .O(N__64216),
            .I(N__64204));
    Span4Mux_v I__15499 (
            .O(N__64213),
            .I(N__64199));
    LocalMux I__15498 (
            .O(N__64208),
            .I(N__64199));
    InMux I__15497 (
            .O(N__64207),
            .I(N__64196));
    Odrv12 I__15496 (
            .O(N__64204),
            .I(\c0.n22849 ));
    Odrv4 I__15495 (
            .O(N__64199),
            .I(\c0.n22849 ));
    LocalMux I__15494 (
            .O(N__64196),
            .I(\c0.n22849 ));
    InMux I__15493 (
            .O(N__64189),
            .I(N__64186));
    LocalMux I__15492 (
            .O(N__64186),
            .I(N__64183));
    Span4Mux_h I__15491 (
            .O(N__64183),
            .I(N__64180));
    Odrv4 I__15490 (
            .O(N__64180),
            .I(\c0.n20406 ));
    InMux I__15489 (
            .O(N__64177),
            .I(N__64174));
    LocalMux I__15488 (
            .O(N__64174),
            .I(N__64170));
    InMux I__15487 (
            .O(N__64173),
            .I(N__64167));
    Span12Mux_s10_h I__15486 (
            .O(N__64170),
            .I(N__64164));
    LocalMux I__15485 (
            .O(N__64167),
            .I(N__64161));
    Odrv12 I__15484 (
            .O(N__64164),
            .I(\c0.n5813 ));
    Odrv4 I__15483 (
            .O(N__64161),
            .I(\c0.n5813 ));
    InMux I__15482 (
            .O(N__64156),
            .I(N__64153));
    LocalMux I__15481 (
            .O(N__64153),
            .I(N__64149));
    InMux I__15480 (
            .O(N__64152),
            .I(N__64146));
    Span4Mux_v I__15479 (
            .O(N__64149),
            .I(N__64141));
    LocalMux I__15478 (
            .O(N__64146),
            .I(N__64141));
    Span4Mux_h I__15477 (
            .O(N__64141),
            .I(N__64138));
    Odrv4 I__15476 (
            .O(N__64138),
            .I(\c0.n21864 ));
    CascadeMux I__15475 (
            .O(N__64135),
            .I(N__64132));
    InMux I__15474 (
            .O(N__64132),
            .I(N__64129));
    LocalMux I__15473 (
            .O(N__64129),
            .I(N__64126));
    Odrv4 I__15472 (
            .O(N__64126),
            .I(\c0.n13768 ));
    InMux I__15471 (
            .O(N__64123),
            .I(N__64119));
    InMux I__15470 (
            .O(N__64122),
            .I(N__64116));
    LocalMux I__15469 (
            .O(N__64119),
            .I(\c0.n22458 ));
    LocalMux I__15468 (
            .O(N__64116),
            .I(\c0.n22458 ));
    InMux I__15467 (
            .O(N__64111),
            .I(N__64106));
    InMux I__15466 (
            .O(N__64110),
            .I(N__64101));
    InMux I__15465 (
            .O(N__64109),
            .I(N__64101));
    LocalMux I__15464 (
            .O(N__64106),
            .I(N__64098));
    LocalMux I__15463 (
            .O(N__64101),
            .I(N__64095));
    Span4Mux_v I__15462 (
            .O(N__64098),
            .I(N__64092));
    Span4Mux_v I__15461 (
            .O(N__64095),
            .I(N__64089));
    Odrv4 I__15460 (
            .O(N__64092),
            .I(\c0.n21114 ));
    Odrv4 I__15459 (
            .O(N__64089),
            .I(\c0.n21114 ));
    InMux I__15458 (
            .O(N__64084),
            .I(N__64081));
    LocalMux I__15457 (
            .O(N__64081),
            .I(N__64078));
    Span4Mux_v I__15456 (
            .O(N__64078),
            .I(N__64075));
    Odrv4 I__15455 (
            .O(N__64075),
            .I(\c0.n18_adj_4246 ));
    CascadeMux I__15454 (
            .O(N__64072),
            .I(\c0.n21_cascade_ ));
    InMux I__15453 (
            .O(N__64069),
            .I(N__64066));
    LocalMux I__15452 (
            .O(N__64066),
            .I(N__64062));
    InMux I__15451 (
            .O(N__64065),
            .I(N__64059));
    Odrv4 I__15450 (
            .O(N__64062),
            .I(\c0.n22399 ));
    LocalMux I__15449 (
            .O(N__64059),
            .I(\c0.n22399 ));
    InMux I__15448 (
            .O(N__64054),
            .I(N__64051));
    LocalMux I__15447 (
            .O(N__64051),
            .I(\c0.n24 ));
    InMux I__15446 (
            .O(N__64048),
            .I(N__64045));
    LocalMux I__15445 (
            .O(N__64045),
            .I(N__64042));
    Span12Mux_s11_h I__15444 (
            .O(N__64042),
            .I(N__64039));
    Odrv12 I__15443 (
            .O(N__64039),
            .I(\c0.n20 ));
    InMux I__15442 (
            .O(N__64036),
            .I(N__64031));
    CascadeMux I__15441 (
            .O(N__64035),
            .I(N__64027));
    CascadeMux I__15440 (
            .O(N__64034),
            .I(N__64024));
    LocalMux I__15439 (
            .O(N__64031),
            .I(N__64021));
    CascadeMux I__15438 (
            .O(N__64030),
            .I(N__64018));
    InMux I__15437 (
            .O(N__64027),
            .I(N__64014));
    InMux I__15436 (
            .O(N__64024),
            .I(N__64011));
    Span4Mux_h I__15435 (
            .O(N__64021),
            .I(N__64008));
    InMux I__15434 (
            .O(N__64018),
            .I(N__64003));
    InMux I__15433 (
            .O(N__64017),
            .I(N__64003));
    LocalMux I__15432 (
            .O(N__64014),
            .I(\c0.data_in_frame_17_1 ));
    LocalMux I__15431 (
            .O(N__64011),
            .I(\c0.data_in_frame_17_1 ));
    Odrv4 I__15430 (
            .O(N__64008),
            .I(\c0.data_in_frame_17_1 ));
    LocalMux I__15429 (
            .O(N__64003),
            .I(\c0.data_in_frame_17_1 ));
    CascadeMux I__15428 (
            .O(N__63994),
            .I(N__63991));
    InMux I__15427 (
            .O(N__63991),
            .I(N__63988));
    LocalMux I__15426 (
            .O(N__63988),
            .I(N__63985));
    Span4Mux_v I__15425 (
            .O(N__63985),
            .I(N__63982));
    Odrv4 I__15424 (
            .O(N__63982),
            .I(\c0.n16 ));
    InMux I__15423 (
            .O(N__63979),
            .I(N__63976));
    LocalMux I__15422 (
            .O(N__63976),
            .I(N__63973));
    Span4Mux_v I__15421 (
            .O(N__63973),
            .I(N__63970));
    Span4Mux_h I__15420 (
            .O(N__63970),
            .I(N__63966));
    InMux I__15419 (
            .O(N__63969),
            .I(N__63963));
    Odrv4 I__15418 (
            .O(N__63966),
            .I(\c0.n21979 ));
    LocalMux I__15417 (
            .O(N__63963),
            .I(\c0.n21979 ));
    InMux I__15416 (
            .O(N__63958),
            .I(N__63953));
    CascadeMux I__15415 (
            .O(N__63957),
            .I(N__63950));
    InMux I__15414 (
            .O(N__63956),
            .I(N__63947));
    LocalMux I__15413 (
            .O(N__63953),
            .I(N__63944));
    InMux I__15412 (
            .O(N__63950),
            .I(N__63941));
    LocalMux I__15411 (
            .O(N__63947),
            .I(N__63938));
    Span4Mux_v I__15410 (
            .O(N__63944),
            .I(N__63935));
    LocalMux I__15409 (
            .O(N__63941),
            .I(N__63932));
    Span4Mux_h I__15408 (
            .O(N__63938),
            .I(N__63929));
    Odrv4 I__15407 (
            .O(N__63935),
            .I(\c0.n23287 ));
    Odrv12 I__15406 (
            .O(N__63932),
            .I(\c0.n23287 ));
    Odrv4 I__15405 (
            .O(N__63929),
            .I(\c0.n23287 ));
    CascadeMux I__15404 (
            .O(N__63922),
            .I(\c0.n23287_cascade_ ));
    InMux I__15403 (
            .O(N__63919),
            .I(N__63914));
    InMux I__15402 (
            .O(N__63918),
            .I(N__63911));
    CascadeMux I__15401 (
            .O(N__63917),
            .I(N__63908));
    LocalMux I__15400 (
            .O(N__63914),
            .I(N__63905));
    LocalMux I__15399 (
            .O(N__63911),
            .I(N__63902));
    InMux I__15398 (
            .O(N__63908),
            .I(N__63897));
    Span4Mux_v I__15397 (
            .O(N__63905),
            .I(N__63894));
    Sp12to4 I__15396 (
            .O(N__63902),
            .I(N__63891));
    InMux I__15395 (
            .O(N__63901),
            .I(N__63886));
    InMux I__15394 (
            .O(N__63900),
            .I(N__63886));
    LocalMux I__15393 (
            .O(N__63897),
            .I(\c0.data_in_frame_19_3 ));
    Odrv4 I__15392 (
            .O(N__63894),
            .I(\c0.data_in_frame_19_3 ));
    Odrv12 I__15391 (
            .O(N__63891),
            .I(\c0.data_in_frame_19_3 ));
    LocalMux I__15390 (
            .O(N__63886),
            .I(\c0.data_in_frame_19_3 ));
    InMux I__15389 (
            .O(N__63877),
            .I(N__63873));
    InMux I__15388 (
            .O(N__63876),
            .I(N__63870));
    LocalMux I__15387 (
            .O(N__63873),
            .I(\c0.n21921 ));
    LocalMux I__15386 (
            .O(N__63870),
            .I(\c0.n21921 ));
    InMux I__15385 (
            .O(N__63865),
            .I(N__63856));
    InMux I__15384 (
            .O(N__63864),
            .I(N__63846));
    InMux I__15383 (
            .O(N__63863),
            .I(N__63843));
    InMux I__15382 (
            .O(N__63862),
            .I(N__63840));
    InMux I__15381 (
            .O(N__63861),
            .I(N__63835));
    InMux I__15380 (
            .O(N__63860),
            .I(N__63835));
    InMux I__15379 (
            .O(N__63859),
            .I(N__63832));
    LocalMux I__15378 (
            .O(N__63856),
            .I(N__63827));
    InMux I__15377 (
            .O(N__63855),
            .I(N__63820));
    InMux I__15376 (
            .O(N__63854),
            .I(N__63820));
    InMux I__15375 (
            .O(N__63853),
            .I(N__63817));
    InMux I__15374 (
            .O(N__63852),
            .I(N__63810));
    InMux I__15373 (
            .O(N__63851),
            .I(N__63807));
    InMux I__15372 (
            .O(N__63850),
            .I(N__63804));
    InMux I__15371 (
            .O(N__63849),
            .I(N__63801));
    LocalMux I__15370 (
            .O(N__63846),
            .I(N__63797));
    LocalMux I__15369 (
            .O(N__63843),
            .I(N__63794));
    LocalMux I__15368 (
            .O(N__63840),
            .I(N__63790));
    LocalMux I__15367 (
            .O(N__63835),
            .I(N__63785));
    LocalMux I__15366 (
            .O(N__63832),
            .I(N__63785));
    InMux I__15365 (
            .O(N__63831),
            .I(N__63782));
    InMux I__15364 (
            .O(N__63830),
            .I(N__63776));
    Span4Mux_h I__15363 (
            .O(N__63827),
            .I(N__63773));
    InMux I__15362 (
            .O(N__63826),
            .I(N__63770));
    InMux I__15361 (
            .O(N__63825),
            .I(N__63765));
    LocalMux I__15360 (
            .O(N__63820),
            .I(N__63761));
    LocalMux I__15359 (
            .O(N__63817),
            .I(N__63758));
    InMux I__15358 (
            .O(N__63816),
            .I(N__63753));
    InMux I__15357 (
            .O(N__63815),
            .I(N__63753));
    InMux I__15356 (
            .O(N__63814),
            .I(N__63750));
    InMux I__15355 (
            .O(N__63813),
            .I(N__63747));
    LocalMux I__15354 (
            .O(N__63810),
            .I(N__63744));
    LocalMux I__15353 (
            .O(N__63807),
            .I(N__63741));
    LocalMux I__15352 (
            .O(N__63804),
            .I(N__63738));
    LocalMux I__15351 (
            .O(N__63801),
            .I(N__63735));
    InMux I__15350 (
            .O(N__63800),
            .I(N__63732));
    Span4Mux_h I__15349 (
            .O(N__63797),
            .I(N__63727));
    Span4Mux_v I__15348 (
            .O(N__63794),
            .I(N__63727));
    InMux I__15347 (
            .O(N__63793),
            .I(N__63724));
    Span4Mux_v I__15346 (
            .O(N__63790),
            .I(N__63717));
    Span4Mux_v I__15345 (
            .O(N__63785),
            .I(N__63717));
    LocalMux I__15344 (
            .O(N__63782),
            .I(N__63717));
    InMux I__15343 (
            .O(N__63781),
            .I(N__63713));
    InMux I__15342 (
            .O(N__63780),
            .I(N__63710));
    InMux I__15341 (
            .O(N__63779),
            .I(N__63707));
    LocalMux I__15340 (
            .O(N__63776),
            .I(N__63700));
    Span4Mux_h I__15339 (
            .O(N__63773),
            .I(N__63700));
    LocalMux I__15338 (
            .O(N__63770),
            .I(N__63700));
    InMux I__15337 (
            .O(N__63769),
            .I(N__63695));
    InMux I__15336 (
            .O(N__63768),
            .I(N__63695));
    LocalMux I__15335 (
            .O(N__63765),
            .I(N__63692));
    InMux I__15334 (
            .O(N__63764),
            .I(N__63689));
    Span4Mux_v I__15333 (
            .O(N__63761),
            .I(N__63686));
    Span4Mux_h I__15332 (
            .O(N__63758),
            .I(N__63679));
    LocalMux I__15331 (
            .O(N__63753),
            .I(N__63679));
    LocalMux I__15330 (
            .O(N__63750),
            .I(N__63679));
    LocalMux I__15329 (
            .O(N__63747),
            .I(N__63672));
    Span4Mux_v I__15328 (
            .O(N__63744),
            .I(N__63672));
    Span4Mux_v I__15327 (
            .O(N__63741),
            .I(N__63672));
    Span4Mux_h I__15326 (
            .O(N__63738),
            .I(N__63665));
    Span4Mux_v I__15325 (
            .O(N__63735),
            .I(N__63665));
    LocalMux I__15324 (
            .O(N__63732),
            .I(N__63665));
    Sp12to4 I__15323 (
            .O(N__63727),
            .I(N__63660));
    LocalMux I__15322 (
            .O(N__63724),
            .I(N__63660));
    Span4Mux_h I__15321 (
            .O(N__63717),
            .I(N__63657));
    InMux I__15320 (
            .O(N__63716),
            .I(N__63654));
    LocalMux I__15319 (
            .O(N__63713),
            .I(N__63651));
    LocalMux I__15318 (
            .O(N__63710),
            .I(N__63644));
    LocalMux I__15317 (
            .O(N__63707),
            .I(N__63644));
    Span4Mux_h I__15316 (
            .O(N__63700),
            .I(N__63644));
    LocalMux I__15315 (
            .O(N__63695),
            .I(N__63638));
    Span4Mux_v I__15314 (
            .O(N__63692),
            .I(N__63638));
    LocalMux I__15313 (
            .O(N__63689),
            .I(N__63633));
    Span4Mux_h I__15312 (
            .O(N__63686),
            .I(N__63633));
    Span4Mux_h I__15311 (
            .O(N__63679),
            .I(N__63626));
    Span4Mux_h I__15310 (
            .O(N__63672),
            .I(N__63626));
    Span4Mux_v I__15309 (
            .O(N__63665),
            .I(N__63626));
    Span12Mux_h I__15308 (
            .O(N__63660),
            .I(N__63623));
    Sp12to4 I__15307 (
            .O(N__63657),
            .I(N__63620));
    LocalMux I__15306 (
            .O(N__63654),
            .I(N__63617));
    Span4Mux_h I__15305 (
            .O(N__63651),
            .I(N__63612));
    Span4Mux_v I__15304 (
            .O(N__63644),
            .I(N__63612));
    InMux I__15303 (
            .O(N__63643),
            .I(N__63609));
    Span4Mux_v I__15302 (
            .O(N__63638),
            .I(N__63606));
    Span4Mux_v I__15301 (
            .O(N__63633),
            .I(N__63603));
    Span4Mux_v I__15300 (
            .O(N__63626),
            .I(N__63600));
    Span12Mux_v I__15299 (
            .O(N__63623),
            .I(N__63597));
    Span12Mux_s10_v I__15298 (
            .O(N__63620),
            .I(N__63592));
    Span12Mux_h I__15297 (
            .O(N__63617),
            .I(N__63592));
    Span4Mux_v I__15296 (
            .O(N__63612),
            .I(N__63589));
    LocalMux I__15295 (
            .O(N__63609),
            .I(rx_data_1));
    Odrv4 I__15294 (
            .O(N__63606),
            .I(rx_data_1));
    Odrv4 I__15293 (
            .O(N__63603),
            .I(rx_data_1));
    Odrv4 I__15292 (
            .O(N__63600),
            .I(rx_data_1));
    Odrv12 I__15291 (
            .O(N__63597),
            .I(rx_data_1));
    Odrv12 I__15290 (
            .O(N__63592),
            .I(rx_data_1));
    Odrv4 I__15289 (
            .O(N__63589),
            .I(rx_data_1));
    CascadeMux I__15288 (
            .O(N__63574),
            .I(N__63570));
    InMux I__15287 (
            .O(N__63573),
            .I(N__63567));
    InMux I__15286 (
            .O(N__63570),
            .I(N__63564));
    LocalMux I__15285 (
            .O(N__63567),
            .I(N__63561));
    LocalMux I__15284 (
            .O(N__63564),
            .I(N__63555));
    Span4Mux_v I__15283 (
            .O(N__63561),
            .I(N__63555));
    InMux I__15282 (
            .O(N__63560),
            .I(N__63552));
    Odrv4 I__15281 (
            .O(N__63555),
            .I(\c0.data_in_frame_24_0 ));
    LocalMux I__15280 (
            .O(N__63552),
            .I(\c0.data_in_frame_24_0 ));
    InMux I__15279 (
            .O(N__63547),
            .I(N__63543));
    CascadeMux I__15278 (
            .O(N__63546),
            .I(N__63540));
    LocalMux I__15277 (
            .O(N__63543),
            .I(N__63535));
    InMux I__15276 (
            .O(N__63540),
            .I(N__63532));
    CascadeMux I__15275 (
            .O(N__63539),
            .I(N__63529));
    InMux I__15274 (
            .O(N__63538),
            .I(N__63526));
    Span4Mux_h I__15273 (
            .O(N__63535),
            .I(N__63523));
    LocalMux I__15272 (
            .O(N__63532),
            .I(N__63520));
    InMux I__15271 (
            .O(N__63529),
            .I(N__63517));
    LocalMux I__15270 (
            .O(N__63526),
            .I(N__63510));
    Span4Mux_h I__15269 (
            .O(N__63523),
            .I(N__63510));
    Span4Mux_h I__15268 (
            .O(N__63520),
            .I(N__63510));
    LocalMux I__15267 (
            .O(N__63517),
            .I(\c0.data_in_frame_24_5 ));
    Odrv4 I__15266 (
            .O(N__63510),
            .I(\c0.data_in_frame_24_5 ));
    CascadeMux I__15265 (
            .O(N__63505),
            .I(N__63502));
    InMux I__15264 (
            .O(N__63502),
            .I(N__63498));
    InMux I__15263 (
            .O(N__63501),
            .I(N__63495));
    LocalMux I__15262 (
            .O(N__63498),
            .I(\c0.n13320 ));
    LocalMux I__15261 (
            .O(N__63495),
            .I(\c0.n13320 ));
    InMux I__15260 (
            .O(N__63490),
            .I(N__63487));
    LocalMux I__15259 (
            .O(N__63487),
            .I(N__63482));
    InMux I__15258 (
            .O(N__63486),
            .I(N__63479));
    InMux I__15257 (
            .O(N__63485),
            .I(N__63476));
    Span4Mux_h I__15256 (
            .O(N__63482),
            .I(N__63470));
    LocalMux I__15255 (
            .O(N__63479),
            .I(N__63470));
    LocalMux I__15254 (
            .O(N__63476),
            .I(N__63467));
    CascadeMux I__15253 (
            .O(N__63475),
            .I(N__63464));
    Span4Mux_v I__15252 (
            .O(N__63470),
            .I(N__63459));
    Span4Mux_v I__15251 (
            .O(N__63467),
            .I(N__63459));
    InMux I__15250 (
            .O(N__63464),
            .I(N__63456));
    Sp12to4 I__15249 (
            .O(N__63459),
            .I(N__63450));
    LocalMux I__15248 (
            .O(N__63456),
            .I(N__63450));
    InMux I__15247 (
            .O(N__63455),
            .I(N__63447));
    Span12Mux_h I__15246 (
            .O(N__63450),
            .I(N__63444));
    LocalMux I__15245 (
            .O(N__63447),
            .I(data_in_frame_22_5));
    Odrv12 I__15244 (
            .O(N__63444),
            .I(data_in_frame_22_5));
    InMux I__15243 (
            .O(N__63439),
            .I(N__63436));
    LocalMux I__15242 (
            .O(N__63436),
            .I(N__63433));
    Span4Mux_h I__15241 (
            .O(N__63433),
            .I(N__63429));
    InMux I__15240 (
            .O(N__63432),
            .I(N__63426));
    Odrv4 I__15239 (
            .O(N__63429),
            .I(\c0.n22255 ));
    LocalMux I__15238 (
            .O(N__63426),
            .I(\c0.n22255 ));
    CascadeMux I__15237 (
            .O(N__63421),
            .I(N__63418));
    InMux I__15236 (
            .O(N__63418),
            .I(N__63413));
    CascadeMux I__15235 (
            .O(N__63417),
            .I(N__63410));
    CascadeMux I__15234 (
            .O(N__63416),
            .I(N__63407));
    LocalMux I__15233 (
            .O(N__63413),
            .I(N__63404));
    InMux I__15232 (
            .O(N__63410),
            .I(N__63401));
    InMux I__15231 (
            .O(N__63407),
            .I(N__63398));
    Span4Mux_h I__15230 (
            .O(N__63404),
            .I(N__63395));
    LocalMux I__15229 (
            .O(N__63401),
            .I(\c0.data_in_frame_19_1 ));
    LocalMux I__15228 (
            .O(N__63398),
            .I(\c0.data_in_frame_19_1 ));
    Odrv4 I__15227 (
            .O(N__63395),
            .I(\c0.data_in_frame_19_1 ));
    InMux I__15226 (
            .O(N__63388),
            .I(N__63384));
    InMux I__15225 (
            .O(N__63387),
            .I(N__63381));
    LocalMux I__15224 (
            .O(N__63384),
            .I(N__63378));
    LocalMux I__15223 (
            .O(N__63381),
            .I(N__63375));
    Span4Mux_h I__15222 (
            .O(N__63378),
            .I(N__63372));
    Span4Mux_h I__15221 (
            .O(N__63375),
            .I(N__63369));
    Odrv4 I__15220 (
            .O(N__63372),
            .I(\c0.n22084 ));
    Odrv4 I__15219 (
            .O(N__63369),
            .I(\c0.n22084 ));
    InMux I__15218 (
            .O(N__63364),
            .I(N__63361));
    LocalMux I__15217 (
            .O(N__63361),
            .I(\c0.n22364 ));
    CascadeMux I__15216 (
            .O(N__63358),
            .I(N__63352));
    InMux I__15215 (
            .O(N__63357),
            .I(N__63348));
    InMux I__15214 (
            .O(N__63356),
            .I(N__63345));
    CascadeMux I__15213 (
            .O(N__63355),
            .I(N__63342));
    InMux I__15212 (
            .O(N__63352),
            .I(N__63339));
    InMux I__15211 (
            .O(N__63351),
            .I(N__63336));
    LocalMux I__15210 (
            .O(N__63348),
            .I(N__63331));
    LocalMux I__15209 (
            .O(N__63345),
            .I(N__63331));
    InMux I__15208 (
            .O(N__63342),
            .I(N__63328));
    LocalMux I__15207 (
            .O(N__63339),
            .I(N__63321));
    LocalMux I__15206 (
            .O(N__63336),
            .I(N__63321));
    Span4Mux_h I__15205 (
            .O(N__63331),
            .I(N__63321));
    LocalMux I__15204 (
            .O(N__63328),
            .I(\c0.data_in_frame_19_7 ));
    Odrv4 I__15203 (
            .O(N__63321),
            .I(\c0.data_in_frame_19_7 ));
    InMux I__15202 (
            .O(N__63316),
            .I(N__63313));
    LocalMux I__15201 (
            .O(N__63313),
            .I(\c0.n15 ));
    CascadeMux I__15200 (
            .O(N__63310),
            .I(N__63305));
    CascadeMux I__15199 (
            .O(N__63309),
            .I(N__63301));
    InMux I__15198 (
            .O(N__63308),
            .I(N__63296));
    InMux I__15197 (
            .O(N__63305),
            .I(N__63296));
    InMux I__15196 (
            .O(N__63304),
            .I(N__63292));
    InMux I__15195 (
            .O(N__63301),
            .I(N__63289));
    LocalMux I__15194 (
            .O(N__63296),
            .I(N__63286));
    InMux I__15193 (
            .O(N__63295),
            .I(N__63283));
    LocalMux I__15192 (
            .O(N__63292),
            .I(N__63280));
    LocalMux I__15191 (
            .O(N__63289),
            .I(N__63275));
    Span4Mux_v I__15190 (
            .O(N__63286),
            .I(N__63275));
    LocalMux I__15189 (
            .O(N__63283),
            .I(\c0.data_in_frame_20_5 ));
    Odrv12 I__15188 (
            .O(N__63280),
            .I(\c0.data_in_frame_20_5 ));
    Odrv4 I__15187 (
            .O(N__63275),
            .I(\c0.data_in_frame_20_5 ));
    CascadeMux I__15186 (
            .O(N__63268),
            .I(N__63264));
    InMux I__15185 (
            .O(N__63267),
            .I(N__63261));
    InMux I__15184 (
            .O(N__63264),
            .I(N__63258));
    LocalMux I__15183 (
            .O(N__63261),
            .I(N__63254));
    LocalMux I__15182 (
            .O(N__63258),
            .I(N__63251));
    InMux I__15181 (
            .O(N__63257),
            .I(N__63248));
    Span4Mux_h I__15180 (
            .O(N__63254),
            .I(N__63245));
    Odrv4 I__15179 (
            .O(N__63251),
            .I(\c0.data_in_frame_23_0 ));
    LocalMux I__15178 (
            .O(N__63248),
            .I(\c0.data_in_frame_23_0 ));
    Odrv4 I__15177 (
            .O(N__63245),
            .I(\c0.data_in_frame_23_0 ));
    InMux I__15176 (
            .O(N__63238),
            .I(N__63235));
    LocalMux I__15175 (
            .O(N__63235),
            .I(N__63232));
    Span4Mux_h I__15174 (
            .O(N__63232),
            .I(N__63229));
    Odrv4 I__15173 (
            .O(N__63229),
            .I(\c0.n26_adj_4281 ));
    InMux I__15172 (
            .O(N__63226),
            .I(N__63222));
    InMux I__15171 (
            .O(N__63225),
            .I(N__63219));
    LocalMux I__15170 (
            .O(N__63222),
            .I(N__63213));
    LocalMux I__15169 (
            .O(N__63219),
            .I(N__63210));
    InMux I__15168 (
            .O(N__63218),
            .I(N__63207));
    CascadeMux I__15167 (
            .O(N__63217),
            .I(N__63201));
    CascadeMux I__15166 (
            .O(N__63216),
            .I(N__63198));
    Span4Mux_v I__15165 (
            .O(N__63213),
            .I(N__63195));
    Span4Mux_h I__15164 (
            .O(N__63210),
            .I(N__63192));
    LocalMux I__15163 (
            .O(N__63207),
            .I(N__63189));
    InMux I__15162 (
            .O(N__63206),
            .I(N__63185));
    InMux I__15161 (
            .O(N__63205),
            .I(N__63182));
    InMux I__15160 (
            .O(N__63204),
            .I(N__63179));
    InMux I__15159 (
            .O(N__63201),
            .I(N__63165));
    InMux I__15158 (
            .O(N__63198),
            .I(N__63165));
    Span4Mux_h I__15157 (
            .O(N__63195),
            .I(N__63162));
    Span4Mux_v I__15156 (
            .O(N__63192),
            .I(N__63156));
    Span4Mux_h I__15155 (
            .O(N__63189),
            .I(N__63156));
    InMux I__15154 (
            .O(N__63188),
            .I(N__63153));
    LocalMux I__15153 (
            .O(N__63185),
            .I(N__63150));
    LocalMux I__15152 (
            .O(N__63182),
            .I(N__63147));
    LocalMux I__15151 (
            .O(N__63179),
            .I(N__63140));
    InMux I__15150 (
            .O(N__63178),
            .I(N__63136));
    InMux I__15149 (
            .O(N__63177),
            .I(N__63133));
    InMux I__15148 (
            .O(N__63176),
            .I(N__63130));
    InMux I__15147 (
            .O(N__63175),
            .I(N__63125));
    InMux I__15146 (
            .O(N__63174),
            .I(N__63125));
    InMux I__15145 (
            .O(N__63173),
            .I(N__63120));
    CascadeMux I__15144 (
            .O(N__63172),
            .I(N__63117));
    InMux I__15143 (
            .O(N__63171),
            .I(N__63114));
    InMux I__15142 (
            .O(N__63170),
            .I(N__63111));
    LocalMux I__15141 (
            .O(N__63165),
            .I(N__63108));
    Span4Mux_h I__15140 (
            .O(N__63162),
            .I(N__63103));
    InMux I__15139 (
            .O(N__63161),
            .I(N__63100));
    Span4Mux_h I__15138 (
            .O(N__63156),
            .I(N__63093));
    LocalMux I__15137 (
            .O(N__63153),
            .I(N__63093));
    Span4Mux_v I__15136 (
            .O(N__63150),
            .I(N__63093));
    Span4Mux_v I__15135 (
            .O(N__63147),
            .I(N__63089));
    InMux I__15134 (
            .O(N__63146),
            .I(N__63086));
    InMux I__15133 (
            .O(N__63145),
            .I(N__63083));
    InMux I__15132 (
            .O(N__63144),
            .I(N__63078));
    InMux I__15131 (
            .O(N__63143),
            .I(N__63078));
    Span4Mux_v I__15130 (
            .O(N__63140),
            .I(N__63075));
    InMux I__15129 (
            .O(N__63139),
            .I(N__63072));
    LocalMux I__15128 (
            .O(N__63136),
            .I(N__63069));
    LocalMux I__15127 (
            .O(N__63133),
            .I(N__63062));
    LocalMux I__15126 (
            .O(N__63130),
            .I(N__63062));
    LocalMux I__15125 (
            .O(N__63125),
            .I(N__63062));
    InMux I__15124 (
            .O(N__63124),
            .I(N__63059));
    InMux I__15123 (
            .O(N__63123),
            .I(N__63055));
    LocalMux I__15122 (
            .O(N__63120),
            .I(N__63052));
    InMux I__15121 (
            .O(N__63117),
            .I(N__63049));
    LocalMux I__15120 (
            .O(N__63114),
            .I(N__63046));
    LocalMux I__15119 (
            .O(N__63111),
            .I(N__63041));
    Span4Mux_v I__15118 (
            .O(N__63108),
            .I(N__63041));
    InMux I__15117 (
            .O(N__63107),
            .I(N__63038));
    InMux I__15116 (
            .O(N__63106),
            .I(N__63035));
    Span4Mux_v I__15115 (
            .O(N__63103),
            .I(N__63030));
    LocalMux I__15114 (
            .O(N__63100),
            .I(N__63030));
    Span4Mux_v I__15113 (
            .O(N__63093),
            .I(N__63027));
    InMux I__15112 (
            .O(N__63092),
            .I(N__63024));
    Span4Mux_v I__15111 (
            .O(N__63089),
            .I(N__63021));
    LocalMux I__15110 (
            .O(N__63086),
            .I(N__63018));
    LocalMux I__15109 (
            .O(N__63083),
            .I(N__63015));
    LocalMux I__15108 (
            .O(N__63078),
            .I(N__63010));
    Span4Mux_v I__15107 (
            .O(N__63075),
            .I(N__63010));
    LocalMux I__15106 (
            .O(N__63072),
            .I(N__63001));
    Span4Mux_v I__15105 (
            .O(N__63069),
            .I(N__63001));
    Span4Mux_v I__15104 (
            .O(N__63062),
            .I(N__63001));
    LocalMux I__15103 (
            .O(N__63059),
            .I(N__63001));
    InMux I__15102 (
            .O(N__63058),
            .I(N__62997));
    LocalMux I__15101 (
            .O(N__63055),
            .I(N__62990));
    Span4Mux_h I__15100 (
            .O(N__63052),
            .I(N__62990));
    LocalMux I__15099 (
            .O(N__63049),
            .I(N__62990));
    Span4Mux_h I__15098 (
            .O(N__63046),
            .I(N__62985));
    Span4Mux_h I__15097 (
            .O(N__63041),
            .I(N__62985));
    LocalMux I__15096 (
            .O(N__63038),
            .I(N__62982));
    LocalMux I__15095 (
            .O(N__63035),
            .I(N__62979));
    Span4Mux_v I__15094 (
            .O(N__63030),
            .I(N__62976));
    Sp12to4 I__15093 (
            .O(N__63027),
            .I(N__62972));
    LocalMux I__15092 (
            .O(N__63024),
            .I(N__62967));
    Span4Mux_v I__15091 (
            .O(N__63021),
            .I(N__62967));
    Span4Mux_v I__15090 (
            .O(N__63018),
            .I(N__62964));
    Span4Mux_v I__15089 (
            .O(N__63015),
            .I(N__62961));
    Span4Mux_h I__15088 (
            .O(N__63010),
            .I(N__62956));
    Span4Mux_v I__15087 (
            .O(N__63001),
            .I(N__62956));
    InMux I__15086 (
            .O(N__63000),
            .I(N__62953));
    LocalMux I__15085 (
            .O(N__62997),
            .I(N__62944));
    Span4Mux_h I__15084 (
            .O(N__62990),
            .I(N__62944));
    Span4Mux_v I__15083 (
            .O(N__62985),
            .I(N__62944));
    Span4Mux_v I__15082 (
            .O(N__62982),
            .I(N__62944));
    Span4Mux_v I__15081 (
            .O(N__62979),
            .I(N__62941));
    Span4Mux_v I__15080 (
            .O(N__62976),
            .I(N__62938));
    InMux I__15079 (
            .O(N__62975),
            .I(N__62935));
    Span12Mux_h I__15078 (
            .O(N__62972),
            .I(N__62932));
    Sp12to4 I__15077 (
            .O(N__62967),
            .I(N__62929));
    Span4Mux_v I__15076 (
            .O(N__62964),
            .I(N__62922));
    Span4Mux_h I__15075 (
            .O(N__62961),
            .I(N__62922));
    Span4Mux_v I__15074 (
            .O(N__62956),
            .I(N__62922));
    LocalMux I__15073 (
            .O(N__62953),
            .I(N__62913));
    Span4Mux_v I__15072 (
            .O(N__62944),
            .I(N__62913));
    Span4Mux_v I__15071 (
            .O(N__62941),
            .I(N__62913));
    Span4Mux_v I__15070 (
            .O(N__62938),
            .I(N__62913));
    LocalMux I__15069 (
            .O(N__62935),
            .I(rx_data_4));
    Odrv12 I__15068 (
            .O(N__62932),
            .I(rx_data_4));
    Odrv12 I__15067 (
            .O(N__62929),
            .I(rx_data_4));
    Odrv4 I__15066 (
            .O(N__62922),
            .I(rx_data_4));
    Odrv4 I__15065 (
            .O(N__62913),
            .I(rx_data_4));
    InMux I__15064 (
            .O(N__62902),
            .I(N__62897));
    CascadeMux I__15063 (
            .O(N__62901),
            .I(N__62894));
    InMux I__15062 (
            .O(N__62900),
            .I(N__62890));
    LocalMux I__15061 (
            .O(N__62897),
            .I(N__62887));
    InMux I__15060 (
            .O(N__62894),
            .I(N__62884));
    InMux I__15059 (
            .O(N__62893),
            .I(N__62881));
    LocalMux I__15058 (
            .O(N__62890),
            .I(N__62874));
    Span4Mux_v I__15057 (
            .O(N__62887),
            .I(N__62874));
    LocalMux I__15056 (
            .O(N__62884),
            .I(N__62874));
    LocalMux I__15055 (
            .O(N__62881),
            .I(\c0.data_in_frame_18_3 ));
    Odrv4 I__15054 (
            .O(N__62874),
            .I(\c0.data_in_frame_18_3 ));
    InMux I__15053 (
            .O(N__62869),
            .I(N__62866));
    LocalMux I__15052 (
            .O(N__62866),
            .I(\c0.n22095 ));
    InMux I__15051 (
            .O(N__62863),
            .I(N__62860));
    LocalMux I__15050 (
            .O(N__62860),
            .I(\c0.n21124 ));
    CascadeMux I__15049 (
            .O(N__62857),
            .I(\c0.n22095_cascade_ ));
    InMux I__15048 (
            .O(N__62854),
            .I(N__62851));
    LocalMux I__15047 (
            .O(N__62851),
            .I(N__62847));
    InMux I__15046 (
            .O(N__62850),
            .I(N__62844));
    Odrv4 I__15045 (
            .O(N__62847),
            .I(\c0.n14143 ));
    LocalMux I__15044 (
            .O(N__62844),
            .I(\c0.n14143 ));
    InMux I__15043 (
            .O(N__62839),
            .I(N__62836));
    LocalMux I__15042 (
            .O(N__62836),
            .I(N__62833));
    Span4Mux_h I__15041 (
            .O(N__62833),
            .I(N__62830));
    Odrv4 I__15040 (
            .O(N__62830),
            .I(\c0.n29 ));
    CascadeMux I__15039 (
            .O(N__62827),
            .I(N__62823));
    InMux I__15038 (
            .O(N__62826),
            .I(N__62819));
    InMux I__15037 (
            .O(N__62823),
            .I(N__62816));
    CascadeMux I__15036 (
            .O(N__62822),
            .I(N__62812));
    LocalMux I__15035 (
            .O(N__62819),
            .I(N__62807));
    LocalMux I__15034 (
            .O(N__62816),
            .I(N__62807));
    InMux I__15033 (
            .O(N__62815),
            .I(N__62804));
    InMux I__15032 (
            .O(N__62812),
            .I(N__62801));
    Span12Mux_v I__15031 (
            .O(N__62807),
            .I(N__62798));
    LocalMux I__15030 (
            .O(N__62804),
            .I(data_in_frame_22_0));
    LocalMux I__15029 (
            .O(N__62801),
            .I(data_in_frame_22_0));
    Odrv12 I__15028 (
            .O(N__62798),
            .I(data_in_frame_22_0));
    InMux I__15027 (
            .O(N__62791),
            .I(N__62788));
    LocalMux I__15026 (
            .O(N__62788),
            .I(N__62784));
    InMux I__15025 (
            .O(N__62787),
            .I(N__62781));
    Span4Mux_v I__15024 (
            .O(N__62784),
            .I(N__62778));
    LocalMux I__15023 (
            .O(N__62781),
            .I(N__62775));
    Odrv4 I__15022 (
            .O(N__62778),
            .I(\c0.n22267 ));
    Odrv4 I__15021 (
            .O(N__62775),
            .I(\c0.n22267 ));
    InMux I__15020 (
            .O(N__62770),
            .I(N__62767));
    LocalMux I__15019 (
            .O(N__62767),
            .I(N__62762));
    InMux I__15018 (
            .O(N__62766),
            .I(N__62757));
    InMux I__15017 (
            .O(N__62765),
            .I(N__62757));
    Odrv4 I__15016 (
            .O(N__62762),
            .I(\c0.data_in_frame_20_4 ));
    LocalMux I__15015 (
            .O(N__62757),
            .I(\c0.data_in_frame_20_4 ));
    CascadeMux I__15014 (
            .O(N__62752),
            .I(N__62748));
    CascadeMux I__15013 (
            .O(N__62751),
            .I(N__62745));
    InMux I__15012 (
            .O(N__62748),
            .I(N__62742));
    InMux I__15011 (
            .O(N__62745),
            .I(N__62739));
    LocalMux I__15010 (
            .O(N__62742),
            .I(N__62736));
    LocalMux I__15009 (
            .O(N__62739),
            .I(N__62733));
    Span4Mux_v I__15008 (
            .O(N__62736),
            .I(N__62730));
    Span4Mux_v I__15007 (
            .O(N__62733),
            .I(N__62726));
    Span4Mux_h I__15006 (
            .O(N__62730),
            .I(N__62723));
    InMux I__15005 (
            .O(N__62729),
            .I(N__62720));
    Span4Mux_h I__15004 (
            .O(N__62726),
            .I(N__62717));
    Span4Mux_v I__15003 (
            .O(N__62723),
            .I(N__62714));
    LocalMux I__15002 (
            .O(N__62720),
            .I(data_in_frame_22_6));
    Odrv4 I__15001 (
            .O(N__62717),
            .I(data_in_frame_22_6));
    Odrv4 I__15000 (
            .O(N__62714),
            .I(data_in_frame_22_6));
    InMux I__14999 (
            .O(N__62707),
            .I(N__62703));
    CascadeMux I__14998 (
            .O(N__62706),
            .I(N__62699));
    LocalMux I__14997 (
            .O(N__62703),
            .I(N__62695));
    InMux I__14996 (
            .O(N__62702),
            .I(N__62690));
    InMux I__14995 (
            .O(N__62699),
            .I(N__62690));
    InMux I__14994 (
            .O(N__62698),
            .I(N__62687));
    Span4Mux_v I__14993 (
            .O(N__62695),
            .I(N__62682));
    LocalMux I__14992 (
            .O(N__62690),
            .I(N__62682));
    LocalMux I__14991 (
            .O(N__62687),
            .I(\c0.n20246 ));
    Odrv4 I__14990 (
            .O(N__62682),
            .I(\c0.n20246 ));
    InMux I__14989 (
            .O(N__62677),
            .I(N__62673));
    CascadeMux I__14988 (
            .O(N__62676),
            .I(N__62668));
    LocalMux I__14987 (
            .O(N__62673),
            .I(N__62665));
    InMux I__14986 (
            .O(N__62672),
            .I(N__62662));
    InMux I__14985 (
            .O(N__62671),
            .I(N__62658));
    InMux I__14984 (
            .O(N__62668),
            .I(N__62655));
    Span4Mux_v I__14983 (
            .O(N__62665),
            .I(N__62650));
    LocalMux I__14982 (
            .O(N__62662),
            .I(N__62650));
    InMux I__14981 (
            .O(N__62661),
            .I(N__62647));
    LocalMux I__14980 (
            .O(N__62658),
            .I(N__62644));
    LocalMux I__14979 (
            .O(N__62655),
            .I(\c0.data_in_frame_13_6 ));
    Odrv4 I__14978 (
            .O(N__62650),
            .I(\c0.data_in_frame_13_6 ));
    LocalMux I__14977 (
            .O(N__62647),
            .I(\c0.data_in_frame_13_6 ));
    Odrv12 I__14976 (
            .O(N__62644),
            .I(\c0.data_in_frame_13_6 ));
    InMux I__14975 (
            .O(N__62635),
            .I(N__62632));
    LocalMux I__14974 (
            .O(N__62632),
            .I(N__62627));
    InMux I__14973 (
            .O(N__62631),
            .I(N__62624));
    CascadeMux I__14972 (
            .O(N__62630),
            .I(N__62621));
    Span4Mux_h I__14971 (
            .O(N__62627),
            .I(N__62618));
    LocalMux I__14970 (
            .O(N__62624),
            .I(N__62615));
    InMux I__14969 (
            .O(N__62621),
            .I(N__62612));
    Span4Mux_v I__14968 (
            .O(N__62618),
            .I(N__62609));
    Span4Mux_v I__14967 (
            .O(N__62615),
            .I(N__62606));
    LocalMux I__14966 (
            .O(N__62612),
            .I(\c0.data_in_frame_26_5 ));
    Odrv4 I__14965 (
            .O(N__62609),
            .I(\c0.data_in_frame_26_5 ));
    Odrv4 I__14964 (
            .O(N__62606),
            .I(\c0.data_in_frame_26_5 ));
    InMux I__14963 (
            .O(N__62599),
            .I(N__62595));
    CascadeMux I__14962 (
            .O(N__62598),
            .I(N__62592));
    LocalMux I__14961 (
            .O(N__62595),
            .I(N__62587));
    InMux I__14960 (
            .O(N__62592),
            .I(N__62584));
    CascadeMux I__14959 (
            .O(N__62591),
            .I(N__62581));
    InMux I__14958 (
            .O(N__62590),
            .I(N__62578));
    Span4Mux_v I__14957 (
            .O(N__62587),
            .I(N__62573));
    LocalMux I__14956 (
            .O(N__62584),
            .I(N__62573));
    InMux I__14955 (
            .O(N__62581),
            .I(N__62570));
    LocalMux I__14954 (
            .O(N__62578),
            .I(N__62567));
    Span4Mux_h I__14953 (
            .O(N__62573),
            .I(N__62564));
    LocalMux I__14952 (
            .O(N__62570),
            .I(\c0.data_in_frame_21_6 ));
    Odrv12 I__14951 (
            .O(N__62567),
            .I(\c0.data_in_frame_21_6 ));
    Odrv4 I__14950 (
            .O(N__62564),
            .I(\c0.data_in_frame_21_6 ));
    InMux I__14949 (
            .O(N__62557),
            .I(N__62551));
    InMux I__14948 (
            .O(N__62556),
            .I(N__62546));
    InMux I__14947 (
            .O(N__62555),
            .I(N__62546));
    InMux I__14946 (
            .O(N__62554),
            .I(N__62535));
    LocalMux I__14945 (
            .O(N__62551),
            .I(N__62532));
    LocalMux I__14944 (
            .O(N__62546),
            .I(N__62519));
    InMux I__14943 (
            .O(N__62545),
            .I(N__62514));
    InMux I__14942 (
            .O(N__62544),
            .I(N__62514));
    InMux I__14941 (
            .O(N__62543),
            .I(N__62511));
    InMux I__14940 (
            .O(N__62542),
            .I(N__62487));
    InMux I__14939 (
            .O(N__62541),
            .I(N__62484));
    InMux I__14938 (
            .O(N__62540),
            .I(N__62477));
    InMux I__14937 (
            .O(N__62539),
            .I(N__62477));
    InMux I__14936 (
            .O(N__62538),
            .I(N__62477));
    LocalMux I__14935 (
            .O(N__62535),
            .I(N__62472));
    Span4Mux_v I__14934 (
            .O(N__62532),
            .I(N__62472));
    InMux I__14933 (
            .O(N__62531),
            .I(N__62465));
    InMux I__14932 (
            .O(N__62530),
            .I(N__62465));
    InMux I__14931 (
            .O(N__62529),
            .I(N__62465));
    InMux I__14930 (
            .O(N__62528),
            .I(N__62458));
    InMux I__14929 (
            .O(N__62527),
            .I(N__62458));
    InMux I__14928 (
            .O(N__62526),
            .I(N__62458));
    InMux I__14927 (
            .O(N__62525),
            .I(N__62449));
    InMux I__14926 (
            .O(N__62524),
            .I(N__62449));
    InMux I__14925 (
            .O(N__62523),
            .I(N__62449));
    InMux I__14924 (
            .O(N__62522),
            .I(N__62449));
    Span4Mux_v I__14923 (
            .O(N__62519),
            .I(N__62444));
    LocalMux I__14922 (
            .O(N__62514),
            .I(N__62444));
    LocalMux I__14921 (
            .O(N__62511),
            .I(N__62441));
    InMux I__14920 (
            .O(N__62510),
            .I(N__62436));
    InMux I__14919 (
            .O(N__62509),
            .I(N__62436));
    InMux I__14918 (
            .O(N__62508),
            .I(N__62433));
    InMux I__14917 (
            .O(N__62507),
            .I(N__62422));
    InMux I__14916 (
            .O(N__62506),
            .I(N__62422));
    InMux I__14915 (
            .O(N__62505),
            .I(N__62417));
    InMux I__14914 (
            .O(N__62504),
            .I(N__62417));
    InMux I__14913 (
            .O(N__62503),
            .I(N__62412));
    InMux I__14912 (
            .O(N__62502),
            .I(N__62412));
    InMux I__14911 (
            .O(N__62501),
            .I(N__62409));
    InMux I__14910 (
            .O(N__62500),
            .I(N__62406));
    InMux I__14909 (
            .O(N__62499),
            .I(N__62397));
    InMux I__14908 (
            .O(N__62498),
            .I(N__62397));
    InMux I__14907 (
            .O(N__62497),
            .I(N__62397));
    InMux I__14906 (
            .O(N__62496),
            .I(N__62397));
    InMux I__14905 (
            .O(N__62495),
            .I(N__62383));
    InMux I__14904 (
            .O(N__62494),
            .I(N__62383));
    InMux I__14903 (
            .O(N__62493),
            .I(N__62383));
    InMux I__14902 (
            .O(N__62492),
            .I(N__62383));
    InMux I__14901 (
            .O(N__62491),
            .I(N__62383));
    InMux I__14900 (
            .O(N__62490),
            .I(N__62383));
    LocalMux I__14899 (
            .O(N__62487),
            .I(N__62380));
    LocalMux I__14898 (
            .O(N__62484),
            .I(N__62365));
    LocalMux I__14897 (
            .O(N__62477),
            .I(N__62365));
    Span4Mux_h I__14896 (
            .O(N__62472),
            .I(N__62365));
    LocalMux I__14895 (
            .O(N__62465),
            .I(N__62365));
    LocalMux I__14894 (
            .O(N__62458),
            .I(N__62360));
    LocalMux I__14893 (
            .O(N__62449),
            .I(N__62360));
    Span4Mux_v I__14892 (
            .O(N__62444),
            .I(N__62357));
    Span4Mux_v I__14891 (
            .O(N__62441),
            .I(N__62352));
    LocalMux I__14890 (
            .O(N__62436),
            .I(N__62352));
    LocalMux I__14889 (
            .O(N__62433),
            .I(N__62348));
    InMux I__14888 (
            .O(N__62432),
            .I(N__62343));
    InMux I__14887 (
            .O(N__62431),
            .I(N__62343));
    InMux I__14886 (
            .O(N__62430),
            .I(N__62340));
    InMux I__14885 (
            .O(N__62429),
            .I(N__62333));
    InMux I__14884 (
            .O(N__62428),
            .I(N__62333));
    InMux I__14883 (
            .O(N__62427),
            .I(N__62333));
    LocalMux I__14882 (
            .O(N__62422),
            .I(N__62330));
    LocalMux I__14881 (
            .O(N__62417),
            .I(N__62327));
    LocalMux I__14880 (
            .O(N__62412),
            .I(N__62324));
    LocalMux I__14879 (
            .O(N__62409),
            .I(N__62317));
    LocalMux I__14878 (
            .O(N__62406),
            .I(N__62317));
    LocalMux I__14877 (
            .O(N__62397),
            .I(N__62317));
    InMux I__14876 (
            .O(N__62396),
            .I(N__62314));
    LocalMux I__14875 (
            .O(N__62383),
            .I(N__62311));
    Span4Mux_v I__14874 (
            .O(N__62380),
            .I(N__62308));
    InMux I__14873 (
            .O(N__62379),
            .I(N__62305));
    InMux I__14872 (
            .O(N__62378),
            .I(N__62302));
    InMux I__14871 (
            .O(N__62377),
            .I(N__62299));
    InMux I__14870 (
            .O(N__62376),
            .I(N__62292));
    InMux I__14869 (
            .O(N__62375),
            .I(N__62292));
    InMux I__14868 (
            .O(N__62374),
            .I(N__62292));
    Span4Mux_v I__14867 (
            .O(N__62365),
            .I(N__62289));
    Span4Mux_v I__14866 (
            .O(N__62360),
            .I(N__62282));
    Span4Mux_h I__14865 (
            .O(N__62357),
            .I(N__62282));
    Span4Mux_v I__14864 (
            .O(N__62352),
            .I(N__62282));
    InMux I__14863 (
            .O(N__62351),
            .I(N__62279));
    Span4Mux_v I__14862 (
            .O(N__62348),
            .I(N__62276));
    LocalMux I__14861 (
            .O(N__62343),
            .I(N__62273));
    LocalMux I__14860 (
            .O(N__62340),
            .I(N__62260));
    LocalMux I__14859 (
            .O(N__62333),
            .I(N__62260));
    Span4Mux_h I__14858 (
            .O(N__62330),
            .I(N__62260));
    Span4Mux_v I__14857 (
            .O(N__62327),
            .I(N__62260));
    Span4Mux_h I__14856 (
            .O(N__62324),
            .I(N__62260));
    Span4Mux_v I__14855 (
            .O(N__62317),
            .I(N__62260));
    LocalMux I__14854 (
            .O(N__62314),
            .I(N__62257));
    Span4Mux_v I__14853 (
            .O(N__62311),
            .I(N__62252));
    Span4Mux_h I__14852 (
            .O(N__62308),
            .I(N__62252));
    LocalMux I__14851 (
            .O(N__62305),
            .I(N__62249));
    LocalMux I__14850 (
            .O(N__62302),
            .I(N__62236));
    LocalMux I__14849 (
            .O(N__62299),
            .I(N__62236));
    LocalMux I__14848 (
            .O(N__62292),
            .I(N__62236));
    Sp12to4 I__14847 (
            .O(N__62289),
            .I(N__62236));
    Sp12to4 I__14846 (
            .O(N__62282),
            .I(N__62236));
    LocalMux I__14845 (
            .O(N__62279),
            .I(N__62236));
    Span4Mux_h I__14844 (
            .O(N__62276),
            .I(N__62233));
    Span12Mux_v I__14843 (
            .O(N__62273),
            .I(N__62230));
    Span4Mux_h I__14842 (
            .O(N__62260),
            .I(N__62227));
    Span4Mux_v I__14841 (
            .O(N__62257),
            .I(N__62222));
    Span4Mux_v I__14840 (
            .O(N__62252),
            .I(N__62222));
    Sp12to4 I__14839 (
            .O(N__62249),
            .I(N__62217));
    Span12Mux_h I__14838 (
            .O(N__62236),
            .I(N__62217));
    Odrv4 I__14837 (
            .O(N__62233),
            .I(\c0.n21749 ));
    Odrv12 I__14836 (
            .O(N__62230),
            .I(\c0.n21749 ));
    Odrv4 I__14835 (
            .O(N__62227),
            .I(\c0.n21749 ));
    Odrv4 I__14834 (
            .O(N__62222),
            .I(\c0.n21749 ));
    Odrv12 I__14833 (
            .O(N__62217),
            .I(\c0.n21749 ));
    CascadeMux I__14832 (
            .O(N__62206),
            .I(N__62199));
    CascadeMux I__14831 (
            .O(N__62205),
            .I(N__62194));
    CascadeMux I__14830 (
            .O(N__62204),
            .I(N__62191));
    CascadeMux I__14829 (
            .O(N__62203),
            .I(N__62178));
    CascadeMux I__14828 (
            .O(N__62202),
            .I(N__62174));
    InMux I__14827 (
            .O(N__62199),
            .I(N__62171));
    InMux I__14826 (
            .O(N__62198),
            .I(N__62168));
    InMux I__14825 (
            .O(N__62197),
            .I(N__62161));
    InMux I__14824 (
            .O(N__62194),
            .I(N__62161));
    InMux I__14823 (
            .O(N__62191),
            .I(N__62157));
    CascadeMux I__14822 (
            .O(N__62190),
            .I(N__62154));
    InMux I__14821 (
            .O(N__62189),
            .I(N__62151));
    InMux I__14820 (
            .O(N__62188),
            .I(N__62145));
    InMux I__14819 (
            .O(N__62187),
            .I(N__62142));
    InMux I__14818 (
            .O(N__62186),
            .I(N__62137));
    InMux I__14817 (
            .O(N__62185),
            .I(N__62137));
    InMux I__14816 (
            .O(N__62184),
            .I(N__62132));
    InMux I__14815 (
            .O(N__62183),
            .I(N__62132));
    InMux I__14814 (
            .O(N__62182),
            .I(N__62125));
    InMux I__14813 (
            .O(N__62181),
            .I(N__62125));
    InMux I__14812 (
            .O(N__62178),
            .I(N__62125));
    CascadeMux I__14811 (
            .O(N__62177),
            .I(N__62122));
    InMux I__14810 (
            .O(N__62174),
            .I(N__62117));
    LocalMux I__14809 (
            .O(N__62171),
            .I(N__62112));
    LocalMux I__14808 (
            .O(N__62168),
            .I(N__62112));
    InMux I__14807 (
            .O(N__62167),
            .I(N__62107));
    InMux I__14806 (
            .O(N__62166),
            .I(N__62107));
    LocalMux I__14805 (
            .O(N__62161),
            .I(N__62104));
    InMux I__14804 (
            .O(N__62160),
            .I(N__62101));
    LocalMux I__14803 (
            .O(N__62157),
            .I(N__62098));
    InMux I__14802 (
            .O(N__62154),
            .I(N__62095));
    LocalMux I__14801 (
            .O(N__62151),
            .I(N__62092));
    InMux I__14800 (
            .O(N__62150),
            .I(N__62089));
    CascadeMux I__14799 (
            .O(N__62149),
            .I(N__62083));
    InMux I__14798 (
            .O(N__62148),
            .I(N__62080));
    LocalMux I__14797 (
            .O(N__62145),
            .I(N__62077));
    LocalMux I__14796 (
            .O(N__62142),
            .I(N__62074));
    LocalMux I__14795 (
            .O(N__62137),
            .I(N__62071));
    LocalMux I__14794 (
            .O(N__62132),
            .I(N__62068));
    LocalMux I__14793 (
            .O(N__62125),
            .I(N__62065));
    InMux I__14792 (
            .O(N__62122),
            .I(N__62062));
    CascadeMux I__14791 (
            .O(N__62121),
            .I(N__62059));
    InMux I__14790 (
            .O(N__62120),
            .I(N__62055));
    LocalMux I__14789 (
            .O(N__62117),
            .I(N__62052));
    Span4Mux_v I__14788 (
            .O(N__62112),
            .I(N__62049));
    LocalMux I__14787 (
            .O(N__62107),
            .I(N__62046));
    Span4Mux_h I__14786 (
            .O(N__62104),
            .I(N__62043));
    LocalMux I__14785 (
            .O(N__62101),
            .I(N__62038));
    Span4Mux_h I__14784 (
            .O(N__62098),
            .I(N__62038));
    LocalMux I__14783 (
            .O(N__62095),
            .I(N__62033));
    Span4Mux_h I__14782 (
            .O(N__62092),
            .I(N__62033));
    LocalMux I__14781 (
            .O(N__62089),
            .I(N__62030));
    InMux I__14780 (
            .O(N__62088),
            .I(N__62027));
    InMux I__14779 (
            .O(N__62087),
            .I(N__62024));
    InMux I__14778 (
            .O(N__62086),
            .I(N__62021));
    InMux I__14777 (
            .O(N__62083),
            .I(N__62018));
    LocalMux I__14776 (
            .O(N__62080),
            .I(N__62015));
    Span4Mux_v I__14775 (
            .O(N__62077),
            .I(N__62010));
    Span4Mux_h I__14774 (
            .O(N__62074),
            .I(N__62010));
    Span4Mux_h I__14773 (
            .O(N__62071),
            .I(N__62007));
    Span4Mux_h I__14772 (
            .O(N__62068),
            .I(N__62004));
    Span4Mux_h I__14771 (
            .O(N__62065),
            .I(N__62001));
    LocalMux I__14770 (
            .O(N__62062),
            .I(N__61998));
    InMux I__14769 (
            .O(N__62059),
            .I(N__61995));
    InMux I__14768 (
            .O(N__62058),
            .I(N__61992));
    LocalMux I__14767 (
            .O(N__62055),
            .I(N__61989));
    Span4Mux_h I__14766 (
            .O(N__62052),
            .I(N__61982));
    Span4Mux_h I__14765 (
            .O(N__62049),
            .I(N__61982));
    Span4Mux_h I__14764 (
            .O(N__62046),
            .I(N__61982));
    Span4Mux_h I__14763 (
            .O(N__62043),
            .I(N__61977));
    Span4Mux_h I__14762 (
            .O(N__62038),
            .I(N__61977));
    Span4Mux_v I__14761 (
            .O(N__62033),
            .I(N__61974));
    Span4Mux_h I__14760 (
            .O(N__62030),
            .I(N__61971));
    LocalMux I__14759 (
            .O(N__62027),
            .I(N__61966));
    LocalMux I__14758 (
            .O(N__62024),
            .I(N__61961));
    LocalMux I__14757 (
            .O(N__62021),
            .I(N__61961));
    LocalMux I__14756 (
            .O(N__62018),
            .I(N__61950));
    Span4Mux_h I__14755 (
            .O(N__62015),
            .I(N__61950));
    Span4Mux_h I__14754 (
            .O(N__62010),
            .I(N__61950));
    Span4Mux_h I__14753 (
            .O(N__62007),
            .I(N__61950));
    Span4Mux_v I__14752 (
            .O(N__62004),
            .I(N__61950));
    Span4Mux_v I__14751 (
            .O(N__62001),
            .I(N__61945));
    Span4Mux_h I__14750 (
            .O(N__61998),
            .I(N__61945));
    LocalMux I__14749 (
            .O(N__61995),
            .I(N__61934));
    LocalMux I__14748 (
            .O(N__61992),
            .I(N__61934));
    Span12Mux_s9_h I__14747 (
            .O(N__61989),
            .I(N__61934));
    Sp12to4 I__14746 (
            .O(N__61982),
            .I(N__61934));
    Sp12to4 I__14745 (
            .O(N__61977),
            .I(N__61934));
    Span4Mux_v I__14744 (
            .O(N__61974),
            .I(N__61929));
    Span4Mux_v I__14743 (
            .O(N__61971),
            .I(N__61929));
    InMux I__14742 (
            .O(N__61970),
            .I(N__61924));
    InMux I__14741 (
            .O(N__61969),
            .I(N__61924));
    Span4Mux_h I__14740 (
            .O(N__61966),
            .I(N__61921));
    Span4Mux_v I__14739 (
            .O(N__61961),
            .I(N__61918));
    Span4Mux_v I__14738 (
            .O(N__61950),
            .I(N__61915));
    Sp12to4 I__14737 (
            .O(N__61945),
            .I(N__61910));
    Span12Mux_v I__14736 (
            .O(N__61934),
            .I(N__61910));
    Span4Mux_h I__14735 (
            .O(N__61929),
            .I(N__61907));
    LocalMux I__14734 (
            .O(N__61924),
            .I(\c0.n9_adj_4237 ));
    Odrv4 I__14733 (
            .O(N__61921),
            .I(\c0.n9_adj_4237 ));
    Odrv4 I__14732 (
            .O(N__61918),
            .I(\c0.n9_adj_4237 ));
    Odrv4 I__14731 (
            .O(N__61915),
            .I(\c0.n9_adj_4237 ));
    Odrv12 I__14730 (
            .O(N__61910),
            .I(\c0.n9_adj_4237 ));
    Odrv4 I__14729 (
            .O(N__61907),
            .I(\c0.n9_adj_4237 ));
    CascadeMux I__14728 (
            .O(N__61894),
            .I(N__61891));
    InMux I__14727 (
            .O(N__61891),
            .I(N__61888));
    LocalMux I__14726 (
            .O(N__61888),
            .I(N__61881));
    InMux I__14725 (
            .O(N__61887),
            .I(N__61878));
    InMux I__14724 (
            .O(N__61886),
            .I(N__61875));
    InMux I__14723 (
            .O(N__61885),
            .I(N__61872));
    InMux I__14722 (
            .O(N__61884),
            .I(N__61869));
    Span12Mux_v I__14721 (
            .O(N__61881),
            .I(N__61866));
    LocalMux I__14720 (
            .O(N__61878),
            .I(N__61861));
    LocalMux I__14719 (
            .O(N__61875),
            .I(N__61861));
    LocalMux I__14718 (
            .O(N__61872),
            .I(\c0.data_in_frame_13_7 ));
    LocalMux I__14717 (
            .O(N__61869),
            .I(\c0.data_in_frame_13_7 ));
    Odrv12 I__14716 (
            .O(N__61866),
            .I(\c0.data_in_frame_13_7 ));
    Odrv12 I__14715 (
            .O(N__61861),
            .I(\c0.data_in_frame_13_7 ));
    InMux I__14714 (
            .O(N__61852),
            .I(N__61849));
    LocalMux I__14713 (
            .O(N__61849),
            .I(N__61845));
    InMux I__14712 (
            .O(N__61848),
            .I(N__61842));
    Span4Mux_v I__14711 (
            .O(N__61845),
            .I(N__61839));
    LocalMux I__14710 (
            .O(N__61842),
            .I(N__61836));
    Span4Mux_v I__14709 (
            .O(N__61839),
            .I(N__61833));
    Odrv12 I__14708 (
            .O(N__61836),
            .I(\c0.n22388 ));
    Odrv4 I__14707 (
            .O(N__61833),
            .I(\c0.n22388 ));
    InMux I__14706 (
            .O(N__61828),
            .I(N__61825));
    LocalMux I__14705 (
            .O(N__61825),
            .I(N__61820));
    InMux I__14704 (
            .O(N__61824),
            .I(N__61817));
    CascadeMux I__14703 (
            .O(N__61823),
            .I(N__61814));
    Span4Mux_v I__14702 (
            .O(N__61820),
            .I(N__61808));
    LocalMux I__14701 (
            .O(N__61817),
            .I(N__61808));
    InMux I__14700 (
            .O(N__61814),
            .I(N__61804));
    InMux I__14699 (
            .O(N__61813),
            .I(N__61801));
    Span4Mux_h I__14698 (
            .O(N__61808),
            .I(N__61798));
    InMux I__14697 (
            .O(N__61807),
            .I(N__61795));
    LocalMux I__14696 (
            .O(N__61804),
            .I(\c0.data_in_frame_17_6 ));
    LocalMux I__14695 (
            .O(N__61801),
            .I(\c0.data_in_frame_17_6 ));
    Odrv4 I__14694 (
            .O(N__61798),
            .I(\c0.data_in_frame_17_6 ));
    LocalMux I__14693 (
            .O(N__61795),
            .I(\c0.data_in_frame_17_6 ));
    InMux I__14692 (
            .O(N__61786),
            .I(N__61783));
    LocalMux I__14691 (
            .O(N__61783),
            .I(N__61780));
    Span4Mux_v I__14690 (
            .O(N__61780),
            .I(N__61777));
    Odrv4 I__14689 (
            .O(N__61777),
            .I(\c0.n20_adj_4247 ));
    InMux I__14688 (
            .O(N__61774),
            .I(N__61770));
    CascadeMux I__14687 (
            .O(N__61773),
            .I(N__61767));
    LocalMux I__14686 (
            .O(N__61770),
            .I(N__61764));
    InMux I__14685 (
            .O(N__61767),
            .I(N__61760));
    Span4Mux_h I__14684 (
            .O(N__61764),
            .I(N__61757));
    InMux I__14683 (
            .O(N__61763),
            .I(N__61754));
    LocalMux I__14682 (
            .O(N__61760),
            .I(\c0.data_in_frame_20_2 ));
    Odrv4 I__14681 (
            .O(N__61757),
            .I(\c0.data_in_frame_20_2 ));
    LocalMux I__14680 (
            .O(N__61754),
            .I(\c0.data_in_frame_20_2 ));
    InMux I__14679 (
            .O(N__61747),
            .I(N__61742));
    InMux I__14678 (
            .O(N__61746),
            .I(N__61738));
    InMux I__14677 (
            .O(N__61745),
            .I(N__61734));
    LocalMux I__14676 (
            .O(N__61742),
            .I(N__61731));
    InMux I__14675 (
            .O(N__61741),
            .I(N__61728));
    LocalMux I__14674 (
            .O(N__61738),
            .I(N__61725));
    InMux I__14673 (
            .O(N__61737),
            .I(N__61722));
    LocalMux I__14672 (
            .O(N__61734),
            .I(N__61715));
    Span4Mux_h I__14671 (
            .O(N__61731),
            .I(N__61715));
    LocalMux I__14670 (
            .O(N__61728),
            .I(N__61715));
    Odrv4 I__14669 (
            .O(N__61725),
            .I(\c0.n13544 ));
    LocalMux I__14668 (
            .O(N__61722),
            .I(\c0.n13544 ));
    Odrv4 I__14667 (
            .O(N__61715),
            .I(\c0.n13544 ));
    CascadeMux I__14666 (
            .O(N__61708),
            .I(N__61705));
    InMux I__14665 (
            .O(N__61705),
            .I(N__61702));
    LocalMux I__14664 (
            .O(N__61702),
            .I(N__61699));
    Span4Mux_v I__14663 (
            .O(N__61699),
            .I(N__61696));
    Span4Mux_v I__14662 (
            .O(N__61696),
            .I(N__61691));
    InMux I__14661 (
            .O(N__61695),
            .I(N__61688));
    InMux I__14660 (
            .O(N__61694),
            .I(N__61685));
    Span4Mux_h I__14659 (
            .O(N__61691),
            .I(N__61682));
    LocalMux I__14658 (
            .O(N__61688),
            .I(N__61679));
    LocalMux I__14657 (
            .O(N__61685),
            .I(data_in_frame_22_3));
    Odrv4 I__14656 (
            .O(N__61682),
            .I(data_in_frame_22_3));
    Odrv4 I__14655 (
            .O(N__61679),
            .I(data_in_frame_22_3));
    InMux I__14654 (
            .O(N__61672),
            .I(N__61669));
    LocalMux I__14653 (
            .O(N__61669),
            .I(N__61663));
    InMux I__14652 (
            .O(N__61668),
            .I(N__61660));
    InMux I__14651 (
            .O(N__61667),
            .I(N__61655));
    InMux I__14650 (
            .O(N__61666),
            .I(N__61655));
    Span4Mux_v I__14649 (
            .O(N__61663),
            .I(N__61652));
    LocalMux I__14648 (
            .O(N__61660),
            .I(N__61647));
    LocalMux I__14647 (
            .O(N__61655),
            .I(N__61647));
    Odrv4 I__14646 (
            .O(N__61652),
            .I(\c0.n23426 ));
    Odrv12 I__14645 (
            .O(N__61647),
            .I(\c0.n23426 ));
    InMux I__14644 (
            .O(N__61642),
            .I(N__61638));
    InMux I__14643 (
            .O(N__61641),
            .I(N__61635));
    LocalMux I__14642 (
            .O(N__61638),
            .I(N__61632));
    LocalMux I__14641 (
            .O(N__61635),
            .I(N__61629));
    Span4Mux_v I__14640 (
            .O(N__61632),
            .I(N__61626));
    Span4Mux_v I__14639 (
            .O(N__61629),
            .I(N__61623));
    Odrv4 I__14638 (
            .O(N__61626),
            .I(\c0.n22007 ));
    Odrv4 I__14637 (
            .O(N__61623),
            .I(\c0.n22007 ));
    InMux I__14636 (
            .O(N__61618),
            .I(N__61612));
    CascadeMux I__14635 (
            .O(N__61617),
            .I(N__61609));
    InMux I__14634 (
            .O(N__61616),
            .I(N__61604));
    InMux I__14633 (
            .O(N__61615),
            .I(N__61604));
    LocalMux I__14632 (
            .O(N__61612),
            .I(N__61600));
    InMux I__14631 (
            .O(N__61609),
            .I(N__61597));
    LocalMux I__14630 (
            .O(N__61604),
            .I(N__61594));
    InMux I__14629 (
            .O(N__61603),
            .I(N__61591));
    Span4Mux_h I__14628 (
            .O(N__61600),
            .I(N__61588));
    LocalMux I__14627 (
            .O(N__61597),
            .I(\c0.data_in_frame_19_6 ));
    Odrv12 I__14626 (
            .O(N__61594),
            .I(\c0.data_in_frame_19_6 ));
    LocalMux I__14625 (
            .O(N__61591),
            .I(\c0.data_in_frame_19_6 ));
    Odrv4 I__14624 (
            .O(N__61588),
            .I(\c0.data_in_frame_19_6 ));
    CascadeMux I__14623 (
            .O(N__61579),
            .I(N__61575));
    InMux I__14622 (
            .O(N__61578),
            .I(N__61572));
    InMux I__14621 (
            .O(N__61575),
            .I(N__61569));
    LocalMux I__14620 (
            .O(N__61572),
            .I(N__61566));
    LocalMux I__14619 (
            .O(N__61569),
            .I(\c0.data_in_frame_18_5 ));
    Odrv12 I__14618 (
            .O(N__61566),
            .I(\c0.data_in_frame_18_5 ));
    InMux I__14617 (
            .O(N__61561),
            .I(N__61558));
    LocalMux I__14616 (
            .O(N__61558),
            .I(N__61555));
    Span4Mux_h I__14615 (
            .O(N__61555),
            .I(N__61552));
    Span4Mux_v I__14614 (
            .O(N__61552),
            .I(N__61549));
    Odrv4 I__14613 (
            .O(N__61549),
            .I(\c0.n22385 ));
    InMux I__14612 (
            .O(N__61546),
            .I(N__61543));
    LocalMux I__14611 (
            .O(N__61543),
            .I(N__61539));
    InMux I__14610 (
            .O(N__61542),
            .I(N__61536));
    Span12Mux_v I__14609 (
            .O(N__61539),
            .I(N__61533));
    LocalMux I__14608 (
            .O(N__61536),
            .I(N__61530));
    Odrv12 I__14607 (
            .O(N__61533),
            .I(\c0.n21126 ));
    Odrv12 I__14606 (
            .O(N__61530),
            .I(\c0.n21126 ));
    CascadeMux I__14605 (
            .O(N__61525),
            .I(N__61522));
    InMux I__14604 (
            .O(N__61522),
            .I(N__61519));
    LocalMux I__14603 (
            .O(N__61519),
            .I(N__61514));
    InMux I__14602 (
            .O(N__61518),
            .I(N__61511));
    InMux I__14601 (
            .O(N__61517),
            .I(N__61508));
    Odrv4 I__14600 (
            .O(N__61514),
            .I(\c0.data_in_frame_16_1 ));
    LocalMux I__14599 (
            .O(N__61511),
            .I(\c0.data_in_frame_16_1 ));
    LocalMux I__14598 (
            .O(N__61508),
            .I(\c0.data_in_frame_16_1 ));
    CascadeMux I__14597 (
            .O(N__61501),
            .I(N__61497));
    CascadeMux I__14596 (
            .O(N__61500),
            .I(N__61493));
    InMux I__14595 (
            .O(N__61497),
            .I(N__61488));
    InMux I__14594 (
            .O(N__61496),
            .I(N__61488));
    InMux I__14593 (
            .O(N__61493),
            .I(N__61485));
    LocalMux I__14592 (
            .O(N__61488),
            .I(N__61482));
    LocalMux I__14591 (
            .O(N__61485),
            .I(N__61476));
    Span4Mux_v I__14590 (
            .O(N__61482),
            .I(N__61476));
    InMux I__14589 (
            .O(N__61481),
            .I(N__61473));
    Odrv4 I__14588 (
            .O(N__61476),
            .I(\c0.data_in_frame_12_3 ));
    LocalMux I__14587 (
            .O(N__61473),
            .I(\c0.data_in_frame_12_3 ));
    InMux I__14586 (
            .O(N__61468),
            .I(N__61464));
    InMux I__14585 (
            .O(N__61467),
            .I(N__61461));
    LocalMux I__14584 (
            .O(N__61464),
            .I(N__61458));
    LocalMux I__14583 (
            .O(N__61461),
            .I(N__61455));
    Span4Mux_v I__14582 (
            .O(N__61458),
            .I(N__61452));
    Span4Mux_h I__14581 (
            .O(N__61455),
            .I(N__61449));
    Span4Mux_h I__14580 (
            .O(N__61452),
            .I(N__61443));
    Span4Mux_v I__14579 (
            .O(N__61449),
            .I(N__61443));
    InMux I__14578 (
            .O(N__61448),
            .I(N__61440));
    Odrv4 I__14577 (
            .O(N__61443),
            .I(\c0.n21975 ));
    LocalMux I__14576 (
            .O(N__61440),
            .I(\c0.n21975 ));
    InMux I__14575 (
            .O(N__61435),
            .I(N__61431));
    InMux I__14574 (
            .O(N__61434),
            .I(N__61427));
    LocalMux I__14573 (
            .O(N__61431),
            .I(N__61424));
    InMux I__14572 (
            .O(N__61430),
            .I(N__61421));
    LocalMux I__14571 (
            .O(N__61427),
            .I(N__61417));
    Span4Mux_v I__14570 (
            .O(N__61424),
            .I(N__61410));
    LocalMux I__14569 (
            .O(N__61421),
            .I(N__61410));
    InMux I__14568 (
            .O(N__61420),
            .I(N__61407));
    Span4Mux_h I__14567 (
            .O(N__61417),
            .I(N__61404));
    InMux I__14566 (
            .O(N__61416),
            .I(N__61399));
    InMux I__14565 (
            .O(N__61415),
            .I(N__61399));
    Odrv4 I__14564 (
            .O(N__61410),
            .I(\c0.data_in_frame_17_2 ));
    LocalMux I__14563 (
            .O(N__61407),
            .I(\c0.data_in_frame_17_2 ));
    Odrv4 I__14562 (
            .O(N__61404),
            .I(\c0.data_in_frame_17_2 ));
    LocalMux I__14561 (
            .O(N__61399),
            .I(\c0.data_in_frame_17_2 ));
    InMux I__14560 (
            .O(N__61390),
            .I(N__61386));
    InMux I__14559 (
            .O(N__61389),
            .I(N__61383));
    LocalMux I__14558 (
            .O(N__61386),
            .I(N__61379));
    LocalMux I__14557 (
            .O(N__61383),
            .I(N__61376));
    InMux I__14556 (
            .O(N__61382),
            .I(N__61373));
    Span4Mux_h I__14555 (
            .O(N__61379),
            .I(N__61370));
    Span12Mux_v I__14554 (
            .O(N__61376),
            .I(N__61367));
    LocalMux I__14553 (
            .O(N__61373),
            .I(\c0.data_in_frame_15_1 ));
    Odrv4 I__14552 (
            .O(N__61370),
            .I(\c0.data_in_frame_15_1 ));
    Odrv12 I__14551 (
            .O(N__61367),
            .I(\c0.data_in_frame_15_1 ));
    CascadeMux I__14550 (
            .O(N__61360),
            .I(N__61356));
    CascadeMux I__14549 (
            .O(N__61359),
            .I(N__61353));
    InMux I__14548 (
            .O(N__61356),
            .I(N__61350));
    InMux I__14547 (
            .O(N__61353),
            .I(N__61347));
    LocalMux I__14546 (
            .O(N__61350),
            .I(N__61344));
    LocalMux I__14545 (
            .O(N__61347),
            .I(N__61338));
    Span4Mux_h I__14544 (
            .O(N__61344),
            .I(N__61338));
    InMux I__14543 (
            .O(N__61343),
            .I(N__61335));
    Odrv4 I__14542 (
            .O(N__61338),
            .I(\c0.data_in_frame_12_4 ));
    LocalMux I__14541 (
            .O(N__61335),
            .I(\c0.data_in_frame_12_4 ));
    CascadeMux I__14540 (
            .O(N__61330),
            .I(N__61326));
    InMux I__14539 (
            .O(N__61329),
            .I(N__61323));
    InMux I__14538 (
            .O(N__61326),
            .I(N__61319));
    LocalMux I__14537 (
            .O(N__61323),
            .I(N__61316));
    InMux I__14536 (
            .O(N__61322),
            .I(N__61313));
    LocalMux I__14535 (
            .O(N__61319),
            .I(N__61307));
    Span4Mux_v I__14534 (
            .O(N__61316),
            .I(N__61307));
    LocalMux I__14533 (
            .O(N__61313),
            .I(N__61304));
    InMux I__14532 (
            .O(N__61312),
            .I(N__61301));
    Odrv4 I__14531 (
            .O(N__61307),
            .I(\c0.data_in_frame_13_3 ));
    Odrv4 I__14530 (
            .O(N__61304),
            .I(\c0.data_in_frame_13_3 ));
    LocalMux I__14529 (
            .O(N__61301),
            .I(\c0.data_in_frame_13_3 ));
    InMux I__14528 (
            .O(N__61294),
            .I(N__61291));
    LocalMux I__14527 (
            .O(N__61291),
            .I(N__61286));
    CascadeMux I__14526 (
            .O(N__61290),
            .I(N__61281));
    InMux I__14525 (
            .O(N__61289),
            .I(N__61278));
    Span4Mux_h I__14524 (
            .O(N__61286),
            .I(N__61275));
    InMux I__14523 (
            .O(N__61285),
            .I(N__61268));
    InMux I__14522 (
            .O(N__61284),
            .I(N__61268));
    InMux I__14521 (
            .O(N__61281),
            .I(N__61268));
    LocalMux I__14520 (
            .O(N__61278),
            .I(\c0.data_in_frame_13_5 ));
    Odrv4 I__14519 (
            .O(N__61275),
            .I(\c0.data_in_frame_13_5 ));
    LocalMux I__14518 (
            .O(N__61268),
            .I(\c0.data_in_frame_13_5 ));
    CascadeMux I__14517 (
            .O(N__61261),
            .I(N__61258));
    InMux I__14516 (
            .O(N__61258),
            .I(N__61255));
    LocalMux I__14515 (
            .O(N__61255),
            .I(N__61251));
    InMux I__14514 (
            .O(N__61254),
            .I(N__61248));
    Odrv12 I__14513 (
            .O(N__61251),
            .I(\c0.n14081 ));
    LocalMux I__14512 (
            .O(N__61248),
            .I(\c0.n14081 ));
    CascadeMux I__14511 (
            .O(N__61243),
            .I(N__61239));
    InMux I__14510 (
            .O(N__61242),
            .I(N__61236));
    InMux I__14509 (
            .O(N__61239),
            .I(N__61232));
    LocalMux I__14508 (
            .O(N__61236),
            .I(N__61229));
    InMux I__14507 (
            .O(N__61235),
            .I(N__61226));
    LocalMux I__14506 (
            .O(N__61232),
            .I(N__61219));
    Span4Mux_h I__14505 (
            .O(N__61229),
            .I(N__61219));
    LocalMux I__14504 (
            .O(N__61226),
            .I(N__61219));
    Odrv4 I__14503 (
            .O(N__61219),
            .I(\c0.data_in_frame_16_0 ));
    CascadeMux I__14502 (
            .O(N__61216),
            .I(N__61213));
    InMux I__14501 (
            .O(N__61213),
            .I(N__61210));
    LocalMux I__14500 (
            .O(N__61210),
            .I(N__61206));
    CascadeMux I__14499 (
            .O(N__61209),
            .I(N__61203));
    Span4Mux_v I__14498 (
            .O(N__61206),
            .I(N__61199));
    InMux I__14497 (
            .O(N__61203),
            .I(N__61196));
    CascadeMux I__14496 (
            .O(N__61202),
            .I(N__61193));
    Span4Mux_h I__14495 (
            .O(N__61199),
            .I(N__61188));
    LocalMux I__14494 (
            .O(N__61196),
            .I(N__61188));
    InMux I__14493 (
            .O(N__61193),
            .I(N__61185));
    Span4Mux_v I__14492 (
            .O(N__61188),
            .I(N__61182));
    LocalMux I__14491 (
            .O(N__61185),
            .I(\c0.data_in_frame_21_7 ));
    Odrv4 I__14490 (
            .O(N__61182),
            .I(\c0.data_in_frame_21_7 ));
    InMux I__14489 (
            .O(N__61177),
            .I(N__61173));
    InMux I__14488 (
            .O(N__61176),
            .I(N__61169));
    LocalMux I__14487 (
            .O(N__61173),
            .I(N__61166));
    InMux I__14486 (
            .O(N__61172),
            .I(N__61163));
    LocalMux I__14485 (
            .O(N__61169),
            .I(\c0.n13210 ));
    Odrv4 I__14484 (
            .O(N__61166),
            .I(\c0.n13210 ));
    LocalMux I__14483 (
            .O(N__61163),
            .I(\c0.n13210 ));
    InMux I__14482 (
            .O(N__61156),
            .I(N__61153));
    LocalMux I__14481 (
            .O(N__61153),
            .I(N__61150));
    Span4Mux_h I__14480 (
            .O(N__61150),
            .I(N__61146));
    InMux I__14479 (
            .O(N__61149),
            .I(N__61143));
    Odrv4 I__14478 (
            .O(N__61146),
            .I(\c0.n22091 ));
    LocalMux I__14477 (
            .O(N__61143),
            .I(\c0.n22091 ));
    InMux I__14476 (
            .O(N__61138),
            .I(N__61135));
    LocalMux I__14475 (
            .O(N__61135),
            .I(N__61132));
    Span4Mux_v I__14474 (
            .O(N__61132),
            .I(N__61128));
    InMux I__14473 (
            .O(N__61131),
            .I(N__61125));
    Sp12to4 I__14472 (
            .O(N__61128),
            .I(N__61119));
    LocalMux I__14471 (
            .O(N__61125),
            .I(N__61119));
    InMux I__14470 (
            .O(N__61124),
            .I(N__61116));
    Odrv12 I__14469 (
            .O(N__61119),
            .I(\c0.n21934 ));
    LocalMux I__14468 (
            .O(N__61116),
            .I(\c0.n21934 ));
    InMux I__14467 (
            .O(N__61111),
            .I(N__61108));
    LocalMux I__14466 (
            .O(N__61108),
            .I(N__61104));
    InMux I__14465 (
            .O(N__61107),
            .I(N__61100));
    Span4Mux_h I__14464 (
            .O(N__61104),
            .I(N__61097));
    InMux I__14463 (
            .O(N__61103),
            .I(N__61094));
    LocalMux I__14462 (
            .O(N__61100),
            .I(N__61089));
    Span4Mux_h I__14461 (
            .O(N__61097),
            .I(N__61084));
    LocalMux I__14460 (
            .O(N__61094),
            .I(N__61084));
    InMux I__14459 (
            .O(N__61093),
            .I(N__61079));
    InMux I__14458 (
            .O(N__61092),
            .I(N__61079));
    Odrv12 I__14457 (
            .O(N__61089),
            .I(\c0.data_in_frame_4_5 ));
    Odrv4 I__14456 (
            .O(N__61084),
            .I(\c0.data_in_frame_4_5 ));
    LocalMux I__14455 (
            .O(N__61079),
            .I(\c0.data_in_frame_4_5 ));
    CascadeMux I__14454 (
            .O(N__61072),
            .I(N__61069));
    InMux I__14453 (
            .O(N__61069),
            .I(N__61066));
    LocalMux I__14452 (
            .O(N__61066),
            .I(N__61063));
    Span4Mux_v I__14451 (
            .O(N__61063),
            .I(N__61059));
    InMux I__14450 (
            .O(N__61062),
            .I(N__61056));
    Span4Mux_h I__14449 (
            .O(N__61059),
            .I(N__61051));
    LocalMux I__14448 (
            .O(N__61056),
            .I(N__61051));
    Span4Mux_h I__14447 (
            .O(N__61051),
            .I(N__61048));
    Odrv4 I__14446 (
            .O(N__61048),
            .I(\c0.n13421 ));
    CascadeMux I__14445 (
            .O(N__61045),
            .I(N__61041));
    InMux I__14444 (
            .O(N__61044),
            .I(N__61037));
    InMux I__14443 (
            .O(N__61041),
            .I(N__61032));
    InMux I__14442 (
            .O(N__61040),
            .I(N__61032));
    LocalMux I__14441 (
            .O(N__61037),
            .I(\c0.data_in_frame_11_4 ));
    LocalMux I__14440 (
            .O(N__61032),
            .I(\c0.data_in_frame_11_4 ));
    CascadeMux I__14439 (
            .O(N__61027),
            .I(\c0.n13421_cascade_ ));
    InMux I__14438 (
            .O(N__61024),
            .I(N__61020));
    InMux I__14437 (
            .O(N__61023),
            .I(N__61017));
    LocalMux I__14436 (
            .O(N__61020),
            .I(N__61014));
    LocalMux I__14435 (
            .O(N__61017),
            .I(N__61011));
    Span4Mux_h I__14434 (
            .O(N__61014),
            .I(N__61008));
    Odrv12 I__14433 (
            .O(N__61011),
            .I(\c0.n22069 ));
    Odrv4 I__14432 (
            .O(N__61008),
            .I(\c0.n22069 ));
    InMux I__14431 (
            .O(N__61003),
            .I(N__61000));
    LocalMux I__14430 (
            .O(N__61000),
            .I(\c0.n10_adj_4252 ));
    CascadeMux I__14429 (
            .O(N__60997),
            .I(N__60993));
    InMux I__14428 (
            .O(N__60996),
            .I(N__60990));
    InMux I__14427 (
            .O(N__60993),
            .I(N__60986));
    LocalMux I__14426 (
            .O(N__60990),
            .I(N__60983));
    InMux I__14425 (
            .O(N__60989),
            .I(N__60980));
    LocalMux I__14424 (
            .O(N__60986),
            .I(\c0.data_in_frame_7_2 ));
    Odrv4 I__14423 (
            .O(N__60983),
            .I(\c0.data_in_frame_7_2 ));
    LocalMux I__14422 (
            .O(N__60980),
            .I(\c0.data_in_frame_7_2 ));
    InMux I__14421 (
            .O(N__60973),
            .I(N__60969));
    InMux I__14420 (
            .O(N__60972),
            .I(N__60966));
    LocalMux I__14419 (
            .O(N__60969),
            .I(N__60963));
    LocalMux I__14418 (
            .O(N__60966),
            .I(\c0.n22343 ));
    Odrv12 I__14417 (
            .O(N__60963),
            .I(\c0.n22343 ));
    InMux I__14416 (
            .O(N__60958),
            .I(N__60955));
    LocalMux I__14415 (
            .O(N__60955),
            .I(N__60952));
    Odrv4 I__14414 (
            .O(N__60952),
            .I(\c0.n10_adj_4267 ));
    CascadeMux I__14413 (
            .O(N__60949),
            .I(N__60944));
    CascadeMux I__14412 (
            .O(N__60948),
            .I(N__60941));
    InMux I__14411 (
            .O(N__60947),
            .I(N__60938));
    InMux I__14410 (
            .O(N__60944),
            .I(N__60934));
    InMux I__14409 (
            .O(N__60941),
            .I(N__60931));
    LocalMux I__14408 (
            .O(N__60938),
            .I(N__60928));
    InMux I__14407 (
            .O(N__60937),
            .I(N__60925));
    LocalMux I__14406 (
            .O(N__60934),
            .I(N__60922));
    LocalMux I__14405 (
            .O(N__60931),
            .I(N__60915));
    Span4Mux_v I__14404 (
            .O(N__60928),
            .I(N__60915));
    LocalMux I__14403 (
            .O(N__60925),
            .I(N__60915));
    Span4Mux_h I__14402 (
            .O(N__60922),
            .I(N__60912));
    Odrv4 I__14401 (
            .O(N__60915),
            .I(\c0.data_in_frame_12_5 ));
    Odrv4 I__14400 (
            .O(N__60912),
            .I(\c0.data_in_frame_12_5 ));
    InMux I__14399 (
            .O(N__60907),
            .I(N__60904));
    LocalMux I__14398 (
            .O(N__60904),
            .I(N__60901));
    Odrv4 I__14397 (
            .O(N__60901),
            .I(\c0.n16_adj_4268 ));
    InMux I__14396 (
            .O(N__60898),
            .I(N__60884));
    InMux I__14395 (
            .O(N__60897),
            .I(N__60878));
    InMux I__14394 (
            .O(N__60896),
            .I(N__60871));
    InMux I__14393 (
            .O(N__60895),
            .I(N__60871));
    InMux I__14392 (
            .O(N__60894),
            .I(N__60871));
    CascadeMux I__14391 (
            .O(N__60893),
            .I(N__60864));
    InMux I__14390 (
            .O(N__60892),
            .I(N__60856));
    InMux I__14389 (
            .O(N__60891),
            .I(N__60856));
    InMux I__14388 (
            .O(N__60890),
            .I(N__60856));
    InMux I__14387 (
            .O(N__60889),
            .I(N__60853));
    InMux I__14386 (
            .O(N__60888),
            .I(N__60839));
    CascadeMux I__14385 (
            .O(N__60887),
            .I(N__60836));
    LocalMux I__14384 (
            .O(N__60884),
            .I(N__60831));
    InMux I__14383 (
            .O(N__60883),
            .I(N__60824));
    InMux I__14382 (
            .O(N__60882),
            .I(N__60824));
    InMux I__14381 (
            .O(N__60881),
            .I(N__60824));
    LocalMux I__14380 (
            .O(N__60878),
            .I(N__60820));
    LocalMux I__14379 (
            .O(N__60871),
            .I(N__60817));
    InMux I__14378 (
            .O(N__60870),
            .I(N__60808));
    InMux I__14377 (
            .O(N__60869),
            .I(N__60808));
    InMux I__14376 (
            .O(N__60868),
            .I(N__60808));
    InMux I__14375 (
            .O(N__60867),
            .I(N__60808));
    InMux I__14374 (
            .O(N__60864),
            .I(N__60803));
    InMux I__14373 (
            .O(N__60863),
            .I(N__60800));
    LocalMux I__14372 (
            .O(N__60856),
            .I(N__60795));
    LocalMux I__14371 (
            .O(N__60853),
            .I(N__60795));
    InMux I__14370 (
            .O(N__60852),
            .I(N__60784));
    InMux I__14369 (
            .O(N__60851),
            .I(N__60784));
    InMux I__14368 (
            .O(N__60850),
            .I(N__60784));
    InMux I__14367 (
            .O(N__60849),
            .I(N__60784));
    InMux I__14366 (
            .O(N__60848),
            .I(N__60784));
    InMux I__14365 (
            .O(N__60847),
            .I(N__60777));
    InMux I__14364 (
            .O(N__60846),
            .I(N__60777));
    InMux I__14363 (
            .O(N__60845),
            .I(N__60777));
    InMux I__14362 (
            .O(N__60844),
            .I(N__60770));
    InMux I__14361 (
            .O(N__60843),
            .I(N__60770));
    InMux I__14360 (
            .O(N__60842),
            .I(N__60770));
    LocalMux I__14359 (
            .O(N__60839),
            .I(N__60767));
    InMux I__14358 (
            .O(N__60836),
            .I(N__60752));
    InMux I__14357 (
            .O(N__60835),
            .I(N__60747));
    InMux I__14356 (
            .O(N__60834),
            .I(N__60747));
    Span4Mux_h I__14355 (
            .O(N__60831),
            .I(N__60742));
    LocalMux I__14354 (
            .O(N__60824),
            .I(N__60742));
    InMux I__14353 (
            .O(N__60823),
            .I(N__60739));
    Span4Mux_h I__14352 (
            .O(N__60820),
            .I(N__60734));
    Span4Mux_v I__14351 (
            .O(N__60817),
            .I(N__60734));
    LocalMux I__14350 (
            .O(N__60808),
            .I(N__60731));
    InMux I__14349 (
            .O(N__60807),
            .I(N__60728));
    InMux I__14348 (
            .O(N__60806),
            .I(N__60724));
    LocalMux I__14347 (
            .O(N__60803),
            .I(N__60719));
    LocalMux I__14346 (
            .O(N__60800),
            .I(N__60719));
    Span4Mux_v I__14345 (
            .O(N__60795),
            .I(N__60716));
    LocalMux I__14344 (
            .O(N__60784),
            .I(N__60708));
    LocalMux I__14343 (
            .O(N__60777),
            .I(N__60708));
    LocalMux I__14342 (
            .O(N__60770),
            .I(N__60703));
    Span4Mux_h I__14341 (
            .O(N__60767),
            .I(N__60703));
    InMux I__14340 (
            .O(N__60766),
            .I(N__60688));
    InMux I__14339 (
            .O(N__60765),
            .I(N__60688));
    InMux I__14338 (
            .O(N__60764),
            .I(N__60688));
    InMux I__14337 (
            .O(N__60763),
            .I(N__60688));
    InMux I__14336 (
            .O(N__60762),
            .I(N__60688));
    InMux I__14335 (
            .O(N__60761),
            .I(N__60688));
    InMux I__14334 (
            .O(N__60760),
            .I(N__60688));
    InMux I__14333 (
            .O(N__60759),
            .I(N__60685));
    InMux I__14332 (
            .O(N__60758),
            .I(N__60676));
    InMux I__14331 (
            .O(N__60757),
            .I(N__60676));
    InMux I__14330 (
            .O(N__60756),
            .I(N__60676));
    InMux I__14329 (
            .O(N__60755),
            .I(N__60676));
    LocalMux I__14328 (
            .O(N__60752),
            .I(N__60673));
    LocalMux I__14327 (
            .O(N__60747),
            .I(N__60668));
    Span4Mux_h I__14326 (
            .O(N__60742),
            .I(N__60668));
    LocalMux I__14325 (
            .O(N__60739),
            .I(N__60661));
    Span4Mux_h I__14324 (
            .O(N__60734),
            .I(N__60661));
    Span4Mux_v I__14323 (
            .O(N__60731),
            .I(N__60661));
    LocalMux I__14322 (
            .O(N__60728),
            .I(N__60658));
    InMux I__14321 (
            .O(N__60727),
            .I(N__60655));
    LocalMux I__14320 (
            .O(N__60724),
            .I(N__60652));
    Span4Mux_v I__14319 (
            .O(N__60719),
            .I(N__60649));
    Span4Mux_v I__14318 (
            .O(N__60716),
            .I(N__60646));
    InMux I__14317 (
            .O(N__60715),
            .I(N__60639));
    InMux I__14316 (
            .O(N__60714),
            .I(N__60634));
    InMux I__14315 (
            .O(N__60713),
            .I(N__60634));
    Span4Mux_v I__14314 (
            .O(N__60708),
            .I(N__60629));
    Span4Mux_v I__14313 (
            .O(N__60703),
            .I(N__60629));
    LocalMux I__14312 (
            .O(N__60688),
            .I(N__60624));
    LocalMux I__14311 (
            .O(N__60685),
            .I(N__60624));
    LocalMux I__14310 (
            .O(N__60676),
            .I(N__60617));
    Span4Mux_h I__14309 (
            .O(N__60673),
            .I(N__60617));
    Span4Mux_v I__14308 (
            .O(N__60668),
            .I(N__60617));
    Span4Mux_v I__14307 (
            .O(N__60661),
            .I(N__60614));
    Span12Mux_v I__14306 (
            .O(N__60658),
            .I(N__60611));
    LocalMux I__14305 (
            .O(N__60655),
            .I(N__60602));
    Span4Mux_v I__14304 (
            .O(N__60652),
            .I(N__60602));
    Span4Mux_h I__14303 (
            .O(N__60649),
            .I(N__60602));
    Span4Mux_h I__14302 (
            .O(N__60646),
            .I(N__60602));
    InMux I__14301 (
            .O(N__60645),
            .I(N__60593));
    InMux I__14300 (
            .O(N__60644),
            .I(N__60593));
    InMux I__14299 (
            .O(N__60643),
            .I(N__60593));
    InMux I__14298 (
            .O(N__60642),
            .I(N__60593));
    LocalMux I__14297 (
            .O(N__60639),
            .I(\c0.n21740 ));
    LocalMux I__14296 (
            .O(N__60634),
            .I(\c0.n21740 ));
    Odrv4 I__14295 (
            .O(N__60629),
            .I(\c0.n21740 ));
    Odrv12 I__14294 (
            .O(N__60624),
            .I(\c0.n21740 ));
    Odrv4 I__14293 (
            .O(N__60617),
            .I(\c0.n21740 ));
    Odrv4 I__14292 (
            .O(N__60614),
            .I(\c0.n21740 ));
    Odrv12 I__14291 (
            .O(N__60611),
            .I(\c0.n21740 ));
    Odrv4 I__14290 (
            .O(N__60602),
            .I(\c0.n21740 ));
    LocalMux I__14289 (
            .O(N__60593),
            .I(\c0.n21740 ));
    InMux I__14288 (
            .O(N__60574),
            .I(N__60571));
    LocalMux I__14287 (
            .O(N__60571),
            .I(N__60568));
    Span4Mux_h I__14286 (
            .O(N__60568),
            .I(N__60563));
    InMux I__14285 (
            .O(N__60567),
            .I(N__60558));
    InMux I__14284 (
            .O(N__60566),
            .I(N__60558));
    Odrv4 I__14283 (
            .O(N__60563),
            .I(\c0.data_in_frame_7_0 ));
    LocalMux I__14282 (
            .O(N__60558),
            .I(\c0.data_in_frame_7_0 ));
    InMux I__14281 (
            .O(N__60553),
            .I(N__60550));
    LocalMux I__14280 (
            .O(N__60550),
            .I(N__60547));
    Span4Mux_h I__14279 (
            .O(N__60547),
            .I(N__60543));
    InMux I__14278 (
            .O(N__60546),
            .I(N__60540));
    Odrv4 I__14277 (
            .O(N__60543),
            .I(\c0.n21845 ));
    LocalMux I__14276 (
            .O(N__60540),
            .I(\c0.n21845 ));
    InMux I__14275 (
            .O(N__60535),
            .I(N__60532));
    LocalMux I__14274 (
            .O(N__60532),
            .I(N__60528));
    InMux I__14273 (
            .O(N__60531),
            .I(N__60525));
    Odrv4 I__14272 (
            .O(N__60528),
            .I(\c0.n22781 ));
    LocalMux I__14271 (
            .O(N__60525),
            .I(\c0.n22781 ));
    InMux I__14270 (
            .O(N__60520),
            .I(N__60516));
    CascadeMux I__14269 (
            .O(N__60519),
            .I(N__60513));
    LocalMux I__14268 (
            .O(N__60516),
            .I(N__60508));
    InMux I__14267 (
            .O(N__60513),
            .I(N__60503));
    InMux I__14266 (
            .O(N__60512),
            .I(N__60503));
    InMux I__14265 (
            .O(N__60511),
            .I(N__60500));
    Span4Mux_h I__14264 (
            .O(N__60508),
            .I(N__60497));
    LocalMux I__14263 (
            .O(N__60503),
            .I(\c0.data_in_frame_11_1 ));
    LocalMux I__14262 (
            .O(N__60500),
            .I(\c0.data_in_frame_11_1 ));
    Odrv4 I__14261 (
            .O(N__60497),
            .I(\c0.data_in_frame_11_1 ));
    InMux I__14260 (
            .O(N__60490),
            .I(N__60486));
    InMux I__14259 (
            .O(N__60489),
            .I(N__60483));
    LocalMux I__14258 (
            .O(N__60486),
            .I(N__60479));
    LocalMux I__14257 (
            .O(N__60483),
            .I(N__60476));
    CascadeMux I__14256 (
            .O(N__60482),
            .I(N__60473));
    Span4Mux_v I__14255 (
            .O(N__60479),
            .I(N__60470));
    Span4Mux_v I__14254 (
            .O(N__60476),
            .I(N__60467));
    InMux I__14253 (
            .O(N__60473),
            .I(N__60464));
    Span4Mux_v I__14252 (
            .O(N__60470),
            .I(N__60461));
    Span4Mux_v I__14251 (
            .O(N__60467),
            .I(N__60458));
    LocalMux I__14250 (
            .O(N__60464),
            .I(\c0.data_in_frame_23_3 ));
    Odrv4 I__14249 (
            .O(N__60461),
            .I(\c0.data_in_frame_23_3 ));
    Odrv4 I__14248 (
            .O(N__60458),
            .I(\c0.data_in_frame_23_3 ));
    InMux I__14247 (
            .O(N__60451),
            .I(N__60447));
    InMux I__14246 (
            .O(N__60450),
            .I(N__60444));
    LocalMux I__14245 (
            .O(N__60447),
            .I(N__60441));
    LocalMux I__14244 (
            .O(N__60444),
            .I(\c0.n22236 ));
    Odrv4 I__14243 (
            .O(N__60441),
            .I(\c0.n22236 ));
    InMux I__14242 (
            .O(N__60436),
            .I(N__60432));
    InMux I__14241 (
            .O(N__60435),
            .I(N__60429));
    LocalMux I__14240 (
            .O(N__60432),
            .I(N__60426));
    LocalMux I__14239 (
            .O(N__60429),
            .I(\c0.n4 ));
    Odrv12 I__14238 (
            .O(N__60426),
            .I(\c0.n4 ));
    CascadeMux I__14237 (
            .O(N__60421),
            .I(N__60418));
    InMux I__14236 (
            .O(N__60418),
            .I(N__60415));
    LocalMux I__14235 (
            .O(N__60415),
            .I(\c0.n5965 ));
    InMux I__14234 (
            .O(N__60412),
            .I(N__60409));
    LocalMux I__14233 (
            .O(N__60409),
            .I(\c0.n8_adj_4275 ));
    InMux I__14232 (
            .O(N__60406),
            .I(N__60403));
    LocalMux I__14231 (
            .O(N__60403),
            .I(\c0.n8_adj_4276 ));
    InMux I__14230 (
            .O(N__60400),
            .I(N__60395));
    InMux I__14229 (
            .O(N__60399),
            .I(N__60392));
    CascadeMux I__14228 (
            .O(N__60398),
            .I(N__60389));
    LocalMux I__14227 (
            .O(N__60395),
            .I(N__60384));
    LocalMux I__14226 (
            .O(N__60392),
            .I(N__60384));
    InMux I__14225 (
            .O(N__60389),
            .I(N__60380));
    Span4Mux_v I__14224 (
            .O(N__60384),
            .I(N__60377));
    InMux I__14223 (
            .O(N__60383),
            .I(N__60374));
    LocalMux I__14222 (
            .O(N__60380),
            .I(\c0.data_in_frame_13_0 ));
    Odrv4 I__14221 (
            .O(N__60377),
            .I(\c0.data_in_frame_13_0 ));
    LocalMux I__14220 (
            .O(N__60374),
            .I(\c0.data_in_frame_13_0 ));
    InMux I__14219 (
            .O(N__60367),
            .I(N__60364));
    LocalMux I__14218 (
            .O(N__60364),
            .I(N__60360));
    InMux I__14217 (
            .O(N__60363),
            .I(N__60357));
    Span4Mux_v I__14216 (
            .O(N__60360),
            .I(N__60351));
    LocalMux I__14215 (
            .O(N__60357),
            .I(N__60351));
    InMux I__14214 (
            .O(N__60356),
            .I(N__60348));
    Span4Mux_h I__14213 (
            .O(N__60351),
            .I(N__60345));
    LocalMux I__14212 (
            .O(N__60348),
            .I(\c0.data_in_frame_12_7 ));
    Odrv4 I__14211 (
            .O(N__60345),
            .I(\c0.data_in_frame_12_7 ));
    InMux I__14210 (
            .O(N__60340),
            .I(N__60337));
    LocalMux I__14209 (
            .O(N__60337),
            .I(N__60334));
    Span4Mux_h I__14208 (
            .O(N__60334),
            .I(N__60330));
    InMux I__14207 (
            .O(N__60333),
            .I(N__60326));
    Span4Mux_v I__14206 (
            .O(N__60330),
            .I(N__60323));
    InMux I__14205 (
            .O(N__60329),
            .I(N__60320));
    LocalMux I__14204 (
            .O(N__60326),
            .I(\c0.data_in_frame_23_1 ));
    Odrv4 I__14203 (
            .O(N__60323),
            .I(\c0.data_in_frame_23_1 ));
    LocalMux I__14202 (
            .O(N__60320),
            .I(\c0.data_in_frame_23_1 ));
    InMux I__14201 (
            .O(N__60313),
            .I(N__60305));
    InMux I__14200 (
            .O(N__60312),
            .I(N__60305));
    InMux I__14199 (
            .O(N__60311),
            .I(N__60302));
    InMux I__14198 (
            .O(N__60310),
            .I(N__60299));
    LocalMux I__14197 (
            .O(N__60305),
            .I(N__60296));
    LocalMux I__14196 (
            .O(N__60302),
            .I(N__60293));
    LocalMux I__14195 (
            .O(N__60299),
            .I(N__60290));
    Span4Mux_v I__14194 (
            .O(N__60296),
            .I(N__60287));
    Span4Mux_h I__14193 (
            .O(N__60293),
            .I(N__60284));
    Odrv4 I__14192 (
            .O(N__60290),
            .I(data_in_frame_22_7));
    Odrv4 I__14191 (
            .O(N__60287),
            .I(data_in_frame_22_7));
    Odrv4 I__14190 (
            .O(N__60284),
            .I(data_in_frame_22_7));
    CascadeMux I__14189 (
            .O(N__60277),
            .I(N__60274));
    InMux I__14188 (
            .O(N__60274),
            .I(N__60271));
    LocalMux I__14187 (
            .O(N__60271),
            .I(N__60268));
    Span4Mux_h I__14186 (
            .O(N__60268),
            .I(N__60265));
    Span4Mux_v I__14185 (
            .O(N__60265),
            .I(N__60262));
    Odrv4 I__14184 (
            .O(N__60262),
            .I(\c0.n21995 ));
    CascadeMux I__14183 (
            .O(N__60259),
            .I(N__60256));
    InMux I__14182 (
            .O(N__60256),
            .I(N__60250));
    InMux I__14181 (
            .O(N__60255),
            .I(N__60245));
    InMux I__14180 (
            .O(N__60254),
            .I(N__60245));
    InMux I__14179 (
            .O(N__60253),
            .I(N__60242));
    LocalMux I__14178 (
            .O(N__60250),
            .I(\c0.data_in_frame_12_1 ));
    LocalMux I__14177 (
            .O(N__60245),
            .I(\c0.data_in_frame_12_1 ));
    LocalMux I__14176 (
            .O(N__60242),
            .I(\c0.data_in_frame_12_1 ));
    InMux I__14175 (
            .O(N__60235),
            .I(N__60229));
    InMux I__14174 (
            .O(N__60234),
            .I(N__60226));
    InMux I__14173 (
            .O(N__60233),
            .I(N__60223));
    InMux I__14172 (
            .O(N__60232),
            .I(N__60220));
    LocalMux I__14171 (
            .O(N__60229),
            .I(\c0.data_in_frame_12_2 ));
    LocalMux I__14170 (
            .O(N__60226),
            .I(\c0.data_in_frame_12_2 ));
    LocalMux I__14169 (
            .O(N__60223),
            .I(\c0.data_in_frame_12_2 ));
    LocalMux I__14168 (
            .O(N__60220),
            .I(\c0.data_in_frame_12_2 ));
    CascadeMux I__14167 (
            .O(N__60211),
            .I(N__60208));
    InMux I__14166 (
            .O(N__60208),
            .I(N__60204));
    InMux I__14165 (
            .O(N__60207),
            .I(N__60201));
    LocalMux I__14164 (
            .O(N__60204),
            .I(\c0.data_in_frame_13_2 ));
    LocalMux I__14163 (
            .O(N__60201),
            .I(\c0.data_in_frame_13_2 ));
    InMux I__14162 (
            .O(N__60196),
            .I(N__60192));
    CascadeMux I__14161 (
            .O(N__60195),
            .I(N__60188));
    LocalMux I__14160 (
            .O(N__60192),
            .I(N__60185));
    InMux I__14159 (
            .O(N__60191),
            .I(N__60182));
    InMux I__14158 (
            .O(N__60188),
            .I(N__60179));
    Span4Mux_h I__14157 (
            .O(N__60185),
            .I(N__60176));
    LocalMux I__14156 (
            .O(N__60182),
            .I(N__60173));
    LocalMux I__14155 (
            .O(N__60179),
            .I(N__60169));
    Span4Mux_v I__14154 (
            .O(N__60176),
            .I(N__60164));
    Span4Mux_h I__14153 (
            .O(N__60173),
            .I(N__60164));
    InMux I__14152 (
            .O(N__60172),
            .I(N__60161));
    Odrv4 I__14151 (
            .O(N__60169),
            .I(\c0.data_in_frame_13_1 ));
    Odrv4 I__14150 (
            .O(N__60164),
            .I(\c0.data_in_frame_13_1 ));
    LocalMux I__14149 (
            .O(N__60161),
            .I(\c0.data_in_frame_13_1 ));
    CascadeMux I__14148 (
            .O(N__60154),
            .I(N__60151));
    InMux I__14147 (
            .O(N__60151),
            .I(N__60147));
    CascadeMux I__14146 (
            .O(N__60150),
            .I(N__60144));
    LocalMux I__14145 (
            .O(N__60147),
            .I(N__60140));
    InMux I__14144 (
            .O(N__60144),
            .I(N__60134));
    InMux I__14143 (
            .O(N__60143),
            .I(N__60134));
    Span4Mux_h I__14142 (
            .O(N__60140),
            .I(N__60131));
    InMux I__14141 (
            .O(N__60139),
            .I(N__60128));
    LocalMux I__14140 (
            .O(N__60134),
            .I(\c0.data_in_frame_11_0 ));
    Odrv4 I__14139 (
            .O(N__60131),
            .I(\c0.data_in_frame_11_0 ));
    LocalMux I__14138 (
            .O(N__60128),
            .I(\c0.data_in_frame_11_0 ));
    InMux I__14137 (
            .O(N__60121),
            .I(N__60118));
    LocalMux I__14136 (
            .O(N__60118),
            .I(N__60114));
    InMux I__14135 (
            .O(N__60117),
            .I(N__60111));
    Span4Mux_h I__14134 (
            .O(N__60114),
            .I(N__60108));
    LocalMux I__14133 (
            .O(N__60111),
            .I(\c0.n22274 ));
    Odrv4 I__14132 (
            .O(N__60108),
            .I(\c0.n22274 ));
    InMux I__14131 (
            .O(N__60103),
            .I(N__60098));
    InMux I__14130 (
            .O(N__60102),
            .I(N__60095));
    InMux I__14129 (
            .O(N__60101),
            .I(N__60091));
    LocalMux I__14128 (
            .O(N__60098),
            .I(N__60088));
    LocalMux I__14127 (
            .O(N__60095),
            .I(N__60085));
    CascadeMux I__14126 (
            .O(N__60094),
            .I(N__60082));
    LocalMux I__14125 (
            .O(N__60091),
            .I(N__60078));
    Span4Mux_v I__14124 (
            .O(N__60088),
            .I(N__60073));
    Span4Mux_h I__14123 (
            .O(N__60085),
            .I(N__60073));
    InMux I__14122 (
            .O(N__60082),
            .I(N__60068));
    InMux I__14121 (
            .O(N__60081),
            .I(N__60068));
    Odrv12 I__14120 (
            .O(N__60078),
            .I(\c0.data_in_frame_10_6 ));
    Odrv4 I__14119 (
            .O(N__60073),
            .I(\c0.data_in_frame_10_6 ));
    LocalMux I__14118 (
            .O(N__60068),
            .I(\c0.data_in_frame_10_6 ));
    CascadeMux I__14117 (
            .O(N__60061),
            .I(\c0.n13999_cascade_ ));
    InMux I__14116 (
            .O(N__60058),
            .I(N__60055));
    LocalMux I__14115 (
            .O(N__60055),
            .I(N__60051));
    InMux I__14114 (
            .O(N__60054),
            .I(N__60048));
    Span4Mux_h I__14113 (
            .O(N__60051),
            .I(N__60045));
    LocalMux I__14112 (
            .O(N__60048),
            .I(N__60042));
    Odrv4 I__14111 (
            .O(N__60045),
            .I(\c0.n21940 ));
    Odrv4 I__14110 (
            .O(N__60042),
            .I(\c0.n21940 ));
    CascadeMux I__14109 (
            .O(N__60037),
            .I(N__60034));
    InMux I__14108 (
            .O(N__60034),
            .I(N__60031));
    LocalMux I__14107 (
            .O(N__60031),
            .I(N__60027));
    InMux I__14106 (
            .O(N__60030),
            .I(N__60024));
    Span4Mux_h I__14105 (
            .O(N__60027),
            .I(N__60021));
    LocalMux I__14104 (
            .O(N__60024),
            .I(N__60018));
    Span4Mux_v I__14103 (
            .O(N__60021),
            .I(N__60015));
    Span4Mux_h I__14102 (
            .O(N__60018),
            .I(N__60012));
    Odrv4 I__14101 (
            .O(N__60015),
            .I(\c0.n13233 ));
    Odrv4 I__14100 (
            .O(N__60012),
            .I(\c0.n13233 ));
    InMux I__14099 (
            .O(N__60007),
            .I(N__60004));
    LocalMux I__14098 (
            .O(N__60004),
            .I(N__59999));
    InMux I__14097 (
            .O(N__60003),
            .I(N__59996));
    InMux I__14096 (
            .O(N__60002),
            .I(N__59993));
    Span4Mux_h I__14095 (
            .O(N__59999),
            .I(N__59990));
    LocalMux I__14094 (
            .O(N__59996),
            .I(\c0.data_in_frame_9_2 ));
    LocalMux I__14093 (
            .O(N__59993),
            .I(\c0.data_in_frame_9_2 ));
    Odrv4 I__14092 (
            .O(N__59990),
            .I(\c0.data_in_frame_9_2 ));
    InMux I__14091 (
            .O(N__59983),
            .I(N__59980));
    LocalMux I__14090 (
            .O(N__59980),
            .I(N__59977));
    Span4Mux_v I__14089 (
            .O(N__59977),
            .I(N__59973));
    InMux I__14088 (
            .O(N__59976),
            .I(N__59970));
    Odrv4 I__14087 (
            .O(N__59973),
            .I(\c0.n13993 ));
    LocalMux I__14086 (
            .O(N__59970),
            .I(\c0.n13993 ));
    InMux I__14085 (
            .O(N__59965),
            .I(N__59962));
    LocalMux I__14084 (
            .O(N__59962),
            .I(N__59959));
    Span4Mux_h I__14083 (
            .O(N__59959),
            .I(N__59954));
    InMux I__14082 (
            .O(N__59958),
            .I(N__59949));
    InMux I__14081 (
            .O(N__59957),
            .I(N__59949));
    Odrv4 I__14080 (
            .O(N__59954),
            .I(n91));
    LocalMux I__14079 (
            .O(N__59949),
            .I(n91));
    InMux I__14078 (
            .O(N__59944),
            .I(N__59941));
    LocalMux I__14077 (
            .O(N__59941),
            .I(N__59936));
    InMux I__14076 (
            .O(N__59940),
            .I(N__59933));
    InMux I__14075 (
            .O(N__59939),
            .I(N__59930));
    Span4Mux_v I__14074 (
            .O(N__59936),
            .I(N__59925));
    LocalMux I__14073 (
            .O(N__59933),
            .I(N__59925));
    LocalMux I__14072 (
            .O(N__59930),
            .I(N__59922));
    Span4Mux_h I__14071 (
            .O(N__59925),
            .I(N__59919));
    Span4Mux_v I__14070 (
            .O(N__59922),
            .I(N__59914));
    Span4Mux_v I__14069 (
            .O(N__59919),
            .I(N__59914));
    Odrv4 I__14068 (
            .O(N__59914),
            .I(n12973));
    InMux I__14067 (
            .O(N__59911),
            .I(N__59907));
    InMux I__14066 (
            .O(N__59910),
            .I(N__59904));
    LocalMux I__14065 (
            .O(N__59907),
            .I(n14917));
    LocalMux I__14064 (
            .O(N__59904),
            .I(n14917));
    InMux I__14063 (
            .O(N__59899),
            .I(N__59894));
    InMux I__14062 (
            .O(N__59898),
            .I(N__59889));
    InMux I__14061 (
            .O(N__59897),
            .I(N__59889));
    LocalMux I__14060 (
            .O(N__59894),
            .I(n14436));
    LocalMux I__14059 (
            .O(N__59889),
            .I(n14436));
    InMux I__14058 (
            .O(N__59884),
            .I(N__59880));
    InMux I__14057 (
            .O(N__59883),
            .I(N__59877));
    LocalMux I__14056 (
            .O(N__59880),
            .I(N__59874));
    LocalMux I__14055 (
            .O(N__59877),
            .I(N__59869));
    Span4Mux_v I__14054 (
            .O(N__59874),
            .I(N__59869));
    Span4Mux_h I__14053 (
            .O(N__59869),
            .I(N__59865));
    CascadeMux I__14052 (
            .O(N__59868),
            .I(N__59860));
    Span4Mux_v I__14051 (
            .O(N__59865),
            .I(N__59856));
    InMux I__14050 (
            .O(N__59864),
            .I(N__59853));
    InMux I__14049 (
            .O(N__59863),
            .I(N__59850));
    InMux I__14048 (
            .O(N__59860),
            .I(N__59845));
    InMux I__14047 (
            .O(N__59859),
            .I(N__59845));
    Span4Mux_h I__14046 (
            .O(N__59856),
            .I(N__59842));
    LocalMux I__14045 (
            .O(N__59853),
            .I(r_Bit_Index_1));
    LocalMux I__14044 (
            .O(N__59850),
            .I(r_Bit_Index_1));
    LocalMux I__14043 (
            .O(N__59845),
            .I(r_Bit_Index_1));
    Odrv4 I__14042 (
            .O(N__59842),
            .I(r_Bit_Index_1));
    InMux I__14041 (
            .O(N__59833),
            .I(N__59829));
    CascadeMux I__14040 (
            .O(N__59832),
            .I(N__59826));
    LocalMux I__14039 (
            .O(N__59829),
            .I(N__59823));
    InMux I__14038 (
            .O(N__59826),
            .I(N__59820));
    Span4Mux_v I__14037 (
            .O(N__59823),
            .I(N__59817));
    LocalMux I__14036 (
            .O(N__59820),
            .I(N__59812));
    Span4Mux_v I__14035 (
            .O(N__59817),
            .I(N__59812));
    Span4Mux_v I__14034 (
            .O(N__59812),
            .I(N__59808));
    InMux I__14033 (
            .O(N__59811),
            .I(N__59805));
    Span4Mux_h I__14032 (
            .O(N__59808),
            .I(N__59802));
    LocalMux I__14031 (
            .O(N__59805),
            .I(data_in_frame_22_4));
    Odrv4 I__14030 (
            .O(N__59802),
            .I(data_in_frame_22_4));
    CascadeMux I__14029 (
            .O(N__59797),
            .I(N__59794));
    InMux I__14028 (
            .O(N__59794),
            .I(N__59791));
    LocalMux I__14027 (
            .O(N__59791),
            .I(N__59788));
    Span4Mux_h I__14026 (
            .O(N__59788),
            .I(N__59784));
    InMux I__14025 (
            .O(N__59787),
            .I(N__59781));
    Span4Mux_v I__14024 (
            .O(N__59784),
            .I(N__59778));
    LocalMux I__14023 (
            .O(N__59781),
            .I(N__59775));
    Odrv4 I__14022 (
            .O(N__59778),
            .I(\c0.n22191 ));
    Odrv12 I__14021 (
            .O(N__59775),
            .I(\c0.n22191 ));
    InMux I__14020 (
            .O(N__59770),
            .I(N__59767));
    LocalMux I__14019 (
            .O(N__59767),
            .I(N__59764));
    Span4Mux_h I__14018 (
            .O(N__59764),
            .I(N__59761));
    Odrv4 I__14017 (
            .O(N__59761),
            .I(\c0.n25 ));
    CascadeMux I__14016 (
            .O(N__59758),
            .I(N__59753));
    InMux I__14015 (
            .O(N__59757),
            .I(N__59740));
    InMux I__14014 (
            .O(N__59756),
            .I(N__59740));
    InMux I__14013 (
            .O(N__59753),
            .I(N__59740));
    InMux I__14012 (
            .O(N__59752),
            .I(N__59733));
    InMux I__14011 (
            .O(N__59751),
            .I(N__59733));
    InMux I__14010 (
            .O(N__59750),
            .I(N__59733));
    InMux I__14009 (
            .O(N__59749),
            .I(N__59728));
    InMux I__14008 (
            .O(N__59748),
            .I(N__59728));
    InMux I__14007 (
            .O(N__59747),
            .I(N__59725));
    LocalMux I__14006 (
            .O(N__59740),
            .I(r_Bit_Index_0));
    LocalMux I__14005 (
            .O(N__59733),
            .I(r_Bit_Index_0));
    LocalMux I__14004 (
            .O(N__59728),
            .I(r_Bit_Index_0));
    LocalMux I__14003 (
            .O(N__59725),
            .I(r_Bit_Index_0));
    CascadeMux I__14002 (
            .O(N__59716),
            .I(N__59712));
    CascadeMux I__14001 (
            .O(N__59715),
            .I(N__59705));
    InMux I__14000 (
            .O(N__59712),
            .I(N__59700));
    InMux I__13999 (
            .O(N__59711),
            .I(N__59700));
    CascadeMux I__13998 (
            .O(N__59710),
            .I(N__59695));
    CascadeMux I__13997 (
            .O(N__59709),
            .I(N__59691));
    InMux I__13996 (
            .O(N__59708),
            .I(N__59685));
    InMux I__13995 (
            .O(N__59705),
            .I(N__59685));
    LocalMux I__13994 (
            .O(N__59700),
            .I(N__59682));
    InMux I__13993 (
            .O(N__59699),
            .I(N__59677));
    InMux I__13992 (
            .O(N__59698),
            .I(N__59677));
    InMux I__13991 (
            .O(N__59695),
            .I(N__59672));
    InMux I__13990 (
            .O(N__59694),
            .I(N__59672));
    InMux I__13989 (
            .O(N__59691),
            .I(N__59669));
    CascadeMux I__13988 (
            .O(N__59690),
            .I(N__59666));
    LocalMux I__13987 (
            .O(N__59685),
            .I(N__59659));
    Span4Mux_h I__13986 (
            .O(N__59682),
            .I(N__59659));
    LocalMux I__13985 (
            .O(N__59677),
            .I(N__59659));
    LocalMux I__13984 (
            .O(N__59672),
            .I(N__59656));
    LocalMux I__13983 (
            .O(N__59669),
            .I(N__59650));
    InMux I__13982 (
            .O(N__59666),
            .I(N__59647));
    Span4Mux_h I__13981 (
            .O(N__59659),
            .I(N__59644));
    Span4Mux_v I__13980 (
            .O(N__59656),
            .I(N__59641));
    InMux I__13979 (
            .O(N__59655),
            .I(N__59634));
    InMux I__13978 (
            .O(N__59654),
            .I(N__59634));
    InMux I__13977 (
            .O(N__59653),
            .I(N__59634));
    Span4Mux_v I__13976 (
            .O(N__59650),
            .I(N__59631));
    LocalMux I__13975 (
            .O(N__59647),
            .I(N__59628));
    Span4Mux_v I__13974 (
            .O(N__59644),
            .I(N__59625));
    Sp12to4 I__13973 (
            .O(N__59641),
            .I(N__59620));
    LocalMux I__13972 (
            .O(N__59634),
            .I(N__59620));
    Span4Mux_v I__13971 (
            .O(N__59631),
            .I(N__59617));
    Span12Mux_h I__13970 (
            .O(N__59628),
            .I(N__59610));
    Sp12to4 I__13969 (
            .O(N__59625),
            .I(N__59610));
    Span12Mux_v I__13968 (
            .O(N__59620),
            .I(N__59610));
    Span4Mux_v I__13967 (
            .O(N__59617),
            .I(N__59607));
    Span12Mux_h I__13966 (
            .O(N__59610),
            .I(N__59604));
    Span4Mux_v I__13965 (
            .O(N__59607),
            .I(N__59601));
    Span12Mux_v I__13964 (
            .O(N__59604),
            .I(N__59598));
    Odrv4 I__13963 (
            .O(N__59601),
            .I(r_Rx_Data));
    Odrv12 I__13962 (
            .O(N__59598),
            .I(r_Rx_Data));
    CascadeMux I__13961 (
            .O(N__59593),
            .I(N__59589));
    InMux I__13960 (
            .O(N__59592),
            .I(N__59584));
    InMux I__13959 (
            .O(N__59589),
            .I(N__59584));
    LocalMux I__13958 (
            .O(N__59584),
            .I(n12970));
    InMux I__13957 (
            .O(N__59581),
            .I(N__59575));
    InMux I__13956 (
            .O(N__59580),
            .I(N__59572));
    InMux I__13955 (
            .O(N__59579),
            .I(N__59569));
    CascadeMux I__13954 (
            .O(N__59578),
            .I(N__59566));
    LocalMux I__13953 (
            .O(N__59575),
            .I(N__59563));
    LocalMux I__13952 (
            .O(N__59572),
            .I(N__59558));
    LocalMux I__13951 (
            .O(N__59569),
            .I(N__59558));
    InMux I__13950 (
            .O(N__59566),
            .I(N__59555));
    Span4Mux_h I__13949 (
            .O(N__59563),
            .I(N__59552));
    Span4Mux_h I__13948 (
            .O(N__59558),
            .I(N__59549));
    LocalMux I__13947 (
            .O(N__59555),
            .I(\c0.data_in_frame_12_0 ));
    Odrv4 I__13946 (
            .O(N__59552),
            .I(\c0.data_in_frame_12_0 ));
    Odrv4 I__13945 (
            .O(N__59549),
            .I(\c0.data_in_frame_12_0 ));
    InMux I__13944 (
            .O(N__59542),
            .I(N__59538));
    InMux I__13943 (
            .O(N__59541),
            .I(N__59535));
    LocalMux I__13942 (
            .O(N__59538),
            .I(N__59528));
    LocalMux I__13941 (
            .O(N__59535),
            .I(N__59528));
    InMux I__13940 (
            .O(N__59534),
            .I(N__59523));
    InMux I__13939 (
            .O(N__59533),
            .I(N__59523));
    Span4Mux_v I__13938 (
            .O(N__59528),
            .I(N__59517));
    LocalMux I__13937 (
            .O(N__59523),
            .I(N__59517));
    CascadeMux I__13936 (
            .O(N__59522),
            .I(N__59514));
    Span4Mux_v I__13935 (
            .O(N__59517),
            .I(N__59511));
    InMux I__13934 (
            .O(N__59514),
            .I(N__59508));
    Span4Mux_v I__13933 (
            .O(N__59511),
            .I(N__59505));
    LocalMux I__13932 (
            .O(N__59508),
            .I(\c0.data_in_frame_24_7 ));
    Odrv4 I__13931 (
            .O(N__59505),
            .I(\c0.data_in_frame_24_7 ));
    InMux I__13930 (
            .O(N__59500),
            .I(N__59496));
    CascadeMux I__13929 (
            .O(N__59499),
            .I(N__59493));
    LocalMux I__13928 (
            .O(N__59496),
            .I(N__59490));
    InMux I__13927 (
            .O(N__59493),
            .I(N__59485));
    Span4Mux_v I__13926 (
            .O(N__59490),
            .I(N__59482));
    InMux I__13925 (
            .O(N__59489),
            .I(N__59477));
    InMux I__13924 (
            .O(N__59488),
            .I(N__59477));
    LocalMux I__13923 (
            .O(N__59485),
            .I(\c0.data_in_frame_26_4 ));
    Odrv4 I__13922 (
            .O(N__59482),
            .I(\c0.data_in_frame_26_4 ));
    LocalMux I__13921 (
            .O(N__59477),
            .I(\c0.data_in_frame_26_4 ));
    InMux I__13920 (
            .O(N__59470),
            .I(N__59467));
    LocalMux I__13919 (
            .O(N__59467),
            .I(\c0.n22337 ));
    CascadeMux I__13918 (
            .O(N__59464),
            .I(\c0.n10_adj_4285_cascade_ ));
    InMux I__13917 (
            .O(N__59461),
            .I(N__59458));
    LocalMux I__13916 (
            .O(N__59458),
            .I(N__59455));
    Span4Mux_h I__13915 (
            .O(N__59455),
            .I(N__59452));
    Span4Mux_h I__13914 (
            .O(N__59452),
            .I(N__59449));
    Odrv4 I__13913 (
            .O(N__59449),
            .I(\c0.n22995 ));
    InMux I__13912 (
            .O(N__59446),
            .I(N__59440));
    InMux I__13911 (
            .O(N__59445),
            .I(N__59440));
    LocalMux I__13910 (
            .O(N__59440),
            .I(N__59436));
    CascadeMux I__13909 (
            .O(N__59439),
            .I(N__59433));
    Span4Mux_h I__13908 (
            .O(N__59436),
            .I(N__59430));
    InMux I__13907 (
            .O(N__59433),
            .I(N__59427));
    Span4Mux_v I__13906 (
            .O(N__59430),
            .I(N__59424));
    LocalMux I__13905 (
            .O(N__59427),
            .I(\c0.data_in_frame_26_6 ));
    Odrv4 I__13904 (
            .O(N__59424),
            .I(\c0.data_in_frame_26_6 ));
    InMux I__13903 (
            .O(N__59419),
            .I(N__59416));
    LocalMux I__13902 (
            .O(N__59416),
            .I(N__59413));
    Odrv4 I__13901 (
            .O(N__59413),
            .I(\c0.n22054 ));
    InMux I__13900 (
            .O(N__59410),
            .I(N__59402));
    InMux I__13899 (
            .O(N__59409),
            .I(N__59402));
    CascadeMux I__13898 (
            .O(N__59408),
            .I(N__59397));
    CascadeMux I__13897 (
            .O(N__59407),
            .I(N__59394));
    LocalMux I__13896 (
            .O(N__59402),
            .I(N__59390));
    InMux I__13895 (
            .O(N__59401),
            .I(N__59385));
    InMux I__13894 (
            .O(N__59400),
            .I(N__59385));
    InMux I__13893 (
            .O(N__59397),
            .I(N__59382));
    InMux I__13892 (
            .O(N__59394),
            .I(N__59377));
    InMux I__13891 (
            .O(N__59393),
            .I(N__59377));
    Span4Mux_v I__13890 (
            .O(N__59390),
            .I(N__59372));
    LocalMux I__13889 (
            .O(N__59385),
            .I(N__59372));
    LocalMux I__13888 (
            .O(N__59382),
            .I(\c0.data_in_frame_24_6 ));
    LocalMux I__13887 (
            .O(N__59377),
            .I(\c0.data_in_frame_24_6 ));
    Odrv4 I__13886 (
            .O(N__59372),
            .I(\c0.data_in_frame_24_6 ));
    CascadeMux I__13885 (
            .O(N__59365),
            .I(N__59362));
    InMux I__13884 (
            .O(N__59362),
            .I(N__59359));
    LocalMux I__13883 (
            .O(N__59359),
            .I(N__59356));
    Odrv12 I__13882 (
            .O(N__59356),
            .I(\c0.n22434 ));
    InMux I__13881 (
            .O(N__59353),
            .I(N__59349));
    InMux I__13880 (
            .O(N__59352),
            .I(N__59346));
    LocalMux I__13879 (
            .O(N__59349),
            .I(N__59343));
    LocalMux I__13878 (
            .O(N__59346),
            .I(N__59340));
    Span4Mux_v I__13877 (
            .O(N__59343),
            .I(N__59337));
    Span4Mux_v I__13876 (
            .O(N__59340),
            .I(N__59332));
    Sp12to4 I__13875 (
            .O(N__59337),
            .I(N__59329));
    InMux I__13874 (
            .O(N__59336),
            .I(N__59324));
    InMux I__13873 (
            .O(N__59335),
            .I(N__59324));
    Odrv4 I__13872 (
            .O(N__59332),
            .I(\c0.data_in_frame_20_0 ));
    Odrv12 I__13871 (
            .O(N__59329),
            .I(\c0.data_in_frame_20_0 ));
    LocalMux I__13870 (
            .O(N__59324),
            .I(\c0.data_in_frame_20_0 ));
    CascadeMux I__13869 (
            .O(N__59317),
            .I(N__59314));
    InMux I__13868 (
            .O(N__59314),
            .I(N__59311));
    LocalMux I__13867 (
            .O(N__59311),
            .I(N__59307));
    InMux I__13866 (
            .O(N__59310),
            .I(N__59303));
    Span12Mux_h I__13865 (
            .O(N__59307),
            .I(N__59300));
    InMux I__13864 (
            .O(N__59306),
            .I(N__59297));
    LocalMux I__13863 (
            .O(N__59303),
            .I(data_in_frame_22_2));
    Odrv12 I__13862 (
            .O(N__59300),
            .I(data_in_frame_22_2));
    LocalMux I__13861 (
            .O(N__59297),
            .I(data_in_frame_22_2));
    InMux I__13860 (
            .O(N__59290),
            .I(N__59286));
    InMux I__13859 (
            .O(N__59289),
            .I(N__59283));
    LocalMux I__13858 (
            .O(N__59286),
            .I(N__59280));
    LocalMux I__13857 (
            .O(N__59283),
            .I(N__59275));
    Span4Mux_v I__13856 (
            .O(N__59280),
            .I(N__59272));
    InMux I__13855 (
            .O(N__59279),
            .I(N__59269));
    InMux I__13854 (
            .O(N__59278),
            .I(N__59266));
    Odrv4 I__13853 (
            .O(N__59275),
            .I(\c0.n12594 ));
    Odrv4 I__13852 (
            .O(N__59272),
            .I(\c0.n12594 ));
    LocalMux I__13851 (
            .O(N__59269),
            .I(\c0.n12594 ));
    LocalMux I__13850 (
            .O(N__59266),
            .I(\c0.n12594 ));
    InMux I__13849 (
            .O(N__59257),
            .I(N__59253));
    InMux I__13848 (
            .O(N__59256),
            .I(N__59250));
    LocalMux I__13847 (
            .O(N__59253),
            .I(\c0.n20596 ));
    LocalMux I__13846 (
            .O(N__59250),
            .I(\c0.n20596 ));
    InMux I__13845 (
            .O(N__59245),
            .I(N__59241));
    InMux I__13844 (
            .O(N__59244),
            .I(N__59238));
    LocalMux I__13843 (
            .O(N__59241),
            .I(N__59235));
    LocalMux I__13842 (
            .O(N__59238),
            .I(N__59232));
    Span4Mux_v I__13841 (
            .O(N__59235),
            .I(N__59227));
    Span4Mux_h I__13840 (
            .O(N__59232),
            .I(N__59227));
    Span4Mux_v I__13839 (
            .O(N__59227),
            .I(N__59223));
    InMux I__13838 (
            .O(N__59226),
            .I(N__59220));
    Span4Mux_v I__13837 (
            .O(N__59223),
            .I(N__59217));
    LocalMux I__13836 (
            .O(N__59220),
            .I(\c0.data_in_frame_11_7 ));
    Odrv4 I__13835 (
            .O(N__59217),
            .I(\c0.data_in_frame_11_7 ));
    InMux I__13834 (
            .O(N__59212),
            .I(N__59207));
    InMux I__13833 (
            .O(N__59211),
            .I(N__59204));
    InMux I__13832 (
            .O(N__59210),
            .I(N__59201));
    LocalMux I__13831 (
            .O(N__59207),
            .I(N__59195));
    LocalMux I__13830 (
            .O(N__59204),
            .I(N__59190));
    LocalMux I__13829 (
            .O(N__59201),
            .I(N__59190));
    InMux I__13828 (
            .O(N__59200),
            .I(N__59187));
    InMux I__13827 (
            .O(N__59199),
            .I(N__59184));
    InMux I__13826 (
            .O(N__59198),
            .I(N__59181));
    Span4Mux_v I__13825 (
            .O(N__59195),
            .I(N__59178));
    Span4Mux_v I__13824 (
            .O(N__59190),
            .I(N__59173));
    LocalMux I__13823 (
            .O(N__59187),
            .I(N__59173));
    LocalMux I__13822 (
            .O(N__59184),
            .I(N__59170));
    LocalMux I__13821 (
            .O(N__59181),
            .I(N__59165));
    Span4Mux_v I__13820 (
            .O(N__59178),
            .I(N__59162));
    Span4Mux_v I__13819 (
            .O(N__59173),
            .I(N__59157));
    Span4Mux_v I__13818 (
            .O(N__59170),
            .I(N__59157));
    InMux I__13817 (
            .O(N__59169),
            .I(N__59154));
    InMux I__13816 (
            .O(N__59168),
            .I(N__59151));
    Span4Mux_v I__13815 (
            .O(N__59165),
            .I(N__59148));
    Sp12to4 I__13814 (
            .O(N__59162),
            .I(N__59141));
    Sp12to4 I__13813 (
            .O(N__59157),
            .I(N__59141));
    LocalMux I__13812 (
            .O(N__59154),
            .I(N__59141));
    LocalMux I__13811 (
            .O(N__59151),
            .I(N__59138));
    Sp12to4 I__13810 (
            .O(N__59148),
            .I(N__59135));
    Span12Mux_h I__13809 (
            .O(N__59141),
            .I(N__59130));
    Span12Mux_h I__13808 (
            .O(N__59138),
            .I(N__59130));
    Odrv12 I__13807 (
            .O(N__59135),
            .I(n21760));
    Odrv12 I__13806 (
            .O(N__59130),
            .I(n21760));
    CascadeMux I__13805 (
            .O(N__59125),
            .I(N__59122));
    InMux I__13804 (
            .O(N__59122),
            .I(N__59119));
    LocalMux I__13803 (
            .O(N__59119),
            .I(N__59114));
    InMux I__13802 (
            .O(N__59118),
            .I(N__59109));
    InMux I__13801 (
            .O(N__59117),
            .I(N__59109));
    Odrv12 I__13800 (
            .O(N__59114),
            .I(\c0.data_in_frame_26_2 ));
    LocalMux I__13799 (
            .O(N__59109),
            .I(\c0.data_in_frame_26_2 ));
    InMux I__13798 (
            .O(N__59104),
            .I(N__59101));
    LocalMux I__13797 (
            .O(N__59101),
            .I(N__59098));
    Odrv4 I__13796 (
            .O(N__59098),
            .I(\c0.n10_adj_4483 ));
    CascadeMux I__13795 (
            .O(N__59095),
            .I(\c0.n20537_cascade_ ));
    InMux I__13794 (
            .O(N__59092),
            .I(N__59089));
    LocalMux I__13793 (
            .O(N__59089),
            .I(N__59086));
    Span4Mux_v I__13792 (
            .O(N__59086),
            .I(N__59083));
    Odrv4 I__13791 (
            .O(N__59083),
            .I(\c0.n14_adj_4484 ));
    InMux I__13790 (
            .O(N__59080),
            .I(N__59074));
    InMux I__13789 (
            .O(N__59079),
            .I(N__59074));
    LocalMux I__13788 (
            .O(N__59074),
            .I(\c0.n21890 ));
    InMux I__13787 (
            .O(N__59071),
            .I(N__59068));
    LocalMux I__13786 (
            .O(N__59068),
            .I(N__59062));
    InMux I__13785 (
            .O(N__59067),
            .I(N__59059));
    InMux I__13784 (
            .O(N__59066),
            .I(N__59054));
    InMux I__13783 (
            .O(N__59065),
            .I(N__59054));
    Odrv4 I__13782 (
            .O(N__59062),
            .I(\c0.n21087 ));
    LocalMux I__13781 (
            .O(N__59059),
            .I(\c0.n21087 ));
    LocalMux I__13780 (
            .O(N__59054),
            .I(\c0.n21087 ));
    CascadeMux I__13779 (
            .O(N__59047),
            .I(\c0.n13320_cascade_ ));
    InMux I__13778 (
            .O(N__59044),
            .I(N__59038));
    InMux I__13777 (
            .O(N__59043),
            .I(N__59038));
    LocalMux I__13776 (
            .O(N__59038),
            .I(\c0.n22468 ));
    CascadeMux I__13775 (
            .O(N__59035),
            .I(\c0.n10_cascade_ ));
    InMux I__13774 (
            .O(N__59032),
            .I(N__59026));
    InMux I__13773 (
            .O(N__59031),
            .I(N__59026));
    LocalMux I__13772 (
            .O(N__59026),
            .I(\c0.n20537 ));
    InMux I__13771 (
            .O(N__59023),
            .I(N__59020));
    LocalMux I__13770 (
            .O(N__59020),
            .I(N__59016));
    InMux I__13769 (
            .O(N__59019),
            .I(N__59013));
    Odrv4 I__13768 (
            .O(N__59016),
            .I(\c0.n22314 ));
    LocalMux I__13767 (
            .O(N__59013),
            .I(\c0.n22314 ));
    InMux I__13766 (
            .O(N__59008),
            .I(N__59003));
    InMux I__13765 (
            .O(N__59007),
            .I(N__59000));
    CascadeMux I__13764 (
            .O(N__59006),
            .I(N__58997));
    LocalMux I__13763 (
            .O(N__59003),
            .I(N__58993));
    LocalMux I__13762 (
            .O(N__59000),
            .I(N__58990));
    InMux I__13761 (
            .O(N__58997),
            .I(N__58987));
    InMux I__13760 (
            .O(N__58996),
            .I(N__58984));
    Span4Mux_v I__13759 (
            .O(N__58993),
            .I(N__58979));
    Span4Mux_v I__13758 (
            .O(N__58990),
            .I(N__58979));
    LocalMux I__13757 (
            .O(N__58987),
            .I(\c0.data_in_frame_24_3 ));
    LocalMux I__13756 (
            .O(N__58984),
            .I(\c0.data_in_frame_24_3 ));
    Odrv4 I__13755 (
            .O(N__58979),
            .I(\c0.data_in_frame_24_3 ));
    InMux I__13754 (
            .O(N__58972),
            .I(N__58969));
    LocalMux I__13753 (
            .O(N__58969),
            .I(N__58966));
    Span4Mux_v I__13752 (
            .O(N__58966),
            .I(N__58963));
    Odrv4 I__13751 (
            .O(N__58963),
            .I(\c0.n22142 ));
    InMux I__13750 (
            .O(N__58960),
            .I(N__58957));
    LocalMux I__13749 (
            .O(N__58957),
            .I(N__58954));
    Span4Mux_v I__13748 (
            .O(N__58954),
            .I(N__58949));
    InMux I__13747 (
            .O(N__58953),
            .I(N__58944));
    InMux I__13746 (
            .O(N__58952),
            .I(N__58944));
    Span4Mux_h I__13745 (
            .O(N__58949),
            .I(N__58939));
    LocalMux I__13744 (
            .O(N__58944),
            .I(N__58939));
    Span4Mux_v I__13743 (
            .O(N__58939),
            .I(N__58935));
    CascadeMux I__13742 (
            .O(N__58938),
            .I(N__58932));
    Span4Mux_h I__13741 (
            .O(N__58935),
            .I(N__58929));
    InMux I__13740 (
            .O(N__58932),
            .I(N__58926));
    Span4Mux_h I__13739 (
            .O(N__58929),
            .I(N__58923));
    LocalMux I__13738 (
            .O(N__58926),
            .I(\c0.data_in_frame_24_4 ));
    Odrv4 I__13737 (
            .O(N__58923),
            .I(\c0.data_in_frame_24_4 ));
    InMux I__13736 (
            .O(N__58918),
            .I(N__58915));
    LocalMux I__13735 (
            .O(N__58915),
            .I(N__58912));
    Span4Mux_h I__13734 (
            .O(N__58912),
            .I(N__58909));
    Odrv4 I__13733 (
            .O(N__58909),
            .I(\c0.n22028 ));
    CascadeMux I__13732 (
            .O(N__58906),
            .I(\c0.n22337_cascade_ ));
    InMux I__13731 (
            .O(N__58903),
            .I(N__58900));
    LocalMux I__13730 (
            .O(N__58900),
            .I(N__58893));
    InMux I__13729 (
            .O(N__58899),
            .I(N__58890));
    InMux I__13728 (
            .O(N__58898),
            .I(N__58885));
    InMux I__13727 (
            .O(N__58897),
            .I(N__58885));
    InMux I__13726 (
            .O(N__58896),
            .I(N__58882));
    Span4Mux_h I__13725 (
            .O(N__58893),
            .I(N__58873));
    LocalMux I__13724 (
            .O(N__58890),
            .I(N__58873));
    LocalMux I__13723 (
            .O(N__58885),
            .I(N__58873));
    LocalMux I__13722 (
            .O(N__58882),
            .I(N__58873));
    Span4Mux_v I__13721 (
            .O(N__58873),
            .I(N__58870));
    Odrv4 I__13720 (
            .O(N__58870),
            .I(\c0.n22020 ));
    InMux I__13719 (
            .O(N__58867),
            .I(N__58861));
    InMux I__13718 (
            .O(N__58866),
            .I(N__58861));
    LocalMux I__13717 (
            .O(N__58861),
            .I(N__58858));
    Span12Mux_v I__13716 (
            .O(N__58858),
            .I(N__58855));
    Odrv12 I__13715 (
            .O(N__58855),
            .I(\c0.n21095 ));
    InMux I__13714 (
            .O(N__58852),
            .I(N__58849));
    LocalMux I__13713 (
            .O(N__58849),
            .I(\c0.n6_adj_4418 ));
    CascadeMux I__13712 (
            .O(N__58846),
            .I(N__58842));
    CascadeMux I__13711 (
            .O(N__58845),
            .I(N__58839));
    InMux I__13710 (
            .O(N__58842),
            .I(N__58832));
    InMux I__13709 (
            .O(N__58839),
            .I(N__58829));
    InMux I__13708 (
            .O(N__58838),
            .I(N__58826));
    InMux I__13707 (
            .O(N__58837),
            .I(N__58823));
    CascadeMux I__13706 (
            .O(N__58836),
            .I(N__58819));
    CascadeMux I__13705 (
            .O(N__58835),
            .I(N__58816));
    LocalMux I__13704 (
            .O(N__58832),
            .I(N__58813));
    LocalMux I__13703 (
            .O(N__58829),
            .I(N__58810));
    LocalMux I__13702 (
            .O(N__58826),
            .I(N__58807));
    LocalMux I__13701 (
            .O(N__58823),
            .I(N__58804));
    InMux I__13700 (
            .O(N__58822),
            .I(N__58799));
    InMux I__13699 (
            .O(N__58819),
            .I(N__58799));
    InMux I__13698 (
            .O(N__58816),
            .I(N__58796));
    Span4Mux_h I__13697 (
            .O(N__58813),
            .I(N__58793));
    Span4Mux_h I__13696 (
            .O(N__58810),
            .I(N__58788));
    Span4Mux_v I__13695 (
            .O(N__58807),
            .I(N__58788));
    Span4Mux_v I__13694 (
            .O(N__58804),
            .I(N__58783));
    LocalMux I__13693 (
            .O(N__58799),
            .I(N__58783));
    LocalMux I__13692 (
            .O(N__58796),
            .I(\c0.data_in_frame_19_5 ));
    Odrv4 I__13691 (
            .O(N__58793),
            .I(\c0.data_in_frame_19_5 ));
    Odrv4 I__13690 (
            .O(N__58788),
            .I(\c0.data_in_frame_19_5 ));
    Odrv4 I__13689 (
            .O(N__58783),
            .I(\c0.data_in_frame_19_5 ));
    InMux I__13688 (
            .O(N__58774),
            .I(N__58771));
    LocalMux I__13687 (
            .O(N__58771),
            .I(N__58767));
    InMux I__13686 (
            .O(N__58770),
            .I(N__58763));
    Span4Mux_h I__13685 (
            .O(N__58767),
            .I(N__58760));
    InMux I__13684 (
            .O(N__58766),
            .I(N__58757));
    LocalMux I__13683 (
            .O(N__58763),
            .I(N__58754));
    Span4Mux_h I__13682 (
            .O(N__58760),
            .I(N__58751));
    LocalMux I__13681 (
            .O(N__58757),
            .I(N__58746));
    Span4Mux_v I__13680 (
            .O(N__58754),
            .I(N__58746));
    Odrv4 I__13679 (
            .O(N__58751),
            .I(\c0.data_in_frame_26_1 ));
    Odrv4 I__13678 (
            .O(N__58746),
            .I(\c0.data_in_frame_26_1 ));
    InMux I__13677 (
            .O(N__58741),
            .I(N__58737));
    InMux I__13676 (
            .O(N__58740),
            .I(N__58734));
    LocalMux I__13675 (
            .O(N__58737),
            .I(\c0.n21039 ));
    LocalMux I__13674 (
            .O(N__58734),
            .I(\c0.n21039 ));
    CascadeMux I__13673 (
            .O(N__58729),
            .I(\c0.n24_adj_4282_cascade_ ));
    InMux I__13672 (
            .O(N__58726),
            .I(N__58723));
    LocalMux I__13671 (
            .O(N__58723),
            .I(\c0.n22711 ));
    CascadeMux I__13670 (
            .O(N__58720),
            .I(\c0.n22711_cascade_ ));
    InMux I__13669 (
            .O(N__58717),
            .I(N__58714));
    LocalMux I__13668 (
            .O(N__58714),
            .I(N__58709));
    InMux I__13667 (
            .O(N__58713),
            .I(N__58706));
    InMux I__13666 (
            .O(N__58712),
            .I(N__58703));
    Odrv4 I__13665 (
            .O(N__58709),
            .I(\c0.n21200 ));
    LocalMux I__13664 (
            .O(N__58706),
            .I(\c0.n21200 ));
    LocalMux I__13663 (
            .O(N__58703),
            .I(\c0.n21200 ));
    InMux I__13662 (
            .O(N__58696),
            .I(N__58693));
    LocalMux I__13661 (
            .O(N__58693),
            .I(N__58688));
    InMux I__13660 (
            .O(N__58692),
            .I(N__58685));
    InMux I__13659 (
            .O(N__58691),
            .I(N__58682));
    Odrv4 I__13658 (
            .O(N__58688),
            .I(\c0.n12596 ));
    LocalMux I__13657 (
            .O(N__58685),
            .I(\c0.n12596 ));
    LocalMux I__13656 (
            .O(N__58682),
            .I(\c0.n12596 ));
    CascadeMux I__13655 (
            .O(N__58675),
            .I(N__58672));
    InMux I__13654 (
            .O(N__58672),
            .I(N__58669));
    LocalMux I__13653 (
            .O(N__58669),
            .I(N__58666));
    Span12Mux_s10_h I__13652 (
            .O(N__58666),
            .I(N__58663));
    Odrv12 I__13651 (
            .O(N__58663),
            .I(\c0.n6707 ));
    CascadeMux I__13650 (
            .O(N__58660),
            .I(\c0.n15_adj_4284_cascade_ ));
    InMux I__13649 (
            .O(N__58657),
            .I(N__58654));
    LocalMux I__13648 (
            .O(N__58654),
            .I(\c0.n14_adj_4283 ));
    InMux I__13647 (
            .O(N__58651),
            .I(N__58648));
    LocalMux I__13646 (
            .O(N__58648),
            .I(\c0.n22437 ));
    InMux I__13645 (
            .O(N__58645),
            .I(N__58638));
    InMux I__13644 (
            .O(N__58644),
            .I(N__58638));
    InMux I__13643 (
            .O(N__58643),
            .I(N__58634));
    LocalMux I__13642 (
            .O(N__58638),
            .I(N__58631));
    InMux I__13641 (
            .O(N__58637),
            .I(N__58628));
    LocalMux I__13640 (
            .O(N__58634),
            .I(N__58623));
    Sp12to4 I__13639 (
            .O(N__58631),
            .I(N__58623));
    LocalMux I__13638 (
            .O(N__58628),
            .I(\c0.data_in_frame_25_0 ));
    Odrv12 I__13637 (
            .O(N__58623),
            .I(\c0.data_in_frame_25_0 ));
    InMux I__13636 (
            .O(N__58618),
            .I(N__58615));
    LocalMux I__13635 (
            .O(N__58615),
            .I(N__58611));
    InMux I__13634 (
            .O(N__58614),
            .I(N__58606));
    Span4Mux_v I__13633 (
            .O(N__58611),
            .I(N__58603));
    CascadeMux I__13632 (
            .O(N__58610),
            .I(N__58600));
    InMux I__13631 (
            .O(N__58609),
            .I(N__58597));
    LocalMux I__13630 (
            .O(N__58606),
            .I(N__58594));
    Span4Mux_h I__13629 (
            .O(N__58603),
            .I(N__58591));
    InMux I__13628 (
            .O(N__58600),
            .I(N__58588));
    LocalMux I__13627 (
            .O(N__58597),
            .I(N__58583));
    Span4Mux_v I__13626 (
            .O(N__58594),
            .I(N__58583));
    Span4Mux_v I__13625 (
            .O(N__58591),
            .I(N__58580));
    LocalMux I__13624 (
            .O(N__58588),
            .I(\c0.data_in_frame_25_6 ));
    Odrv4 I__13623 (
            .O(N__58583),
            .I(\c0.data_in_frame_25_6 ));
    Odrv4 I__13622 (
            .O(N__58580),
            .I(\c0.data_in_frame_25_6 ));
    CascadeMux I__13621 (
            .O(N__58573),
            .I(\c0.n22437_cascade_ ));
    CascadeMux I__13620 (
            .O(N__58570),
            .I(N__58567));
    InMux I__13619 (
            .O(N__58567),
            .I(N__58564));
    LocalMux I__13618 (
            .O(N__58564),
            .I(\c0.n50_adj_4487 ));
    InMux I__13617 (
            .O(N__58561),
            .I(N__58557));
    InMux I__13616 (
            .O(N__58560),
            .I(N__58554));
    LocalMux I__13615 (
            .O(N__58557),
            .I(N__58551));
    LocalMux I__13614 (
            .O(N__58554),
            .I(N__58548));
    Odrv12 I__13613 (
            .O(N__58551),
            .I(\c0.n22323 ));
    Odrv4 I__13612 (
            .O(N__58548),
            .I(\c0.n22323 ));
    InMux I__13611 (
            .O(N__58543),
            .I(N__58536));
    InMux I__13610 (
            .O(N__58542),
            .I(N__58536));
    InMux I__13609 (
            .O(N__58541),
            .I(N__58533));
    LocalMux I__13608 (
            .O(N__58536),
            .I(\c0.n20203 ));
    LocalMux I__13607 (
            .O(N__58533),
            .I(\c0.n20203 ));
    InMux I__13606 (
            .O(N__58528),
            .I(N__58525));
    LocalMux I__13605 (
            .O(N__58525),
            .I(N__58522));
    Span4Mux_v I__13604 (
            .O(N__58522),
            .I(N__58519));
    Odrv4 I__13603 (
            .O(N__58519),
            .I(\c0.n21870 ));
    CascadeMux I__13602 (
            .O(N__58516),
            .I(\c0.n18_adj_4249_cascade_ ));
    InMux I__13601 (
            .O(N__58513),
            .I(N__58510));
    LocalMux I__13600 (
            .O(N__58510),
            .I(N__58507));
    Odrv4 I__13599 (
            .O(N__58507),
            .I(\c0.n24_adj_4248 ));
    InMux I__13598 (
            .O(N__58504),
            .I(N__58501));
    LocalMux I__13597 (
            .O(N__58501),
            .I(\c0.n26_adj_4250 ));
    CascadeMux I__13596 (
            .O(N__58498),
            .I(N__58494));
    InMux I__13595 (
            .O(N__58497),
            .I(N__58491));
    InMux I__13594 (
            .O(N__58494),
            .I(N__58487));
    LocalMux I__13593 (
            .O(N__58491),
            .I(N__58484));
    InMux I__13592 (
            .O(N__58490),
            .I(N__58480));
    LocalMux I__13591 (
            .O(N__58487),
            .I(N__58475));
    Span4Mux_h I__13590 (
            .O(N__58484),
            .I(N__58475));
    InMux I__13589 (
            .O(N__58483),
            .I(N__58472));
    LocalMux I__13588 (
            .O(N__58480),
            .I(N__58469));
    Span4Mux_v I__13587 (
            .O(N__58475),
            .I(N__58466));
    LocalMux I__13586 (
            .O(N__58472),
            .I(\c0.data_in_frame_15_4 ));
    Odrv4 I__13585 (
            .O(N__58469),
            .I(\c0.data_in_frame_15_4 ));
    Odrv4 I__13584 (
            .O(N__58466),
            .I(\c0.data_in_frame_15_4 ));
    InMux I__13583 (
            .O(N__58459),
            .I(N__58455));
    InMux I__13582 (
            .O(N__58458),
            .I(N__58452));
    LocalMux I__13581 (
            .O(N__58455),
            .I(\c0.n23072 ));
    LocalMux I__13580 (
            .O(N__58452),
            .I(\c0.n23072 ));
    InMux I__13579 (
            .O(N__58447),
            .I(N__58441));
    InMux I__13578 (
            .O(N__58446),
            .I(N__58441));
    LocalMux I__13577 (
            .O(N__58441),
            .I(N__58438));
    Span4Mux_h I__13576 (
            .O(N__58438),
            .I(N__58435));
    Odrv4 I__13575 (
            .O(N__58435),
            .I(\c0.n13457 ));
    CascadeMux I__13574 (
            .O(N__58432),
            .I(\c0.n23072_cascade_ ));
    InMux I__13573 (
            .O(N__58429),
            .I(N__58423));
    InMux I__13572 (
            .O(N__58428),
            .I(N__58420));
    InMux I__13571 (
            .O(N__58427),
            .I(N__58417));
    InMux I__13570 (
            .O(N__58426),
            .I(N__58414));
    LocalMux I__13569 (
            .O(N__58423),
            .I(N__58409));
    LocalMux I__13568 (
            .O(N__58420),
            .I(N__58409));
    LocalMux I__13567 (
            .O(N__58417),
            .I(N__58404));
    LocalMux I__13566 (
            .O(N__58414),
            .I(N__58404));
    Span4Mux_v I__13565 (
            .O(N__58409),
            .I(N__58401));
    Odrv12 I__13564 (
            .O(N__58404),
            .I(\c0.n21067 ));
    Odrv4 I__13563 (
            .O(N__58401),
            .I(\c0.n21067 ));
    InMux I__13562 (
            .O(N__58396),
            .I(N__58393));
    LocalMux I__13561 (
            .O(N__58393),
            .I(\c0.n14_adj_4251 ));
    InMux I__13560 (
            .O(N__58390),
            .I(N__58387));
    LocalMux I__13559 (
            .O(N__58387),
            .I(\c0.n21054 ));
    CascadeMux I__13558 (
            .O(N__58384),
            .I(\c0.n6_adj_4292_cascade_ ));
    InMux I__13557 (
            .O(N__58381),
            .I(N__58378));
    LocalMux I__13556 (
            .O(N__58378),
            .I(N__58374));
    CascadeMux I__13555 (
            .O(N__58377),
            .I(N__58371));
    Span4Mux_v I__13554 (
            .O(N__58374),
            .I(N__58368));
    InMux I__13553 (
            .O(N__58371),
            .I(N__58365));
    Span4Mux_h I__13552 (
            .O(N__58368),
            .I(N__58362));
    LocalMux I__13551 (
            .O(N__58365),
            .I(\c0.data_in_frame_28_5 ));
    Odrv4 I__13550 (
            .O(N__58362),
            .I(\c0.data_in_frame_28_5 ));
    InMux I__13549 (
            .O(N__58357),
            .I(N__58354));
    LocalMux I__13548 (
            .O(N__58354),
            .I(N__58351));
    Span4Mux_v I__13547 (
            .O(N__58351),
            .I(N__58348));
    Span4Mux_h I__13546 (
            .O(N__58348),
            .I(N__58345));
    Odrv4 I__13545 (
            .O(N__58345),
            .I(\c0.n23073 ));
    InMux I__13544 (
            .O(N__58342),
            .I(N__58338));
    InMux I__13543 (
            .O(N__58341),
            .I(N__58334));
    LocalMux I__13542 (
            .O(N__58338),
            .I(N__58331));
    CascadeMux I__13541 (
            .O(N__58337),
            .I(N__58328));
    LocalMux I__13540 (
            .O(N__58334),
            .I(N__58324));
    Span4Mux_h I__13539 (
            .O(N__58331),
            .I(N__58321));
    InMux I__13538 (
            .O(N__58328),
            .I(N__58318));
    InMux I__13537 (
            .O(N__58327),
            .I(N__58315));
    Span4Mux_h I__13536 (
            .O(N__58324),
            .I(N__58312));
    Span4Mux_v I__13535 (
            .O(N__58321),
            .I(N__58309));
    LocalMux I__13534 (
            .O(N__58318),
            .I(\c0.data_in_frame_21_4 ));
    LocalMux I__13533 (
            .O(N__58315),
            .I(\c0.data_in_frame_21_4 ));
    Odrv4 I__13532 (
            .O(N__58312),
            .I(\c0.data_in_frame_21_4 ));
    Odrv4 I__13531 (
            .O(N__58309),
            .I(\c0.data_in_frame_21_4 ));
    InMux I__13530 (
            .O(N__58300),
            .I(N__58297));
    LocalMux I__13529 (
            .O(N__58297),
            .I(\c0.n21905 ));
    CascadeMux I__13528 (
            .O(N__58294),
            .I(\c0.n21905_cascade_ ));
    InMux I__13527 (
            .O(N__58291),
            .I(N__58288));
    LocalMux I__13526 (
            .O(N__58288),
            .I(N__58285));
    Span12Mux_v I__13525 (
            .O(N__58285),
            .I(N__58282));
    Odrv12 I__13524 (
            .O(N__58282),
            .I(\c0.n21069 ));
    InMux I__13523 (
            .O(N__58279),
            .I(N__58275));
    InMux I__13522 (
            .O(N__58278),
            .I(N__58272));
    LocalMux I__13521 (
            .O(N__58275),
            .I(N__58269));
    LocalMux I__13520 (
            .O(N__58272),
            .I(N__58266));
    Odrv4 I__13519 (
            .O(N__58269),
            .I(\c0.n22113 ));
    Odrv4 I__13518 (
            .O(N__58266),
            .I(\c0.n22113 ));
    CascadeMux I__13517 (
            .O(N__58261),
            .I(N__58258));
    InMux I__13516 (
            .O(N__58258),
            .I(N__58253));
    InMux I__13515 (
            .O(N__58257),
            .I(N__58248));
    InMux I__13514 (
            .O(N__58256),
            .I(N__58248));
    LocalMux I__13513 (
            .O(N__58253),
            .I(\c0.data_in_frame_20_3 ));
    LocalMux I__13512 (
            .O(N__58248),
            .I(\c0.data_in_frame_20_3 ));
    InMux I__13511 (
            .O(N__58243),
            .I(N__58240));
    LocalMux I__13510 (
            .O(N__58240),
            .I(\c0.n22352 ));
    CascadeMux I__13509 (
            .O(N__58237),
            .I(N__58233));
    CascadeMux I__13508 (
            .O(N__58236),
            .I(N__58230));
    InMux I__13507 (
            .O(N__58233),
            .I(N__58227));
    InMux I__13506 (
            .O(N__58230),
            .I(N__58224));
    LocalMux I__13505 (
            .O(N__58227),
            .I(N__58221));
    LocalMux I__13504 (
            .O(N__58224),
            .I(\c0.data_in_frame_18_4 ));
    Odrv4 I__13503 (
            .O(N__58221),
            .I(\c0.data_in_frame_18_4 ));
    InMux I__13502 (
            .O(N__58216),
            .I(N__58213));
    LocalMux I__13501 (
            .O(N__58213),
            .I(N__58209));
    InMux I__13500 (
            .O(N__58212),
            .I(N__58206));
    Span4Mux_h I__13499 (
            .O(N__58209),
            .I(N__58200));
    LocalMux I__13498 (
            .O(N__58206),
            .I(N__58200));
    InMux I__13497 (
            .O(N__58205),
            .I(N__58197));
    Span4Mux_v I__13496 (
            .O(N__58200),
            .I(N__58194));
    LocalMux I__13495 (
            .O(N__58197),
            .I(\c0.n13598 ));
    Odrv4 I__13494 (
            .O(N__58194),
            .I(\c0.n13598 ));
    InMux I__13493 (
            .O(N__58189),
            .I(N__58186));
    LocalMux I__13492 (
            .O(N__58186),
            .I(N__58182));
    InMux I__13491 (
            .O(N__58185),
            .I(N__58179));
    Odrv12 I__13490 (
            .O(N__58182),
            .I(\c0.n20374 ));
    LocalMux I__13489 (
            .O(N__58179),
            .I(\c0.n20374 ));
    CascadeMux I__13488 (
            .O(N__58174),
            .I(N__58169));
    CascadeMux I__13487 (
            .O(N__58173),
            .I(N__58166));
    InMux I__13486 (
            .O(N__58172),
            .I(N__58163));
    InMux I__13485 (
            .O(N__58169),
            .I(N__58159));
    InMux I__13484 (
            .O(N__58166),
            .I(N__58156));
    LocalMux I__13483 (
            .O(N__58163),
            .I(N__58153));
    InMux I__13482 (
            .O(N__58162),
            .I(N__58150));
    LocalMux I__13481 (
            .O(N__58159),
            .I(\c0.data_in_frame_16_5 ));
    LocalMux I__13480 (
            .O(N__58156),
            .I(\c0.data_in_frame_16_5 ));
    Odrv4 I__13479 (
            .O(N__58153),
            .I(\c0.data_in_frame_16_5 ));
    LocalMux I__13478 (
            .O(N__58150),
            .I(\c0.data_in_frame_16_5 ));
    InMux I__13477 (
            .O(N__58141),
            .I(N__58138));
    LocalMux I__13476 (
            .O(N__58138),
            .I(N__58134));
    InMux I__13475 (
            .O(N__58137),
            .I(N__58131));
    Span4Mux_v I__13474 (
            .O(N__58134),
            .I(N__58127));
    LocalMux I__13473 (
            .O(N__58131),
            .I(N__58124));
    CascadeMux I__13472 (
            .O(N__58130),
            .I(N__58121));
    Span4Mux_v I__13471 (
            .O(N__58127),
            .I(N__58118));
    Span4Mux_h I__13470 (
            .O(N__58124),
            .I(N__58115));
    InMux I__13469 (
            .O(N__58121),
            .I(N__58112));
    Span4Mux_h I__13468 (
            .O(N__58118),
            .I(N__58109));
    Span4Mux_h I__13467 (
            .O(N__58115),
            .I(N__58106));
    LocalMux I__13466 (
            .O(N__58112),
            .I(\c0.data_in_frame_16_3 ));
    Odrv4 I__13465 (
            .O(N__58109),
            .I(\c0.data_in_frame_16_3 ));
    Odrv4 I__13464 (
            .O(N__58106),
            .I(\c0.data_in_frame_16_3 ));
    CascadeMux I__13463 (
            .O(N__58099),
            .I(N__58095));
    InMux I__13462 (
            .O(N__58098),
            .I(N__58091));
    InMux I__13461 (
            .O(N__58095),
            .I(N__58088));
    InMux I__13460 (
            .O(N__58094),
            .I(N__58085));
    LocalMux I__13459 (
            .O(N__58091),
            .I(N__58082));
    LocalMux I__13458 (
            .O(N__58088),
            .I(\c0.data_in_frame_16_2 ));
    LocalMux I__13457 (
            .O(N__58085),
            .I(\c0.data_in_frame_16_2 ));
    Odrv4 I__13456 (
            .O(N__58082),
            .I(\c0.data_in_frame_16_2 ));
    InMux I__13455 (
            .O(N__58075),
            .I(N__58072));
    LocalMux I__13454 (
            .O(N__58072),
            .I(\c0.n10_adj_4230 ));
    CascadeMux I__13453 (
            .O(N__58069),
            .I(N__58064));
    InMux I__13452 (
            .O(N__58068),
            .I(N__58056));
    InMux I__13451 (
            .O(N__58067),
            .I(N__58056));
    InMux I__13450 (
            .O(N__58064),
            .I(N__58051));
    InMux I__13449 (
            .O(N__58063),
            .I(N__58051));
    InMux I__13448 (
            .O(N__58062),
            .I(N__58046));
    InMux I__13447 (
            .O(N__58061),
            .I(N__58046));
    LocalMux I__13446 (
            .O(N__58056),
            .I(N__58043));
    LocalMux I__13445 (
            .O(N__58051),
            .I(\c0.data_in_frame_13_4 ));
    LocalMux I__13444 (
            .O(N__58046),
            .I(\c0.data_in_frame_13_4 ));
    Odrv12 I__13443 (
            .O(N__58043),
            .I(\c0.data_in_frame_13_4 ));
    CascadeMux I__13442 (
            .O(N__58036),
            .I(N__58033));
    InMux I__13441 (
            .O(N__58033),
            .I(N__58030));
    LocalMux I__13440 (
            .O(N__58030),
            .I(N__58025));
    InMux I__13439 (
            .O(N__58029),
            .I(N__58022));
    CascadeMux I__13438 (
            .O(N__58028),
            .I(N__58019));
    Span4Mux_v I__13437 (
            .O(N__58025),
            .I(N__58013));
    LocalMux I__13436 (
            .O(N__58022),
            .I(N__58013));
    InMux I__13435 (
            .O(N__58019),
            .I(N__58010));
    InMux I__13434 (
            .O(N__58018),
            .I(N__58007));
    Span4Mux_h I__13433 (
            .O(N__58013),
            .I(N__58004));
    LocalMux I__13432 (
            .O(N__58010),
            .I(\c0.data_in_frame_15_5 ));
    LocalMux I__13431 (
            .O(N__58007),
            .I(\c0.data_in_frame_15_5 ));
    Odrv4 I__13430 (
            .O(N__58004),
            .I(\c0.data_in_frame_15_5 ));
    CascadeMux I__13429 (
            .O(N__57997),
            .I(N__57994));
    InMux I__13428 (
            .O(N__57994),
            .I(N__57991));
    LocalMux I__13427 (
            .O(N__57991),
            .I(N__57988));
    Span4Mux_v I__13426 (
            .O(N__57988),
            .I(N__57984));
    InMux I__13425 (
            .O(N__57987),
            .I(N__57981));
    Span4Mux_h I__13424 (
            .O(N__57984),
            .I(N__57978));
    LocalMux I__13423 (
            .O(N__57981),
            .I(\c0.data_in_frame_26_3 ));
    Odrv4 I__13422 (
            .O(N__57978),
            .I(\c0.data_in_frame_26_3 ));
    InMux I__13421 (
            .O(N__57973),
            .I(N__57969));
    CascadeMux I__13420 (
            .O(N__57972),
            .I(N__57966));
    LocalMux I__13419 (
            .O(N__57969),
            .I(N__57963));
    InMux I__13418 (
            .O(N__57966),
            .I(N__57960));
    Odrv4 I__13417 (
            .O(N__57963),
            .I(\c0.n20266 ));
    LocalMux I__13416 (
            .O(N__57960),
            .I(\c0.n20266 ));
    CascadeMux I__13415 (
            .O(N__57955),
            .I(\c0.n22402_cascade_ ));
    InMux I__13414 (
            .O(N__57952),
            .I(N__57949));
    LocalMux I__13413 (
            .O(N__57949),
            .I(N__57946));
    Span4Mux_v I__13412 (
            .O(N__57946),
            .I(N__57943));
    Odrv4 I__13411 (
            .O(N__57943),
            .I(\c0.n33 ));
    InMux I__13410 (
            .O(N__57940),
            .I(N__57937));
    LocalMux I__13409 (
            .O(N__57937),
            .I(N__57933));
    InMux I__13408 (
            .O(N__57936),
            .I(N__57930));
    Odrv4 I__13407 (
            .O(N__57933),
            .I(\c0.n21982 ));
    LocalMux I__13406 (
            .O(N__57930),
            .I(\c0.n21982 ));
    InMux I__13405 (
            .O(N__57925),
            .I(N__57921));
    InMux I__13404 (
            .O(N__57924),
            .I(N__57918));
    LocalMux I__13403 (
            .O(N__57921),
            .I(N__57915));
    LocalMux I__13402 (
            .O(N__57918),
            .I(data_in_frame_14_0));
    Odrv12 I__13401 (
            .O(N__57915),
            .I(data_in_frame_14_0));
    InMux I__13400 (
            .O(N__57910),
            .I(N__57905));
    InMux I__13399 (
            .O(N__57909),
            .I(N__57902));
    InMux I__13398 (
            .O(N__57908),
            .I(N__57899));
    LocalMux I__13397 (
            .O(N__57905),
            .I(N__57896));
    LocalMux I__13396 (
            .O(N__57902),
            .I(N__57893));
    LocalMux I__13395 (
            .O(N__57899),
            .I(N__57890));
    Span4Mux_h I__13394 (
            .O(N__57896),
            .I(N__57882));
    Span4Mux_v I__13393 (
            .O(N__57893),
            .I(N__57882));
    Span4Mux_v I__13392 (
            .O(N__57890),
            .I(N__57882));
    InMux I__13391 (
            .O(N__57889),
            .I(N__57879));
    Odrv4 I__13390 (
            .O(N__57882),
            .I(\c0.n13865 ));
    LocalMux I__13389 (
            .O(N__57879),
            .I(\c0.n13865 ));
    InMux I__13388 (
            .O(N__57874),
            .I(N__57871));
    LocalMux I__13387 (
            .O(N__57871),
            .I(N__57866));
    InMux I__13386 (
            .O(N__57870),
            .I(N__57863));
    InMux I__13385 (
            .O(N__57869),
            .I(N__57860));
    Span4Mux_v I__13384 (
            .O(N__57866),
            .I(N__57857));
    LocalMux I__13383 (
            .O(N__57863),
            .I(\c0.data_in_frame_15_6 ));
    LocalMux I__13382 (
            .O(N__57860),
            .I(\c0.data_in_frame_15_6 ));
    Odrv4 I__13381 (
            .O(N__57857),
            .I(\c0.data_in_frame_15_6 ));
    InMux I__13380 (
            .O(N__57850),
            .I(N__57844));
    InMux I__13379 (
            .O(N__57849),
            .I(N__57844));
    LocalMux I__13378 (
            .O(N__57844),
            .I(N__57839));
    InMux I__13377 (
            .O(N__57843),
            .I(N__57834));
    InMux I__13376 (
            .O(N__57842),
            .I(N__57834));
    Odrv4 I__13375 (
            .O(N__57839),
            .I(\c0.n4_adj_4240 ));
    LocalMux I__13374 (
            .O(N__57834),
            .I(\c0.n4_adj_4240 ));
    CascadeMux I__13373 (
            .O(N__57829),
            .I(\c0.n22352_cascade_ ));
    CascadeMux I__13372 (
            .O(N__57826),
            .I(\c0.n22000_cascade_ ));
    InMux I__13371 (
            .O(N__57823),
            .I(N__57820));
    LocalMux I__13370 (
            .O(N__57820),
            .I(\c0.n31 ));
    InMux I__13369 (
            .O(N__57817),
            .I(N__57814));
    LocalMux I__13368 (
            .O(N__57814),
            .I(N__57811));
    Span4Mux_h I__13367 (
            .O(N__57811),
            .I(N__57806));
    InMux I__13366 (
            .O(N__57810),
            .I(N__57801));
    InMux I__13365 (
            .O(N__57809),
            .I(N__57801));
    Odrv4 I__13364 (
            .O(N__57806),
            .I(\c0.data_in_frame_15_7 ));
    LocalMux I__13363 (
            .O(N__57801),
            .I(\c0.data_in_frame_15_7 ));
    CascadeMux I__13362 (
            .O(N__57796),
            .I(N__57792));
    CascadeMux I__13361 (
            .O(N__57795),
            .I(N__57789));
    InMux I__13360 (
            .O(N__57792),
            .I(N__57786));
    InMux I__13359 (
            .O(N__57789),
            .I(N__57783));
    LocalMux I__13358 (
            .O(N__57786),
            .I(\c0.data_in_frame_18_2 ));
    LocalMux I__13357 (
            .O(N__57783),
            .I(\c0.data_in_frame_18_2 ));
    InMux I__13356 (
            .O(N__57778),
            .I(N__57775));
    LocalMux I__13355 (
            .O(N__57775),
            .I(N__57772));
    Odrv4 I__13354 (
            .O(N__57772),
            .I(\c0.n22000 ));
    CascadeMux I__13353 (
            .O(N__57769),
            .I(\c0.n12_cascade_ ));
    InMux I__13352 (
            .O(N__57766),
            .I(N__57763));
    LocalMux I__13351 (
            .O(N__57763),
            .I(N__57760));
    Odrv12 I__13350 (
            .O(N__57760),
            .I(\c0.n10_adj_4239 ));
    CascadeMux I__13349 (
            .O(N__57757),
            .I(N__57753));
    InMux I__13348 (
            .O(N__57756),
            .I(N__57750));
    InMux I__13347 (
            .O(N__57753),
            .I(N__57747));
    LocalMux I__13346 (
            .O(N__57750),
            .I(\c0.data_in_frame_18_0 ));
    LocalMux I__13345 (
            .O(N__57747),
            .I(\c0.data_in_frame_18_0 ));
    InMux I__13344 (
            .O(N__57742),
            .I(N__57739));
    LocalMux I__13343 (
            .O(N__57739),
            .I(\c0.n14_adj_4238 ));
    CascadeMux I__13342 (
            .O(N__57736),
            .I(\c0.n13210_cascade_ ));
    InMux I__13341 (
            .O(N__57733),
            .I(N__57727));
    InMux I__13340 (
            .O(N__57732),
            .I(N__57724));
    CascadeMux I__13339 (
            .O(N__57731),
            .I(N__57721));
    InMux I__13338 (
            .O(N__57730),
            .I(N__57718));
    LocalMux I__13337 (
            .O(N__57727),
            .I(N__57713));
    LocalMux I__13336 (
            .O(N__57724),
            .I(N__57713));
    InMux I__13335 (
            .O(N__57721),
            .I(N__57709));
    LocalMux I__13334 (
            .O(N__57718),
            .I(N__57706));
    Span4Mux_h I__13333 (
            .O(N__57713),
            .I(N__57703));
    InMux I__13332 (
            .O(N__57712),
            .I(N__57700));
    LocalMux I__13331 (
            .O(N__57709),
            .I(\c0.data_in_frame_8_7 ));
    Odrv12 I__13330 (
            .O(N__57706),
            .I(\c0.data_in_frame_8_7 ));
    Odrv4 I__13329 (
            .O(N__57703),
            .I(\c0.data_in_frame_8_7 ));
    LocalMux I__13328 (
            .O(N__57700),
            .I(\c0.data_in_frame_8_7 ));
    InMux I__13327 (
            .O(N__57691),
            .I(N__57688));
    LocalMux I__13326 (
            .O(N__57688),
            .I(N__57685));
    Odrv4 I__13325 (
            .O(N__57685),
            .I(\c0.n21822 ));
    CascadeMux I__13324 (
            .O(N__57682),
            .I(\c0.n7_adj_4277_cascade_ ));
    CascadeMux I__13323 (
            .O(N__57679),
            .I(N__57676));
    InMux I__13322 (
            .O(N__57676),
            .I(N__57671));
    InMux I__13321 (
            .O(N__57675),
            .I(N__57668));
    InMux I__13320 (
            .O(N__57674),
            .I(N__57665));
    LocalMux I__13319 (
            .O(N__57671),
            .I(\c0.data_in_frame_11_5 ));
    LocalMux I__13318 (
            .O(N__57668),
            .I(\c0.data_in_frame_11_5 ));
    LocalMux I__13317 (
            .O(N__57665),
            .I(\c0.data_in_frame_11_5 ));
    CascadeMux I__13316 (
            .O(N__57658),
            .I(\c0.n10_adj_4264_cascade_ ));
    InMux I__13315 (
            .O(N__57655),
            .I(N__57652));
    LocalMux I__13314 (
            .O(N__57652),
            .I(N__57649));
    Span4Mux_h I__13313 (
            .O(N__57649),
            .I(N__57646));
    Odrv4 I__13312 (
            .O(N__57646),
            .I(\c0.n16_adj_4265 ));
    InMux I__13311 (
            .O(N__57643),
            .I(N__57640));
    LocalMux I__13310 (
            .O(N__57640),
            .I(N__57636));
    CascadeMux I__13309 (
            .O(N__57639),
            .I(N__57633));
    Span4Mux_h I__13308 (
            .O(N__57636),
            .I(N__57629));
    InMux I__13307 (
            .O(N__57633),
            .I(N__57624));
    InMux I__13306 (
            .O(N__57632),
            .I(N__57624));
    Odrv4 I__13305 (
            .O(N__57629),
            .I(\c0.data_in_frame_11_6 ));
    LocalMux I__13304 (
            .O(N__57624),
            .I(\c0.data_in_frame_11_6 ));
    CascadeMux I__13303 (
            .O(N__57619),
            .I(N__57616));
    InMux I__13302 (
            .O(N__57616),
            .I(N__57609));
    InMux I__13301 (
            .O(N__57615),
            .I(N__57609));
    CascadeMux I__13300 (
            .O(N__57614),
            .I(N__57606));
    LocalMux I__13299 (
            .O(N__57609),
            .I(N__57602));
    InMux I__13298 (
            .O(N__57606),
            .I(N__57597));
    InMux I__13297 (
            .O(N__57605),
            .I(N__57597));
    Odrv12 I__13296 (
            .O(N__57602),
            .I(\c0.data_in_frame_11_2 ));
    LocalMux I__13295 (
            .O(N__57597),
            .I(\c0.data_in_frame_11_2 ));
    InMux I__13294 (
            .O(N__57592),
            .I(N__57589));
    LocalMux I__13293 (
            .O(N__57589),
            .I(N__57586));
    Span4Mux_h I__13292 (
            .O(N__57586),
            .I(N__57578));
    InMux I__13291 (
            .O(N__57585),
            .I(N__57573));
    InMux I__13290 (
            .O(N__57584),
            .I(N__57573));
    InMux I__13289 (
            .O(N__57583),
            .I(N__57570));
    InMux I__13288 (
            .O(N__57582),
            .I(N__57567));
    InMux I__13287 (
            .O(N__57581),
            .I(N__57564));
    Odrv4 I__13286 (
            .O(N__57578),
            .I(\c0.n20135 ));
    LocalMux I__13285 (
            .O(N__57573),
            .I(\c0.n20135 ));
    LocalMux I__13284 (
            .O(N__57570),
            .I(\c0.n20135 ));
    LocalMux I__13283 (
            .O(N__57567),
            .I(\c0.n20135 ));
    LocalMux I__13282 (
            .O(N__57564),
            .I(\c0.n20135 ));
    CascadeMux I__13281 (
            .O(N__57553),
            .I(N__57550));
    InMux I__13280 (
            .O(N__57550),
            .I(N__57547));
    LocalMux I__13279 (
            .O(N__57547),
            .I(N__57544));
    Odrv4 I__13278 (
            .O(N__57544),
            .I(\c0.n22464 ));
    InMux I__13277 (
            .O(N__57541),
            .I(N__57537));
    InMux I__13276 (
            .O(N__57540),
            .I(N__57534));
    LocalMux I__13275 (
            .O(N__57537),
            .I(\c0.n21867 ));
    LocalMux I__13274 (
            .O(N__57534),
            .I(\c0.n21867 ));
    InMux I__13273 (
            .O(N__57529),
            .I(N__57526));
    LocalMux I__13272 (
            .O(N__57526),
            .I(\c0.n6_adj_4225 ));
    InMux I__13271 (
            .O(N__57523),
            .I(N__57520));
    LocalMux I__13270 (
            .O(N__57520),
            .I(N__57517));
    Odrv4 I__13269 (
            .O(N__57517),
            .I(\c0.n15_adj_4269 ));
    CascadeMux I__13268 (
            .O(N__57514),
            .I(\c0.n22464_cascade_ ));
    InMux I__13267 (
            .O(N__57511),
            .I(N__57508));
    LocalMux I__13266 (
            .O(N__57508),
            .I(N__57505));
    Span4Mux_h I__13265 (
            .O(N__57505),
            .I(N__57502));
    Odrv4 I__13264 (
            .O(N__57502),
            .I(\c0.n22415 ));
    InMux I__13263 (
            .O(N__57499),
            .I(N__57493));
    InMux I__13262 (
            .O(N__57498),
            .I(N__57493));
    LocalMux I__13261 (
            .O(N__57493),
            .I(\c0.n13728 ));
    InMux I__13260 (
            .O(N__57490),
            .I(N__57486));
    InMux I__13259 (
            .O(N__57489),
            .I(N__57483));
    LocalMux I__13258 (
            .O(N__57486),
            .I(N__57480));
    LocalMux I__13257 (
            .O(N__57483),
            .I(N__57477));
    Span4Mux_h I__13256 (
            .O(N__57480),
            .I(N__57472));
    Span4Mux_v I__13255 (
            .O(N__57477),
            .I(N__57472));
    Odrv4 I__13254 (
            .O(N__57472),
            .I(\c0.n14053 ));
    CascadeMux I__13253 (
            .O(N__57469),
            .I(N__57465));
    InMux I__13252 (
            .O(N__57468),
            .I(N__57462));
    InMux I__13251 (
            .O(N__57465),
            .I(N__57459));
    LocalMux I__13250 (
            .O(N__57462),
            .I(N__57456));
    LocalMux I__13249 (
            .O(N__57459),
            .I(\c0.data_in_frame_18_1 ));
    Odrv4 I__13248 (
            .O(N__57456),
            .I(\c0.data_in_frame_18_1 ));
    CascadeMux I__13247 (
            .O(N__57451),
            .I(\c0.n14053_cascade_ ));
    InMux I__13246 (
            .O(N__57448),
            .I(N__57441));
    InMux I__13245 (
            .O(N__57447),
            .I(N__57438));
    InMux I__13244 (
            .O(N__57446),
            .I(N__57433));
    InMux I__13243 (
            .O(N__57445),
            .I(N__57433));
    CascadeMux I__13242 (
            .O(N__57444),
            .I(N__57430));
    LocalMux I__13241 (
            .O(N__57441),
            .I(N__57425));
    LocalMux I__13240 (
            .O(N__57438),
            .I(N__57425));
    LocalMux I__13239 (
            .O(N__57433),
            .I(N__57422));
    InMux I__13238 (
            .O(N__57430),
            .I(N__57419));
    Span12Mux_v I__13237 (
            .O(N__57425),
            .I(N__57416));
    Span4Mux_h I__13236 (
            .O(N__57422),
            .I(N__57413));
    LocalMux I__13235 (
            .O(N__57419),
            .I(\c0.data_in_frame_17_7 ));
    Odrv12 I__13234 (
            .O(N__57416),
            .I(\c0.data_in_frame_17_7 ));
    Odrv4 I__13233 (
            .O(N__57413),
            .I(\c0.data_in_frame_17_7 ));
    CascadeMux I__13232 (
            .O(N__57406),
            .I(\c0.n23586_cascade_ ));
    InMux I__13231 (
            .O(N__57403),
            .I(N__57400));
    LocalMux I__13230 (
            .O(N__57400),
            .I(N__57397));
    Span4Mux_h I__13229 (
            .O(N__57397),
            .I(N__57392));
    InMux I__13228 (
            .O(N__57396),
            .I(N__57387));
    InMux I__13227 (
            .O(N__57395),
            .I(N__57387));
    Odrv4 I__13226 (
            .O(N__57392),
            .I(\c0.data_in_frame_9_3 ));
    LocalMux I__13225 (
            .O(N__57387),
            .I(\c0.data_in_frame_9_3 ));
    InMux I__13224 (
            .O(N__57382),
            .I(N__57379));
    LocalMux I__13223 (
            .O(N__57379),
            .I(N__57376));
    Span4Mux_h I__13222 (
            .O(N__57376),
            .I(N__57373));
    Odrv4 I__13221 (
            .O(N__57373),
            .I(\c0.n22043 ));
    CascadeMux I__13220 (
            .O(N__57370),
            .I(N__57366));
    InMux I__13219 (
            .O(N__57369),
            .I(N__57362));
    InMux I__13218 (
            .O(N__57366),
            .I(N__57359));
    InMux I__13217 (
            .O(N__57365),
            .I(N__57356));
    LocalMux I__13216 (
            .O(N__57362),
            .I(N__57353));
    LocalMux I__13215 (
            .O(N__57359),
            .I(\c0.data_in_frame_9_7 ));
    LocalMux I__13214 (
            .O(N__57356),
            .I(\c0.data_in_frame_9_7 ));
    Odrv4 I__13213 (
            .O(N__57353),
            .I(\c0.data_in_frame_9_7 ));
    InMux I__13212 (
            .O(N__57346),
            .I(N__57342));
    InMux I__13211 (
            .O(N__57345),
            .I(N__57339));
    LocalMux I__13210 (
            .O(N__57342),
            .I(N__57336));
    LocalMux I__13209 (
            .O(N__57339),
            .I(N__57333));
    Span4Mux_v I__13208 (
            .O(N__57336),
            .I(N__57330));
    Odrv4 I__13207 (
            .O(N__57333),
            .I(\c0.n22471 ));
    Odrv4 I__13206 (
            .O(N__57330),
            .I(\c0.n22471 ));
    InMux I__13205 (
            .O(N__57325),
            .I(N__57321));
    CascadeMux I__13204 (
            .O(N__57324),
            .I(N__57318));
    LocalMux I__13203 (
            .O(N__57321),
            .I(N__57315));
    InMux I__13202 (
            .O(N__57318),
            .I(N__57310));
    Span12Mux_v I__13201 (
            .O(N__57315),
            .I(N__57307));
    InMux I__13200 (
            .O(N__57314),
            .I(N__57304));
    InMux I__13199 (
            .O(N__57313),
            .I(N__57301));
    LocalMux I__13198 (
            .O(N__57310),
            .I(\c0.data_in_frame_16_4 ));
    Odrv12 I__13197 (
            .O(N__57307),
            .I(\c0.data_in_frame_16_4 ));
    LocalMux I__13196 (
            .O(N__57304),
            .I(\c0.data_in_frame_16_4 ));
    LocalMux I__13195 (
            .O(N__57301),
            .I(\c0.data_in_frame_16_4 ));
    InMux I__13194 (
            .O(N__57292),
            .I(N__57286));
    InMux I__13193 (
            .O(N__57291),
            .I(N__57286));
    LocalMux I__13192 (
            .O(N__57286),
            .I(N__57280));
    InMux I__13191 (
            .O(N__57285),
            .I(N__57277));
    InMux I__13190 (
            .O(N__57284),
            .I(N__57274));
    InMux I__13189 (
            .O(N__57283),
            .I(N__57271));
    Span4Mux_v I__13188 (
            .O(N__57280),
            .I(N__57266));
    LocalMux I__13187 (
            .O(N__57277),
            .I(N__57266));
    LocalMux I__13186 (
            .O(N__57274),
            .I(N__57263));
    LocalMux I__13185 (
            .O(N__57271),
            .I(N__57258));
    Span4Mux_v I__13184 (
            .O(N__57266),
            .I(N__57258));
    Odrv12 I__13183 (
            .O(N__57263),
            .I(\c0.n20240 ));
    Odrv4 I__13182 (
            .O(N__57258),
            .I(\c0.n20240 ));
    CascadeMux I__13181 (
            .O(N__57253),
            .I(N__57250));
    InMux I__13180 (
            .O(N__57250),
            .I(N__57247));
    LocalMux I__13179 (
            .O(N__57247),
            .I(\c0.n22446 ));
    CascadeMux I__13178 (
            .O(N__57244),
            .I(N__57241));
    InMux I__13177 (
            .O(N__57241),
            .I(N__57238));
    LocalMux I__13176 (
            .O(N__57238),
            .I(N__57235));
    Span4Mux_h I__13175 (
            .O(N__57235),
            .I(N__57231));
    InMux I__13174 (
            .O(N__57234),
            .I(N__57228));
    Span4Mux_v I__13173 (
            .O(N__57231),
            .I(N__57225));
    LocalMux I__13172 (
            .O(N__57228),
            .I(\c0.n22328 ));
    Odrv4 I__13171 (
            .O(N__57225),
            .I(\c0.n22328 ));
    CascadeMux I__13170 (
            .O(N__57220),
            .I(\c0.n22446_cascade_ ));
    InMux I__13169 (
            .O(N__57217),
            .I(N__57213));
    InMux I__13168 (
            .O(N__57216),
            .I(N__57210));
    LocalMux I__13167 (
            .O(N__57213),
            .I(N__57207));
    LocalMux I__13166 (
            .O(N__57210),
            .I(N__57204));
    Odrv4 I__13165 (
            .O(N__57207),
            .I(\c0.n22424 ));
    Odrv4 I__13164 (
            .O(N__57204),
            .I(\c0.n22424 ));
    InMux I__13163 (
            .O(N__57199),
            .I(N__57196));
    LocalMux I__13162 (
            .O(N__57196),
            .I(N__57193));
    Span4Mux_v I__13161 (
            .O(N__57193),
            .I(N__57190));
    Odrv4 I__13160 (
            .O(N__57190),
            .I(\c0.n30_adj_4233 ));
    CascadeMux I__13159 (
            .O(N__57187),
            .I(N__57183));
    InMux I__13158 (
            .O(N__57186),
            .I(N__57178));
    InMux I__13157 (
            .O(N__57183),
            .I(N__57178));
    LocalMux I__13156 (
            .O(N__57178),
            .I(data_in_frame_14_2));
    InMux I__13155 (
            .O(N__57175),
            .I(N__57172));
    LocalMux I__13154 (
            .O(N__57172),
            .I(N__57169));
    Odrv4 I__13153 (
            .O(N__57169),
            .I(\c0.n22340 ));
    InMux I__13152 (
            .O(N__57166),
            .I(N__57163));
    LocalMux I__13151 (
            .O(N__57163),
            .I(N__57160));
    Span4Mux_v I__13150 (
            .O(N__57160),
            .I(N__57151));
    InMux I__13149 (
            .O(N__57159),
            .I(N__57146));
    InMux I__13148 (
            .O(N__57158),
            .I(N__57146));
    InMux I__13147 (
            .O(N__57157),
            .I(N__57143));
    InMux I__13146 (
            .O(N__57156),
            .I(N__57136));
    InMux I__13145 (
            .O(N__57155),
            .I(N__57136));
    InMux I__13144 (
            .O(N__57154),
            .I(N__57136));
    Odrv4 I__13143 (
            .O(N__57151),
            .I(n21755));
    LocalMux I__13142 (
            .O(N__57146),
            .I(n21755));
    LocalMux I__13141 (
            .O(N__57143),
            .I(n21755));
    LocalMux I__13140 (
            .O(N__57136),
            .I(n21755));
    InMux I__13139 (
            .O(N__57127),
            .I(N__57123));
    InMux I__13138 (
            .O(N__57126),
            .I(N__57120));
    LocalMux I__13137 (
            .O(N__57123),
            .I(data_in_frame_14_4));
    LocalMux I__13136 (
            .O(N__57120),
            .I(data_in_frame_14_4));
    InMux I__13135 (
            .O(N__57115),
            .I(N__57112));
    LocalMux I__13134 (
            .O(N__57112),
            .I(n19619));
    InMux I__13133 (
            .O(N__57109),
            .I(N__57106));
    LocalMux I__13132 (
            .O(N__57106),
            .I(N__57102));
    InMux I__13131 (
            .O(N__57105),
            .I(N__57098));
    Span4Mux_h I__13130 (
            .O(N__57102),
            .I(N__57095));
    CascadeMux I__13129 (
            .O(N__57101),
            .I(N__57092));
    LocalMux I__13128 (
            .O(N__57098),
            .I(N__57085));
    Sp12to4 I__13127 (
            .O(N__57095),
            .I(N__57085));
    InMux I__13126 (
            .O(N__57092),
            .I(N__57082));
    InMux I__13125 (
            .O(N__57091),
            .I(N__57079));
    InMux I__13124 (
            .O(N__57090),
            .I(N__57076));
    Span12Mux_v I__13123 (
            .O(N__57085),
            .I(N__57073));
    LocalMux I__13122 (
            .O(N__57082),
            .I(r_Bit_Index_2));
    LocalMux I__13121 (
            .O(N__57079),
            .I(r_Bit_Index_2));
    LocalMux I__13120 (
            .O(N__57076),
            .I(r_Bit_Index_2));
    Odrv12 I__13119 (
            .O(N__57073),
            .I(r_Bit_Index_2));
    CascadeMux I__13118 (
            .O(N__57064),
            .I(n91_cascade_));
    InMux I__13117 (
            .O(N__57061),
            .I(N__57055));
    InMux I__13116 (
            .O(N__57060),
            .I(N__57051));
    InMux I__13115 (
            .O(N__57059),
            .I(N__57048));
    InMux I__13114 (
            .O(N__57058),
            .I(N__57045));
    LocalMux I__13113 (
            .O(N__57055),
            .I(N__57042));
    InMux I__13112 (
            .O(N__57054),
            .I(N__57039));
    LocalMux I__13111 (
            .O(N__57051),
            .I(r_SM_Main_2_N_3681_2));
    LocalMux I__13110 (
            .O(N__57048),
            .I(r_SM_Main_2_N_3681_2));
    LocalMux I__13109 (
            .O(N__57045),
            .I(r_SM_Main_2_N_3681_2));
    Odrv4 I__13108 (
            .O(N__57042),
            .I(r_SM_Main_2_N_3681_2));
    LocalMux I__13107 (
            .O(N__57039),
            .I(r_SM_Main_2_N_3681_2));
    InMux I__13106 (
            .O(N__57028),
            .I(N__57024));
    InMux I__13105 (
            .O(N__57027),
            .I(N__57021));
    LocalMux I__13104 (
            .O(N__57024),
            .I(N__57018));
    LocalMux I__13103 (
            .O(N__57021),
            .I(N__57015));
    Span4Mux_v I__13102 (
            .O(N__57018),
            .I(N__57012));
    Span4Mux_h I__13101 (
            .O(N__57015),
            .I(N__57009));
    Sp12to4 I__13100 (
            .O(N__57012),
            .I(N__57004));
    Span4Mux_v I__13099 (
            .O(N__57009),
            .I(N__56999));
    InMux I__13098 (
            .O(N__57008),
            .I(N__56994));
    InMux I__13097 (
            .O(N__57007),
            .I(N__56994));
    Span12Mux_v I__13096 (
            .O(N__57004),
            .I(N__56988));
    InMux I__13095 (
            .O(N__57003),
            .I(N__56985));
    InMux I__13094 (
            .O(N__57002),
            .I(N__56982));
    Span4Mux_h I__13093 (
            .O(N__56999),
            .I(N__56979));
    LocalMux I__13092 (
            .O(N__56994),
            .I(N__56976));
    InMux I__13091 (
            .O(N__56993),
            .I(N__56973));
    InMux I__13090 (
            .O(N__56992),
            .I(N__56970));
    InMux I__13089 (
            .O(N__56991),
            .I(N__56967));
    Odrv12 I__13088 (
            .O(N__56988),
            .I(r_SM_Main_2));
    LocalMux I__13087 (
            .O(N__56985),
            .I(r_SM_Main_2));
    LocalMux I__13086 (
            .O(N__56982),
            .I(r_SM_Main_2));
    Odrv4 I__13085 (
            .O(N__56979),
            .I(r_SM_Main_2));
    Odrv4 I__13084 (
            .O(N__56976),
            .I(r_SM_Main_2));
    LocalMux I__13083 (
            .O(N__56973),
            .I(r_SM_Main_2));
    LocalMux I__13082 (
            .O(N__56970),
            .I(r_SM_Main_2));
    LocalMux I__13081 (
            .O(N__56967),
            .I(r_SM_Main_2));
    InMux I__13080 (
            .O(N__56950),
            .I(N__56947));
    LocalMux I__13079 (
            .O(N__56947),
            .I(N__56943));
    CascadeMux I__13078 (
            .O(N__56946),
            .I(N__56940));
    Span4Mux_v I__13077 (
            .O(N__56943),
            .I(N__56935));
    InMux I__13076 (
            .O(N__56940),
            .I(N__56929));
    InMux I__13075 (
            .O(N__56939),
            .I(N__56929));
    CascadeMux I__13074 (
            .O(N__56938),
            .I(N__56924));
    Span4Mux_v I__13073 (
            .O(N__56935),
            .I(N__56921));
    InMux I__13072 (
            .O(N__56934),
            .I(N__56918));
    LocalMux I__13071 (
            .O(N__56929),
            .I(N__56915));
    CascadeMux I__13070 (
            .O(N__56928),
            .I(N__56911));
    InMux I__13069 (
            .O(N__56927),
            .I(N__56905));
    InMux I__13068 (
            .O(N__56924),
            .I(N__56905));
    Span4Mux_v I__13067 (
            .O(N__56921),
            .I(N__56902));
    LocalMux I__13066 (
            .O(N__56918),
            .I(N__56899));
    Span4Mux_v I__13065 (
            .O(N__56915),
            .I(N__56895));
    InMux I__13064 (
            .O(N__56914),
            .I(N__56890));
    InMux I__13063 (
            .O(N__56911),
            .I(N__56890));
    CascadeMux I__13062 (
            .O(N__56910),
            .I(N__56886));
    LocalMux I__13061 (
            .O(N__56905),
            .I(N__56883));
    Span4Mux_h I__13060 (
            .O(N__56902),
            .I(N__56878));
    Span4Mux_v I__13059 (
            .O(N__56899),
            .I(N__56878));
    InMux I__13058 (
            .O(N__56898),
            .I(N__56875));
    Span4Mux_h I__13057 (
            .O(N__56895),
            .I(N__56870));
    LocalMux I__13056 (
            .O(N__56890),
            .I(N__56870));
    InMux I__13055 (
            .O(N__56889),
            .I(N__56867));
    InMux I__13054 (
            .O(N__56886),
            .I(N__56864));
    Span4Mux_h I__13053 (
            .O(N__56883),
            .I(N__56861));
    Span4Mux_h I__13052 (
            .O(N__56878),
            .I(N__56858));
    LocalMux I__13051 (
            .O(N__56875),
            .I(r_SM_Main_1));
    Odrv4 I__13050 (
            .O(N__56870),
            .I(r_SM_Main_1));
    LocalMux I__13049 (
            .O(N__56867),
            .I(r_SM_Main_1));
    LocalMux I__13048 (
            .O(N__56864),
            .I(r_SM_Main_1));
    Odrv4 I__13047 (
            .O(N__56861),
            .I(r_SM_Main_1));
    Odrv4 I__13046 (
            .O(N__56858),
            .I(r_SM_Main_1));
    CascadeMux I__13045 (
            .O(N__56845),
            .I(\c0.rx.n14_cascade_ ));
    InMux I__13044 (
            .O(N__56842),
            .I(N__56839));
    LocalMux I__13043 (
            .O(N__56839),
            .I(\c0.rx.n36 ));
    InMux I__13042 (
            .O(N__56836),
            .I(N__56832));
    InMux I__13041 (
            .O(N__56835),
            .I(N__56829));
    LocalMux I__13040 (
            .O(N__56832),
            .I(N__56823));
    LocalMux I__13039 (
            .O(N__56829),
            .I(N__56819));
    InMux I__13038 (
            .O(N__56828),
            .I(N__56811));
    InMux I__13037 (
            .O(N__56827),
            .I(N__56811));
    InMux I__13036 (
            .O(N__56826),
            .I(N__56811));
    Span12Mux_h I__13035 (
            .O(N__56823),
            .I(N__56805));
    InMux I__13034 (
            .O(N__56822),
            .I(N__56802));
    Span4Mux_h I__13033 (
            .O(N__56819),
            .I(N__56799));
    InMux I__13032 (
            .O(N__56818),
            .I(N__56796));
    LocalMux I__13031 (
            .O(N__56811),
            .I(N__56793));
    InMux I__13030 (
            .O(N__56810),
            .I(N__56788));
    InMux I__13029 (
            .O(N__56809),
            .I(N__56788));
    InMux I__13028 (
            .O(N__56808),
            .I(N__56785));
    Odrv12 I__13027 (
            .O(N__56805),
            .I(r_SM_Main_0));
    LocalMux I__13026 (
            .O(N__56802),
            .I(r_SM_Main_0));
    Odrv4 I__13025 (
            .O(N__56799),
            .I(r_SM_Main_0));
    LocalMux I__13024 (
            .O(N__56796),
            .I(r_SM_Main_0));
    Odrv12 I__13023 (
            .O(N__56793),
            .I(r_SM_Main_0));
    LocalMux I__13022 (
            .O(N__56788),
            .I(r_SM_Main_0));
    LocalMux I__13021 (
            .O(N__56785),
            .I(r_SM_Main_0));
    CascadeMux I__13020 (
            .O(N__56770),
            .I(n21755_cascade_));
    CascadeMux I__13019 (
            .O(N__56767),
            .I(N__56764));
    InMux I__13018 (
            .O(N__56764),
            .I(N__56760));
    InMux I__13017 (
            .O(N__56763),
            .I(N__56757));
    LocalMux I__13016 (
            .O(N__56760),
            .I(N__56754));
    LocalMux I__13015 (
            .O(N__56757),
            .I(data_in_frame_14_1));
    Odrv4 I__13014 (
            .O(N__56754),
            .I(data_in_frame_14_1));
    CascadeMux I__13013 (
            .O(N__56749),
            .I(N__56745));
    CascadeMux I__13012 (
            .O(N__56748),
            .I(N__56739));
    InMux I__13011 (
            .O(N__56745),
            .I(N__56736));
    CascadeMux I__13010 (
            .O(N__56744),
            .I(N__56733));
    CascadeMux I__13009 (
            .O(N__56743),
            .I(N__56730));
    CascadeMux I__13008 (
            .O(N__56742),
            .I(N__56726));
    InMux I__13007 (
            .O(N__56739),
            .I(N__56723));
    LocalMux I__13006 (
            .O(N__56736),
            .I(N__56720));
    InMux I__13005 (
            .O(N__56733),
            .I(N__56715));
    InMux I__13004 (
            .O(N__56730),
            .I(N__56712));
    InMux I__13003 (
            .O(N__56729),
            .I(N__56709));
    InMux I__13002 (
            .O(N__56726),
            .I(N__56705));
    LocalMux I__13001 (
            .O(N__56723),
            .I(N__56700));
    Span4Mux_v I__13000 (
            .O(N__56720),
            .I(N__56700));
    CascadeMux I__12999 (
            .O(N__56719),
            .I(N__56696));
    InMux I__12998 (
            .O(N__56718),
            .I(N__56693));
    LocalMux I__12997 (
            .O(N__56715),
            .I(N__56688));
    LocalMux I__12996 (
            .O(N__56712),
            .I(N__56683));
    LocalMux I__12995 (
            .O(N__56709),
            .I(N__56683));
    InMux I__12994 (
            .O(N__56708),
            .I(N__56680));
    LocalMux I__12993 (
            .O(N__56705),
            .I(N__56675));
    Span4Mux_v I__12992 (
            .O(N__56700),
            .I(N__56675));
    InMux I__12991 (
            .O(N__56699),
            .I(N__56672));
    InMux I__12990 (
            .O(N__56696),
            .I(N__56669));
    LocalMux I__12989 (
            .O(N__56693),
            .I(N__56666));
    InMux I__12988 (
            .O(N__56692),
            .I(N__56661));
    InMux I__12987 (
            .O(N__56691),
            .I(N__56661));
    Span4Mux_v I__12986 (
            .O(N__56688),
            .I(N__56658));
    Span4Mux_v I__12985 (
            .O(N__56683),
            .I(N__56653));
    LocalMux I__12984 (
            .O(N__56680),
            .I(N__56653));
    Span4Mux_v I__12983 (
            .O(N__56675),
            .I(N__56648));
    LocalMux I__12982 (
            .O(N__56672),
            .I(N__56648));
    LocalMux I__12981 (
            .O(N__56669),
            .I(N__56645));
    Span4Mux_v I__12980 (
            .O(N__56666),
            .I(N__56642));
    LocalMux I__12979 (
            .O(N__56661),
            .I(N__56639));
    Sp12to4 I__12978 (
            .O(N__56658),
            .I(N__56636));
    Span4Mux_h I__12977 (
            .O(N__56653),
            .I(N__56631));
    Span4Mux_v I__12976 (
            .O(N__56648),
            .I(N__56631));
    Span4Mux_v I__12975 (
            .O(N__56645),
            .I(N__56625));
    Span4Mux_v I__12974 (
            .O(N__56642),
            .I(N__56625));
    Span12Mux_h I__12973 (
            .O(N__56639),
            .I(N__56620));
    Span12Mux_v I__12972 (
            .O(N__56636),
            .I(N__56620));
    Span4Mux_v I__12971 (
            .O(N__56631),
            .I(N__56617));
    InMux I__12970 (
            .O(N__56630),
            .I(N__56614));
    Odrv4 I__12969 (
            .O(N__56625),
            .I(\c0.FRAME_MATCHER_i_0 ));
    Odrv12 I__12968 (
            .O(N__56620),
            .I(\c0.FRAME_MATCHER_i_0 ));
    Odrv4 I__12967 (
            .O(N__56617),
            .I(\c0.FRAME_MATCHER_i_0 ));
    LocalMux I__12966 (
            .O(N__56614),
            .I(\c0.FRAME_MATCHER_i_0 ));
    InMux I__12965 (
            .O(N__56605),
            .I(N__56602));
    LocalMux I__12964 (
            .O(N__56602),
            .I(N__56593));
    InMux I__12963 (
            .O(N__56601),
            .I(N__56590));
    InMux I__12962 (
            .O(N__56600),
            .I(N__56586));
    InMux I__12961 (
            .O(N__56599),
            .I(N__56583));
    InMux I__12960 (
            .O(N__56598),
            .I(N__56579));
    InMux I__12959 (
            .O(N__56597),
            .I(N__56574));
    InMux I__12958 (
            .O(N__56596),
            .I(N__56574));
    Span4Mux_h I__12957 (
            .O(N__56593),
            .I(N__56570));
    LocalMux I__12956 (
            .O(N__56590),
            .I(N__56565));
    InMux I__12955 (
            .O(N__56589),
            .I(N__56562));
    LocalMux I__12954 (
            .O(N__56586),
            .I(N__56557));
    LocalMux I__12953 (
            .O(N__56583),
            .I(N__56557));
    InMux I__12952 (
            .O(N__56582),
            .I(N__56554));
    LocalMux I__12951 (
            .O(N__56579),
            .I(N__56551));
    LocalMux I__12950 (
            .O(N__56574),
            .I(N__56548));
    InMux I__12949 (
            .O(N__56573),
            .I(N__56545));
    Span4Mux_v I__12948 (
            .O(N__56570),
            .I(N__56541));
    InMux I__12947 (
            .O(N__56569),
            .I(N__56538));
    InMux I__12946 (
            .O(N__56568),
            .I(N__56535));
    Span4Mux_v I__12945 (
            .O(N__56565),
            .I(N__56530));
    LocalMux I__12944 (
            .O(N__56562),
            .I(N__56530));
    Span4Mux_h I__12943 (
            .O(N__56557),
            .I(N__56527));
    LocalMux I__12942 (
            .O(N__56554),
            .I(N__56520));
    Span4Mux_h I__12941 (
            .O(N__56551),
            .I(N__56520));
    Span4Mux_v I__12940 (
            .O(N__56548),
            .I(N__56520));
    LocalMux I__12939 (
            .O(N__56545),
            .I(N__56517));
    CascadeMux I__12938 (
            .O(N__56544),
            .I(N__56514));
    Span4Mux_v I__12937 (
            .O(N__56541),
            .I(N__56507));
    LocalMux I__12936 (
            .O(N__56538),
            .I(N__56507));
    LocalMux I__12935 (
            .O(N__56535),
            .I(N__56507));
    Span4Mux_v I__12934 (
            .O(N__56530),
            .I(N__56504));
    Sp12to4 I__12933 (
            .O(N__56527),
            .I(N__56501));
    Span4Mux_h I__12932 (
            .O(N__56520),
            .I(N__56496));
    Span4Mux_h I__12931 (
            .O(N__56517),
            .I(N__56496));
    InMux I__12930 (
            .O(N__56514),
            .I(N__56492));
    Span4Mux_v I__12929 (
            .O(N__56507),
            .I(N__56487));
    Span4Mux_v I__12928 (
            .O(N__56504),
            .I(N__56487));
    Span12Mux_v I__12927 (
            .O(N__56501),
            .I(N__56484));
    Span4Mux_v I__12926 (
            .O(N__56496),
            .I(N__56481));
    InMux I__12925 (
            .O(N__56495),
            .I(N__56478));
    LocalMux I__12924 (
            .O(N__56492),
            .I(\c0.FRAME_MATCHER_i_1 ));
    Odrv4 I__12923 (
            .O(N__56487),
            .I(\c0.FRAME_MATCHER_i_1 ));
    Odrv12 I__12922 (
            .O(N__56484),
            .I(\c0.FRAME_MATCHER_i_1 ));
    Odrv4 I__12921 (
            .O(N__56481),
            .I(\c0.FRAME_MATCHER_i_1 ));
    LocalMux I__12920 (
            .O(N__56478),
            .I(\c0.FRAME_MATCHER_i_1 ));
    InMux I__12919 (
            .O(N__56467),
            .I(N__56462));
    InMux I__12918 (
            .O(N__56466),
            .I(N__56459));
    InMux I__12917 (
            .O(N__56465),
            .I(N__56452));
    LocalMux I__12916 (
            .O(N__56462),
            .I(N__56449));
    LocalMux I__12915 (
            .O(N__56459),
            .I(N__56446));
    CascadeMux I__12914 (
            .O(N__56458),
            .I(N__56443));
    InMux I__12913 (
            .O(N__56457),
            .I(N__56440));
    InMux I__12912 (
            .O(N__56456),
            .I(N__56436));
    InMux I__12911 (
            .O(N__56455),
            .I(N__56431));
    LocalMux I__12910 (
            .O(N__56452),
            .I(N__56428));
    Span4Mux_v I__12909 (
            .O(N__56449),
            .I(N__56423));
    Span4Mux_v I__12908 (
            .O(N__56446),
            .I(N__56423));
    InMux I__12907 (
            .O(N__56443),
            .I(N__56420));
    LocalMux I__12906 (
            .O(N__56440),
            .I(N__56416));
    InMux I__12905 (
            .O(N__56439),
            .I(N__56413));
    LocalMux I__12904 (
            .O(N__56436),
            .I(N__56410));
    InMux I__12903 (
            .O(N__56435),
            .I(N__56407));
    InMux I__12902 (
            .O(N__56434),
            .I(N__56404));
    LocalMux I__12901 (
            .O(N__56431),
            .I(N__56400));
    Span4Mux_v I__12900 (
            .O(N__56428),
            .I(N__56395));
    Span4Mux_v I__12899 (
            .O(N__56423),
            .I(N__56395));
    LocalMux I__12898 (
            .O(N__56420),
            .I(N__56391));
    InMux I__12897 (
            .O(N__56419),
            .I(N__56388));
    Span4Mux_v I__12896 (
            .O(N__56416),
            .I(N__56383));
    LocalMux I__12895 (
            .O(N__56413),
            .I(N__56383));
    Span4Mux_v I__12894 (
            .O(N__56410),
            .I(N__56376));
    LocalMux I__12893 (
            .O(N__56407),
            .I(N__56376));
    LocalMux I__12892 (
            .O(N__56404),
            .I(N__56376));
    CascadeMux I__12891 (
            .O(N__56403),
            .I(N__56373));
    Span4Mux_v I__12890 (
            .O(N__56400),
            .I(N__56370));
    Span4Mux_v I__12889 (
            .O(N__56395),
            .I(N__56367));
    InMux I__12888 (
            .O(N__56394),
            .I(N__56364));
    Span4Mux_h I__12887 (
            .O(N__56391),
            .I(N__56357));
    LocalMux I__12886 (
            .O(N__56388),
            .I(N__56357));
    Span4Mux_h I__12885 (
            .O(N__56383),
            .I(N__56357));
    Span4Mux_v I__12884 (
            .O(N__56376),
            .I(N__56354));
    InMux I__12883 (
            .O(N__56373),
            .I(N__56350));
    Span4Mux_v I__12882 (
            .O(N__56370),
            .I(N__56345));
    Span4Mux_v I__12881 (
            .O(N__56367),
            .I(N__56345));
    LocalMux I__12880 (
            .O(N__56364),
            .I(N__56338));
    Span4Mux_v I__12879 (
            .O(N__56357),
            .I(N__56338));
    Span4Mux_h I__12878 (
            .O(N__56354),
            .I(N__56338));
    InMux I__12877 (
            .O(N__56353),
            .I(N__56335));
    LocalMux I__12876 (
            .O(N__56350),
            .I(\c0.FRAME_MATCHER_i_2 ));
    Odrv4 I__12875 (
            .O(N__56345),
            .I(\c0.FRAME_MATCHER_i_2 ));
    Odrv4 I__12874 (
            .O(N__56338),
            .I(\c0.FRAME_MATCHER_i_2 ));
    LocalMux I__12873 (
            .O(N__56335),
            .I(\c0.FRAME_MATCHER_i_2 ));
    InMux I__12872 (
            .O(N__56326),
            .I(N__56323));
    LocalMux I__12871 (
            .O(N__56323),
            .I(N__56319));
    InMux I__12870 (
            .O(N__56322),
            .I(N__56316));
    Span4Mux_h I__12869 (
            .O(N__56319),
            .I(N__56311));
    LocalMux I__12868 (
            .O(N__56316),
            .I(N__56311));
    Odrv4 I__12867 (
            .O(N__56311),
            .I(\c0.n20370 ));
    CascadeMux I__12866 (
            .O(N__56308),
            .I(N__56305));
    InMux I__12865 (
            .O(N__56305),
            .I(N__56301));
    InMux I__12864 (
            .O(N__56304),
            .I(N__56298));
    LocalMux I__12863 (
            .O(N__56301),
            .I(\c0.data_in_frame_29_5 ));
    LocalMux I__12862 (
            .O(N__56298),
            .I(\c0.data_in_frame_29_5 ));
    InMux I__12861 (
            .O(N__56293),
            .I(N__56290));
    LocalMux I__12860 (
            .O(N__56290),
            .I(N__56287));
    Odrv4 I__12859 (
            .O(N__56287),
            .I(\c0.n22157 ));
    CascadeMux I__12858 (
            .O(N__56284),
            .I(N__56280));
    CascadeMux I__12857 (
            .O(N__56283),
            .I(N__56275));
    InMux I__12856 (
            .O(N__56280),
            .I(N__56272));
    InMux I__12855 (
            .O(N__56279),
            .I(N__56269));
    InMux I__12854 (
            .O(N__56278),
            .I(N__56266));
    InMux I__12853 (
            .O(N__56275),
            .I(N__56263));
    LocalMux I__12852 (
            .O(N__56272),
            .I(N__56258));
    LocalMux I__12851 (
            .O(N__56269),
            .I(N__56258));
    LocalMux I__12850 (
            .O(N__56266),
            .I(N__56253));
    LocalMux I__12849 (
            .O(N__56263),
            .I(N__56253));
    Odrv4 I__12848 (
            .O(N__56258),
            .I(\c0.data_in_frame_27_3 ));
    Odrv12 I__12847 (
            .O(N__56253),
            .I(\c0.data_in_frame_27_3 ));
    InMux I__12846 (
            .O(N__56248),
            .I(N__56245));
    LocalMux I__12845 (
            .O(N__56245),
            .I(\c0.n22719 ));
    CascadeMux I__12844 (
            .O(N__56242),
            .I(\c0.n8_adj_4291_cascade_ ));
    InMux I__12843 (
            .O(N__56239),
            .I(N__56236));
    LocalMux I__12842 (
            .O(N__56236),
            .I(\c0.n22148 ));
    InMux I__12841 (
            .O(N__56233),
            .I(N__56230));
    LocalMux I__12840 (
            .O(N__56230),
            .I(N__56227));
    Span4Mux_h I__12839 (
            .O(N__56227),
            .I(N__56224));
    Odrv4 I__12838 (
            .O(N__56224),
            .I(\c0.n23811 ));
    InMux I__12837 (
            .O(N__56221),
            .I(N__56217));
    CascadeMux I__12836 (
            .O(N__56220),
            .I(N__56214));
    LocalMux I__12835 (
            .O(N__56217),
            .I(N__56211));
    InMux I__12834 (
            .O(N__56214),
            .I(N__56208));
    Span4Mux_h I__12833 (
            .O(N__56211),
            .I(N__56204));
    LocalMux I__12832 (
            .O(N__56208),
            .I(N__56201));
    InMux I__12831 (
            .O(N__56207),
            .I(N__56198));
    Span4Mux_v I__12830 (
            .O(N__56204),
            .I(N__56195));
    Odrv4 I__12829 (
            .O(N__56201),
            .I(n12977));
    LocalMux I__12828 (
            .O(N__56198),
            .I(n12977));
    Odrv4 I__12827 (
            .O(N__56195),
            .I(n12977));
    InMux I__12826 (
            .O(N__56188),
            .I(N__56181));
    InMux I__12825 (
            .O(N__56187),
            .I(N__56181));
    InMux I__12824 (
            .O(N__56186),
            .I(N__56178));
    LocalMux I__12823 (
            .O(N__56181),
            .I(N__56175));
    LocalMux I__12822 (
            .O(N__56178),
            .I(N__56172));
    Span4Mux_v I__12821 (
            .O(N__56175),
            .I(N__56169));
    Odrv4 I__12820 (
            .O(N__56172),
            .I(\c0.rx.n21704 ));
    Odrv4 I__12819 (
            .O(N__56169),
            .I(\c0.rx.n21704 ));
    CascadeMux I__12818 (
            .O(N__56164),
            .I(n14436_cascade_));
    InMux I__12817 (
            .O(N__56161),
            .I(N__56157));
    InMux I__12816 (
            .O(N__56160),
            .I(N__56154));
    LocalMux I__12815 (
            .O(N__56157),
            .I(\c0.rx.n12862 ));
    LocalMux I__12814 (
            .O(N__56154),
            .I(\c0.rx.n12862 ));
    CascadeMux I__12813 (
            .O(N__56149),
            .I(N__56146));
    InMux I__12812 (
            .O(N__56146),
            .I(N__56143));
    LocalMux I__12811 (
            .O(N__56143),
            .I(N__56139));
    InMux I__12810 (
            .O(N__56142),
            .I(N__56135));
    Span4Mux_v I__12809 (
            .O(N__56139),
            .I(N__56132));
    CascadeMux I__12808 (
            .O(N__56138),
            .I(N__56129));
    LocalMux I__12807 (
            .O(N__56135),
            .I(N__56126));
    Span4Mux_v I__12806 (
            .O(N__56132),
            .I(N__56123));
    InMux I__12805 (
            .O(N__56129),
            .I(N__56120));
    Span12Mux_v I__12804 (
            .O(N__56126),
            .I(N__56117));
    Span4Mux_h I__12803 (
            .O(N__56123),
            .I(N__56114));
    LocalMux I__12802 (
            .O(N__56120),
            .I(\c0.data_in_frame_25_1 ));
    Odrv12 I__12801 (
            .O(N__56117),
            .I(\c0.data_in_frame_25_1 ));
    Odrv4 I__12800 (
            .O(N__56114),
            .I(\c0.data_in_frame_25_1 ));
    InMux I__12799 (
            .O(N__56107),
            .I(N__56104));
    LocalMux I__12798 (
            .O(N__56104),
            .I(N__56101));
    Span4Mux_v I__12797 (
            .O(N__56101),
            .I(N__56098));
    Span4Mux_h I__12796 (
            .O(N__56098),
            .I(N__56095));
    Odrv4 I__12795 (
            .O(N__56095),
            .I(\c0.n49_adj_4488 ));
    InMux I__12794 (
            .O(N__56092),
            .I(N__56089));
    LocalMux I__12793 (
            .O(N__56089),
            .I(\c0.n55 ));
    InMux I__12792 (
            .O(N__56086),
            .I(N__56083));
    LocalMux I__12791 (
            .O(N__56083),
            .I(\c0.n53 ));
    InMux I__12790 (
            .O(N__56080),
            .I(N__56077));
    LocalMux I__12789 (
            .O(N__56077),
            .I(N__56074));
    Span4Mux_h I__12788 (
            .O(N__56074),
            .I(N__56071));
    Odrv4 I__12787 (
            .O(N__56071),
            .I(\c0.n23416 ));
    CascadeMux I__12786 (
            .O(N__56068),
            .I(\c0.n23416_cascade_ ));
    InMux I__12785 (
            .O(N__56065),
            .I(N__56062));
    LocalMux I__12784 (
            .O(N__56062),
            .I(\c0.n12_adj_4296 ));
    InMux I__12783 (
            .O(N__56059),
            .I(N__56054));
    CascadeMux I__12782 (
            .O(N__56058),
            .I(N__56050));
    InMux I__12781 (
            .O(N__56057),
            .I(N__56047));
    LocalMux I__12780 (
            .O(N__56054),
            .I(N__56044));
    InMux I__12779 (
            .O(N__56053),
            .I(N__56041));
    InMux I__12778 (
            .O(N__56050),
            .I(N__56038));
    LocalMux I__12777 (
            .O(N__56047),
            .I(N__56035));
    Span4Mux_h I__12776 (
            .O(N__56044),
            .I(N__56032));
    LocalMux I__12775 (
            .O(N__56041),
            .I(N__56029));
    LocalMux I__12774 (
            .O(N__56038),
            .I(\c0.data_in_frame_27_2 ));
    Odrv4 I__12773 (
            .O(N__56035),
            .I(\c0.data_in_frame_27_2 ));
    Odrv4 I__12772 (
            .O(N__56032),
            .I(\c0.data_in_frame_27_2 ));
    Odrv12 I__12771 (
            .O(N__56029),
            .I(\c0.data_in_frame_27_2 ));
    InMux I__12770 (
            .O(N__56020),
            .I(N__56017));
    LocalMux I__12769 (
            .O(N__56017),
            .I(\c0.n36_adj_4489 ));
    CascadeMux I__12768 (
            .O(N__56014),
            .I(N__56011));
    InMux I__12767 (
            .O(N__56011),
            .I(N__56007));
    InMux I__12766 (
            .O(N__56010),
            .I(N__56003));
    LocalMux I__12765 (
            .O(N__56007),
            .I(N__56000));
    CascadeMux I__12764 (
            .O(N__56006),
            .I(N__55996));
    LocalMux I__12763 (
            .O(N__56003),
            .I(N__55993));
    Span4Mux_h I__12762 (
            .O(N__56000),
            .I(N__55990));
    InMux I__12761 (
            .O(N__55999),
            .I(N__55987));
    InMux I__12760 (
            .O(N__55996),
            .I(N__55984));
    Span4Mux_h I__12759 (
            .O(N__55993),
            .I(N__55981));
    Span4Mux_v I__12758 (
            .O(N__55990),
            .I(N__55978));
    LocalMux I__12757 (
            .O(N__55987),
            .I(N__55975));
    LocalMux I__12756 (
            .O(N__55984),
            .I(\c0.data_in_frame_19_2 ));
    Odrv4 I__12755 (
            .O(N__55981),
            .I(\c0.data_in_frame_19_2 ));
    Odrv4 I__12754 (
            .O(N__55978),
            .I(\c0.data_in_frame_19_2 ));
    Odrv4 I__12753 (
            .O(N__55975),
            .I(\c0.data_in_frame_19_2 ));
    InMux I__12752 (
            .O(N__55966),
            .I(N__55959));
    InMux I__12751 (
            .O(N__55965),
            .I(N__55959));
    InMux I__12750 (
            .O(N__55964),
            .I(N__55956));
    LocalMux I__12749 (
            .O(N__55959),
            .I(N__55953));
    LocalMux I__12748 (
            .O(N__55956),
            .I(N__55948));
    Span4Mux_v I__12747 (
            .O(N__55953),
            .I(N__55948));
    Odrv4 I__12746 (
            .O(N__55948),
            .I(\c0.n6221 ));
    CascadeMux I__12745 (
            .O(N__55945),
            .I(N__55942));
    InMux I__12744 (
            .O(N__55942),
            .I(N__55939));
    LocalMux I__12743 (
            .O(N__55939),
            .I(N__55935));
    InMux I__12742 (
            .O(N__55938),
            .I(N__55932));
    Span4Mux_h I__12741 (
            .O(N__55935),
            .I(N__55929));
    LocalMux I__12740 (
            .O(N__55932),
            .I(\c0.n21037 ));
    Odrv4 I__12739 (
            .O(N__55929),
            .I(\c0.n21037 ));
    InMux I__12738 (
            .O(N__55924),
            .I(N__55921));
    LocalMux I__12737 (
            .O(N__55921),
            .I(N__55916));
    InMux I__12736 (
            .O(N__55920),
            .I(N__55911));
    InMux I__12735 (
            .O(N__55919),
            .I(N__55911));
    Span4Mux_h I__12734 (
            .O(N__55916),
            .I(N__55908));
    LocalMux I__12733 (
            .O(N__55911),
            .I(N__55905));
    Odrv4 I__12732 (
            .O(N__55908),
            .I(\c0.data_in_frame_23_6 ));
    Odrv4 I__12731 (
            .O(N__55905),
            .I(\c0.data_in_frame_23_6 ));
    CascadeMux I__12730 (
            .O(N__55900),
            .I(\c0.n21037_cascade_ ));
    CascadeMux I__12729 (
            .O(N__55897),
            .I(N__55891));
    InMux I__12728 (
            .O(N__55896),
            .I(N__55887));
    InMux I__12727 (
            .O(N__55895),
            .I(N__55884));
    InMux I__12726 (
            .O(N__55894),
            .I(N__55877));
    InMux I__12725 (
            .O(N__55891),
            .I(N__55877));
    InMux I__12724 (
            .O(N__55890),
            .I(N__55877));
    LocalMux I__12723 (
            .O(N__55887),
            .I(N__55873));
    LocalMux I__12722 (
            .O(N__55884),
            .I(N__55870));
    LocalMux I__12721 (
            .O(N__55877),
            .I(N__55867));
    InMux I__12720 (
            .O(N__55876),
            .I(N__55864));
    Span4Mux_v I__12719 (
            .O(N__55873),
            .I(N__55861));
    Span4Mux_h I__12718 (
            .O(N__55870),
            .I(N__55858));
    Span4Mux_h I__12717 (
            .O(N__55867),
            .I(N__55855));
    LocalMux I__12716 (
            .O(N__55864),
            .I(\c0.data_in_frame_19_4 ));
    Odrv4 I__12715 (
            .O(N__55861),
            .I(\c0.data_in_frame_19_4 ));
    Odrv4 I__12714 (
            .O(N__55858),
            .I(\c0.data_in_frame_19_4 ));
    Odrv4 I__12713 (
            .O(N__55855),
            .I(\c0.data_in_frame_19_4 ));
    InMux I__12712 (
            .O(N__55846),
            .I(N__55843));
    LocalMux I__12711 (
            .O(N__55843),
            .I(\c0.n13282 ));
    CascadeMux I__12710 (
            .O(N__55840),
            .I(N__55836));
    CascadeMux I__12709 (
            .O(N__55839),
            .I(N__55833));
    InMux I__12708 (
            .O(N__55836),
            .I(N__55830));
    InMux I__12707 (
            .O(N__55833),
            .I(N__55826));
    LocalMux I__12706 (
            .O(N__55830),
            .I(N__55823));
    InMux I__12705 (
            .O(N__55829),
            .I(N__55820));
    LocalMux I__12704 (
            .O(N__55826),
            .I(N__55815));
    Span4Mux_h I__12703 (
            .O(N__55823),
            .I(N__55815));
    LocalMux I__12702 (
            .O(N__55820),
            .I(\c0.data_in_frame_27_4 ));
    Odrv4 I__12701 (
            .O(N__55815),
            .I(\c0.data_in_frame_27_4 ));
    CascadeMux I__12700 (
            .O(N__55810),
            .I(\c0.n52_cascade_ ));
    InMux I__12699 (
            .O(N__55807),
            .I(N__55804));
    LocalMux I__12698 (
            .O(N__55804),
            .I(N__55801));
    Odrv4 I__12697 (
            .O(N__55801),
            .I(\c0.n13872 ));
    InMux I__12696 (
            .O(N__55798),
            .I(N__55795));
    LocalMux I__12695 (
            .O(N__55795),
            .I(N__55791));
    InMux I__12694 (
            .O(N__55794),
            .I(N__55788));
    Odrv12 I__12693 (
            .O(N__55791),
            .I(\c0.n12420 ));
    LocalMux I__12692 (
            .O(N__55788),
            .I(\c0.n12420 ));
    InMux I__12691 (
            .O(N__55783),
            .I(N__55780));
    LocalMux I__12690 (
            .O(N__55780),
            .I(N__55777));
    Odrv4 I__12689 (
            .O(N__55777),
            .I(\c0.n23615 ));
    InMux I__12688 (
            .O(N__55774),
            .I(N__55771));
    LocalMux I__12687 (
            .O(N__55771),
            .I(\c0.n44_adj_4490 ));
    CascadeMux I__12686 (
            .O(N__55768),
            .I(\c0.n48_adj_4485_cascade_ ));
    InMux I__12685 (
            .O(N__55765),
            .I(N__55762));
    LocalMux I__12684 (
            .O(N__55762),
            .I(N__55759));
    Span4Mux_h I__12683 (
            .O(N__55759),
            .I(N__55756));
    Odrv4 I__12682 (
            .O(N__55756),
            .I(\c0.n12_adj_4290 ));
    InMux I__12681 (
            .O(N__55753),
            .I(N__55750));
    LocalMux I__12680 (
            .O(N__55750),
            .I(N__55746));
    InMux I__12679 (
            .O(N__55749),
            .I(N__55743));
    Span4Mux_v I__12678 (
            .O(N__55746),
            .I(N__55738));
    LocalMux I__12677 (
            .O(N__55743),
            .I(N__55738));
    Span4Mux_v I__12676 (
            .O(N__55738),
            .I(N__55735));
    Odrv4 I__12675 (
            .O(N__55735),
            .I(\c0.n22355 ));
    CascadeMux I__12674 (
            .O(N__55732),
            .I(\c0.n23062_cascade_ ));
    CascadeMux I__12673 (
            .O(N__55729),
            .I(N__55725));
    CascadeMux I__12672 (
            .O(N__55728),
            .I(N__55721));
    InMux I__12671 (
            .O(N__55725),
            .I(N__55718));
    InMux I__12670 (
            .O(N__55724),
            .I(N__55715));
    InMux I__12669 (
            .O(N__55721),
            .I(N__55712));
    LocalMux I__12668 (
            .O(N__55718),
            .I(N__55709));
    LocalMux I__12667 (
            .O(N__55715),
            .I(N__55706));
    LocalMux I__12666 (
            .O(N__55712),
            .I(N__55703));
    Span4Mux_v I__12665 (
            .O(N__55709),
            .I(N__55700));
    Span4Mux_v I__12664 (
            .O(N__55706),
            .I(N__55697));
    Odrv4 I__12663 (
            .O(N__55703),
            .I(\c0.data_in_frame_21_0 ));
    Odrv4 I__12662 (
            .O(N__55700),
            .I(\c0.data_in_frame_21_0 ));
    Odrv4 I__12661 (
            .O(N__55697),
            .I(\c0.data_in_frame_21_0 ));
    InMux I__12660 (
            .O(N__55690),
            .I(N__55687));
    LocalMux I__12659 (
            .O(N__55687),
            .I(\c0.n23062 ));
    InMux I__12658 (
            .O(N__55684),
            .I(N__55681));
    LocalMux I__12657 (
            .O(N__55681),
            .I(\c0.n8 ));
    InMux I__12656 (
            .O(N__55678),
            .I(N__55675));
    LocalMux I__12655 (
            .O(N__55675),
            .I(\c0.n27 ));
    InMux I__12654 (
            .O(N__55672),
            .I(N__55669));
    LocalMux I__12653 (
            .O(N__55669),
            .I(N__55665));
    InMux I__12652 (
            .O(N__55668),
            .I(N__55662));
    Span4Mux_v I__12651 (
            .O(N__55665),
            .I(N__55659));
    LocalMux I__12650 (
            .O(N__55662),
            .I(N__55656));
    Span4Mux_v I__12649 (
            .O(N__55659),
            .I(N__55653));
    Span4Mux_v I__12648 (
            .O(N__55656),
            .I(N__55650));
    Odrv4 I__12647 (
            .O(N__55653),
            .I(\c0.n22296 ));
    Odrv4 I__12646 (
            .O(N__55650),
            .I(\c0.n22296 ));
    InMux I__12645 (
            .O(N__55645),
            .I(N__55642));
    LocalMux I__12644 (
            .O(N__55642),
            .I(N__55638));
    InMux I__12643 (
            .O(N__55641),
            .I(N__55635));
    Span4Mux_v I__12642 (
            .O(N__55638),
            .I(N__55630));
    LocalMux I__12641 (
            .O(N__55635),
            .I(N__55630));
    Odrv4 I__12640 (
            .O(N__55630),
            .I(\c0.n21831 ));
    CascadeMux I__12639 (
            .O(N__55627),
            .I(N__55620));
    InMux I__12638 (
            .O(N__55626),
            .I(N__55617));
    InMux I__12637 (
            .O(N__55625),
            .I(N__55614));
    InMux I__12636 (
            .O(N__55624),
            .I(N__55609));
    InMux I__12635 (
            .O(N__55623),
            .I(N__55609));
    InMux I__12634 (
            .O(N__55620),
            .I(N__55606));
    LocalMux I__12633 (
            .O(N__55617),
            .I(N__55603));
    LocalMux I__12632 (
            .O(N__55614),
            .I(N__55600));
    LocalMux I__12631 (
            .O(N__55609),
            .I(N__55597));
    LocalMux I__12630 (
            .O(N__55606),
            .I(N__55594));
    Span4Mux_h I__12629 (
            .O(N__55603),
            .I(N__55591));
    Span4Mux_h I__12628 (
            .O(N__55600),
            .I(N__55588));
    Span4Mux_h I__12627 (
            .O(N__55597),
            .I(N__55585));
    Odrv4 I__12626 (
            .O(N__55594),
            .I(\c0.data_in_frame_17_0 ));
    Odrv4 I__12625 (
            .O(N__55591),
            .I(\c0.data_in_frame_17_0 ));
    Odrv4 I__12624 (
            .O(N__55588),
            .I(\c0.data_in_frame_17_0 ));
    Odrv4 I__12623 (
            .O(N__55585),
            .I(\c0.data_in_frame_17_0 ));
    CascadeMux I__12622 (
            .O(N__55576),
            .I(\c0.n16_adj_4223_cascade_ ));
    InMux I__12621 (
            .O(N__55573),
            .I(N__55570));
    LocalMux I__12620 (
            .O(N__55570),
            .I(N__55567));
    Odrv12 I__12619 (
            .O(N__55567),
            .I(\c0.n17 ));
    InMux I__12618 (
            .O(N__55564),
            .I(N__55558));
    InMux I__12617 (
            .O(N__55563),
            .I(N__55558));
    LocalMux I__12616 (
            .O(N__55558),
            .I(N__55554));
    InMux I__12615 (
            .O(N__55557),
            .I(N__55551));
    Span4Mux_h I__12614 (
            .O(N__55554),
            .I(N__55548));
    LocalMux I__12613 (
            .O(N__55551),
            .I(\c0.n21187 ));
    Odrv4 I__12612 (
            .O(N__55548),
            .I(\c0.n21187 ));
    CascadeMux I__12611 (
            .O(N__55543),
            .I(\c0.n22211_cascade_ ));
    InMux I__12610 (
            .O(N__55540),
            .I(N__55536));
    InMux I__12609 (
            .O(N__55539),
            .I(N__55531));
    LocalMux I__12608 (
            .O(N__55536),
            .I(N__55528));
    InMux I__12607 (
            .O(N__55535),
            .I(N__55525));
    InMux I__12606 (
            .O(N__55534),
            .I(N__55522));
    LocalMux I__12605 (
            .O(N__55531),
            .I(\c0.n21140 ));
    Odrv4 I__12604 (
            .O(N__55528),
            .I(\c0.n21140 ));
    LocalMux I__12603 (
            .O(N__55525),
            .I(\c0.n21140 ));
    LocalMux I__12602 (
            .O(N__55522),
            .I(\c0.n21140 ));
    InMux I__12601 (
            .O(N__55513),
            .I(N__55510));
    LocalMux I__12600 (
            .O(N__55510),
            .I(N__55506));
    InMux I__12599 (
            .O(N__55509),
            .I(N__55503));
    Odrv4 I__12598 (
            .O(N__55506),
            .I(\c0.n22311 ));
    LocalMux I__12597 (
            .O(N__55503),
            .I(\c0.n22311 ));
    InMux I__12596 (
            .O(N__55498),
            .I(N__55494));
    InMux I__12595 (
            .O(N__55497),
            .I(N__55491));
    LocalMux I__12594 (
            .O(N__55494),
            .I(\c0.n22211 ));
    LocalMux I__12593 (
            .O(N__55491),
            .I(\c0.n22211 ));
    InMux I__12592 (
            .O(N__55486),
            .I(N__55482));
    InMux I__12591 (
            .O(N__55485),
            .I(N__55479));
    LocalMux I__12590 (
            .O(N__55482),
            .I(N__55476));
    LocalMux I__12589 (
            .O(N__55479),
            .I(\c0.n23298 ));
    Odrv4 I__12588 (
            .O(N__55476),
            .I(\c0.n23298 ));
    InMux I__12587 (
            .O(N__55471),
            .I(N__55468));
    LocalMux I__12586 (
            .O(N__55468),
            .I(N__55465));
    Odrv4 I__12585 (
            .O(N__55465),
            .I(\c0.n7 ));
    CascadeMux I__12584 (
            .O(N__55462),
            .I(\c0.n23298_cascade_ ));
    InMux I__12583 (
            .O(N__55459),
            .I(N__55456));
    LocalMux I__12582 (
            .O(N__55456),
            .I(N__55453));
    Span4Mux_h I__12581 (
            .O(N__55453),
            .I(N__55450));
    Odrv4 I__12580 (
            .O(N__55450),
            .I(\c0.n45_adj_4486 ));
    InMux I__12579 (
            .O(N__55447),
            .I(N__55444));
    LocalMux I__12578 (
            .O(N__55444),
            .I(\c0.n22100 ));
    CascadeMux I__12577 (
            .O(N__55441),
            .I(\c0.n21054_cascade_ ));
    InMux I__12576 (
            .O(N__55438),
            .I(N__55435));
    LocalMux I__12575 (
            .O(N__55435),
            .I(\c0.n21043 ));
    InMux I__12574 (
            .O(N__55432),
            .I(N__55426));
    InMux I__12573 (
            .O(N__55431),
            .I(N__55421));
    InMux I__12572 (
            .O(N__55430),
            .I(N__55421));
    CascadeMux I__12571 (
            .O(N__55429),
            .I(N__55418));
    LocalMux I__12570 (
            .O(N__55426),
            .I(N__55412));
    LocalMux I__12569 (
            .O(N__55421),
            .I(N__55412));
    InMux I__12568 (
            .O(N__55418),
            .I(N__55409));
    InMux I__12567 (
            .O(N__55417),
            .I(N__55406));
    Span4Mux_h I__12566 (
            .O(N__55412),
            .I(N__55403));
    LocalMux I__12565 (
            .O(N__55409),
            .I(\c0.data_in_frame_17_3 ));
    LocalMux I__12564 (
            .O(N__55406),
            .I(\c0.data_in_frame_17_3 ));
    Odrv4 I__12563 (
            .O(N__55403),
            .I(\c0.data_in_frame_17_3 ));
    InMux I__12562 (
            .O(N__55396),
            .I(N__55389));
    InMux I__12561 (
            .O(N__55395),
            .I(N__55389));
    InMux I__12560 (
            .O(N__55394),
            .I(N__55386));
    LocalMux I__12559 (
            .O(N__55389),
            .I(N__55382));
    LocalMux I__12558 (
            .O(N__55386),
            .I(N__55379));
    InMux I__12557 (
            .O(N__55385),
            .I(N__55376));
    Span4Mux_v I__12556 (
            .O(N__55382),
            .I(N__55372));
    Span4Mux_h I__12555 (
            .O(N__55379),
            .I(N__55367));
    LocalMux I__12554 (
            .O(N__55376),
            .I(N__55367));
    InMux I__12553 (
            .O(N__55375),
            .I(N__55364));
    Span4Mux_h I__12552 (
            .O(N__55372),
            .I(N__55361));
    Span4Mux_h I__12551 (
            .O(N__55367),
            .I(N__55358));
    LocalMux I__12550 (
            .O(N__55364),
            .I(\c0.data_in_frame_17_4 ));
    Odrv4 I__12549 (
            .O(N__55361),
            .I(\c0.data_in_frame_17_4 ));
    Odrv4 I__12548 (
            .O(N__55358),
            .I(\c0.data_in_frame_17_4 ));
    InMux I__12547 (
            .O(N__55351),
            .I(N__55345));
    InMux I__12546 (
            .O(N__55350),
            .I(N__55345));
    LocalMux I__12545 (
            .O(N__55345),
            .I(N__55342));
    Odrv4 I__12544 (
            .O(N__55342),
            .I(\c0.n22480 ));
    InMux I__12543 (
            .O(N__55339),
            .I(N__55335));
    CascadeMux I__12542 (
            .O(N__55338),
            .I(N__55332));
    LocalMux I__12541 (
            .O(N__55335),
            .I(N__55329));
    InMux I__12540 (
            .O(N__55332),
            .I(N__55323));
    Span4Mux_h I__12539 (
            .O(N__55329),
            .I(N__55320));
    InMux I__12538 (
            .O(N__55328),
            .I(N__55317));
    InMux I__12537 (
            .O(N__55327),
            .I(N__55312));
    InMux I__12536 (
            .O(N__55326),
            .I(N__55312));
    LocalMux I__12535 (
            .O(N__55323),
            .I(\c0.data_in_frame_17_5 ));
    Odrv4 I__12534 (
            .O(N__55320),
            .I(\c0.data_in_frame_17_5 ));
    LocalMux I__12533 (
            .O(N__55317),
            .I(\c0.data_in_frame_17_5 ));
    LocalMux I__12532 (
            .O(N__55312),
            .I(\c0.data_in_frame_17_5 ));
    InMux I__12531 (
            .O(N__55303),
            .I(N__55299));
    InMux I__12530 (
            .O(N__55302),
            .I(N__55296));
    LocalMux I__12529 (
            .O(N__55299),
            .I(N__55293));
    LocalMux I__12528 (
            .O(N__55296),
            .I(N__55290));
    Span4Mux_v I__12527 (
            .O(N__55293),
            .I(N__55287));
    Odrv4 I__12526 (
            .O(N__55290),
            .I(\c0.n13719 ));
    Odrv4 I__12525 (
            .O(N__55287),
            .I(\c0.n13719 ));
    InMux I__12524 (
            .O(N__55282),
            .I(N__55279));
    LocalMux I__12523 (
            .O(N__55279),
            .I(\c0.n18 ));
    CascadeMux I__12522 (
            .O(N__55276),
            .I(N__55273));
    InMux I__12521 (
            .O(N__55273),
            .I(N__55270));
    LocalMux I__12520 (
            .O(N__55270),
            .I(N__55267));
    Span4Mux_h I__12519 (
            .O(N__55267),
            .I(N__55264));
    Odrv4 I__12518 (
            .O(N__55264),
            .I(\c0.n22349 ));
    InMux I__12517 (
            .O(N__55261),
            .I(N__55258));
    LocalMux I__12516 (
            .O(N__55258),
            .I(\c0.n30 ));
    InMux I__12515 (
            .O(N__55255),
            .I(N__55252));
    LocalMux I__12514 (
            .O(N__55252),
            .I(\c0.n22 ));
    InMux I__12513 (
            .O(N__55249),
            .I(N__55246));
    LocalMux I__12512 (
            .O(N__55246),
            .I(N__55243));
    Odrv4 I__12511 (
            .O(N__55243),
            .I(\c0.n7_adj_4235 ));
    InMux I__12510 (
            .O(N__55240),
            .I(N__55237));
    LocalMux I__12509 (
            .O(N__55237),
            .I(N__55234));
    Odrv4 I__12508 (
            .O(N__55234),
            .I(\c0.n8_adj_4236 ));
    CascadeMux I__12507 (
            .O(N__55231),
            .I(\c0.n20203_cascade_ ));
    InMux I__12506 (
            .O(N__55228),
            .I(N__55225));
    LocalMux I__12505 (
            .O(N__55225),
            .I(N__55222));
    Odrv4 I__12504 (
            .O(N__55222),
            .I(\c0.n21120 ));
    InMux I__12503 (
            .O(N__55219),
            .I(N__55214));
    CascadeMux I__12502 (
            .O(N__55218),
            .I(N__55211));
    InMux I__12501 (
            .O(N__55217),
            .I(N__55207));
    LocalMux I__12500 (
            .O(N__55214),
            .I(N__55204));
    InMux I__12499 (
            .O(N__55211),
            .I(N__55201));
    InMux I__12498 (
            .O(N__55210),
            .I(N__55198));
    LocalMux I__12497 (
            .O(N__55207),
            .I(N__55195));
    Sp12to4 I__12496 (
            .O(N__55204),
            .I(N__55192));
    LocalMux I__12495 (
            .O(N__55201),
            .I(\c0.data_in_frame_15_2 ));
    LocalMux I__12494 (
            .O(N__55198),
            .I(\c0.data_in_frame_15_2 ));
    Odrv4 I__12493 (
            .O(N__55195),
            .I(\c0.data_in_frame_15_2 ));
    Odrv12 I__12492 (
            .O(N__55192),
            .I(\c0.data_in_frame_15_2 ));
    InMux I__12491 (
            .O(N__55183),
            .I(N__55180));
    LocalMux I__12490 (
            .O(N__55180),
            .I(N__55177));
    Span4Mux_v I__12489 (
            .O(N__55177),
            .I(N__55174));
    Odrv4 I__12488 (
            .O(N__55174),
            .I(\c0.n22242 ));
    CascadeMux I__12487 (
            .O(N__55171),
            .I(N__55168));
    InMux I__12486 (
            .O(N__55168),
            .I(N__55165));
    LocalMux I__12485 (
            .O(N__55165),
            .I(N__55162));
    Span4Mux_h I__12484 (
            .O(N__55162),
            .I(N__55159));
    Odrv4 I__12483 (
            .O(N__55159),
            .I(\c0.n20402 ));
    InMux I__12482 (
            .O(N__55156),
            .I(N__55152));
    InMux I__12481 (
            .O(N__55155),
            .I(N__55149));
    LocalMux I__12480 (
            .O(N__55152),
            .I(\c0.n20196 ));
    LocalMux I__12479 (
            .O(N__55149),
            .I(\c0.n20196 ));
    CascadeMux I__12478 (
            .O(N__55144),
            .I(\c0.n13719_cascade_ ));
    InMux I__12477 (
            .O(N__55141),
            .I(N__55138));
    LocalMux I__12476 (
            .O(N__55138),
            .I(N__55134));
    InMux I__12475 (
            .O(N__55137),
            .I(N__55131));
    Odrv4 I__12474 (
            .O(N__55134),
            .I(\c0.n22221 ));
    LocalMux I__12473 (
            .O(N__55131),
            .I(\c0.n22221 ));
    InMux I__12472 (
            .O(N__55126),
            .I(N__55123));
    LocalMux I__12471 (
            .O(N__55123),
            .I(N__55120));
    Span4Mux_h I__12470 (
            .O(N__55120),
            .I(N__55115));
    InMux I__12469 (
            .O(N__55119),
            .I(N__55112));
    InMux I__12468 (
            .O(N__55118),
            .I(N__55109));
    Odrv4 I__12467 (
            .O(N__55115),
            .I(\c0.n13786 ));
    LocalMux I__12466 (
            .O(N__55112),
            .I(\c0.n13786 ));
    LocalMux I__12465 (
            .O(N__55109),
            .I(\c0.n13786 ));
    InMux I__12464 (
            .O(N__55102),
            .I(N__55098));
    InMux I__12463 (
            .O(N__55101),
            .I(N__55092));
    LocalMux I__12462 (
            .O(N__55098),
            .I(N__55089));
    InMux I__12461 (
            .O(N__55097),
            .I(N__55084));
    InMux I__12460 (
            .O(N__55096),
            .I(N__55084));
    InMux I__12459 (
            .O(N__55095),
            .I(N__55081));
    LocalMux I__12458 (
            .O(N__55092),
            .I(N__55078));
    Span4Mux_v I__12457 (
            .O(N__55089),
            .I(N__55073));
    LocalMux I__12456 (
            .O(N__55084),
            .I(N__55073));
    LocalMux I__12455 (
            .O(N__55081),
            .I(data_in_frame_14_6));
    Odrv12 I__12454 (
            .O(N__55078),
            .I(data_in_frame_14_6));
    Odrv4 I__12453 (
            .O(N__55073),
            .I(data_in_frame_14_6));
    InMux I__12452 (
            .O(N__55066),
            .I(N__55061));
    CascadeMux I__12451 (
            .O(N__55065),
            .I(N__55058));
    InMux I__12450 (
            .O(N__55064),
            .I(N__55054));
    LocalMux I__12449 (
            .O(N__55061),
            .I(N__55051));
    InMux I__12448 (
            .O(N__55058),
            .I(N__55048));
    InMux I__12447 (
            .O(N__55057),
            .I(N__55044));
    LocalMux I__12446 (
            .O(N__55054),
            .I(N__55037));
    Span4Mux_v I__12445 (
            .O(N__55051),
            .I(N__55037));
    LocalMux I__12444 (
            .O(N__55048),
            .I(N__55037));
    InMux I__12443 (
            .O(N__55047),
            .I(N__55034));
    LocalMux I__12442 (
            .O(N__55044),
            .I(data_in_frame_14_7));
    Odrv4 I__12441 (
            .O(N__55037),
            .I(data_in_frame_14_7));
    LocalMux I__12440 (
            .O(N__55034),
            .I(data_in_frame_14_7));
    CascadeMux I__12439 (
            .O(N__55027),
            .I(N__55024));
    InMux I__12438 (
            .O(N__55024),
            .I(N__55021));
    LocalMux I__12437 (
            .O(N__55021),
            .I(\c0.n5996 ));
    CascadeMux I__12436 (
            .O(N__55018),
            .I(\c0.n20222_cascade_ ));
    InMux I__12435 (
            .O(N__55015),
            .I(N__55012));
    LocalMux I__12434 (
            .O(N__55012),
            .I(N__55008));
    InMux I__12433 (
            .O(N__55011),
            .I(N__55005));
    Span4Mux_h I__12432 (
            .O(N__55008),
            .I(N__55000));
    LocalMux I__12431 (
            .O(N__55005),
            .I(N__55000));
    Span4Mux_v I__12430 (
            .O(N__55000),
            .I(N__54996));
    InMux I__12429 (
            .O(N__54999),
            .I(N__54993));
    Sp12to4 I__12428 (
            .O(N__54996),
            .I(N__54988));
    LocalMux I__12427 (
            .O(N__54993),
            .I(N__54988));
    Odrv12 I__12426 (
            .O(N__54988),
            .I(\c0.n13677 ));
    CascadeMux I__12425 (
            .O(N__54985),
            .I(\c0.n28_adj_4232_cascade_ ));
    CascadeMux I__12424 (
            .O(N__54982),
            .I(\c0.n32_cascade_ ));
    InMux I__12423 (
            .O(N__54979),
            .I(N__54976));
    LocalMux I__12422 (
            .O(N__54976),
            .I(N__54973));
    Odrv12 I__12421 (
            .O(N__54973),
            .I(\c0.n29_adj_4234 ));
    InMux I__12420 (
            .O(N__54970),
            .I(N__54967));
    LocalMux I__12419 (
            .O(N__54967),
            .I(N__54964));
    Span4Mux_h I__12418 (
            .O(N__54964),
            .I(N__54961));
    Odrv4 I__12417 (
            .O(N__54961),
            .I(\c0.n13681 ));
    CascadeMux I__12416 (
            .O(N__54958),
            .I(\c0.n21238_cascade_ ));
    InMux I__12415 (
            .O(N__54955),
            .I(N__54952));
    LocalMux I__12414 (
            .O(N__54952),
            .I(N__54948));
    InMux I__12413 (
            .O(N__54951),
            .I(N__54945));
    Span4Mux_h I__12412 (
            .O(N__54948),
            .I(N__54942));
    LocalMux I__12411 (
            .O(N__54945),
            .I(\c0.n21989 ));
    Odrv4 I__12410 (
            .O(N__54942),
            .I(\c0.n21989 ));
    InMux I__12409 (
            .O(N__54937),
            .I(N__54931));
    InMux I__12408 (
            .O(N__54936),
            .I(N__54931));
    LocalMux I__12407 (
            .O(N__54931),
            .I(\c0.n21238 ));
    InMux I__12406 (
            .O(N__54928),
            .I(N__54924));
    InMux I__12405 (
            .O(N__54927),
            .I(N__54921));
    LocalMux I__12404 (
            .O(N__54924),
            .I(N__54916));
    LocalMux I__12403 (
            .O(N__54921),
            .I(N__54916));
    Span4Mux_v I__12402 (
            .O(N__54916),
            .I(N__54913));
    Odrv4 I__12401 (
            .O(N__54913),
            .I(\c0.n22430 ));
    InMux I__12400 (
            .O(N__54910),
            .I(N__54907));
    LocalMux I__12399 (
            .O(N__54907),
            .I(N__54903));
    InMux I__12398 (
            .O(N__54906),
            .I(N__54900));
    Odrv4 I__12397 (
            .O(N__54903),
            .I(\c0.n5810 ));
    LocalMux I__12396 (
            .O(N__54900),
            .I(\c0.n5810 ));
    CascadeMux I__12395 (
            .O(N__54895),
            .I(N__54890));
    InMux I__12394 (
            .O(N__54894),
            .I(N__54886));
    CascadeMux I__12393 (
            .O(N__54893),
            .I(N__54883));
    InMux I__12392 (
            .O(N__54890),
            .I(N__54880));
    InMux I__12391 (
            .O(N__54889),
            .I(N__54877));
    LocalMux I__12390 (
            .O(N__54886),
            .I(N__54874));
    InMux I__12389 (
            .O(N__54883),
            .I(N__54871));
    LocalMux I__12388 (
            .O(N__54880),
            .I(N__54866));
    LocalMux I__12387 (
            .O(N__54877),
            .I(N__54866));
    Odrv4 I__12386 (
            .O(N__54874),
            .I(\c0.data_in_frame_7_1 ));
    LocalMux I__12385 (
            .O(N__54871),
            .I(\c0.data_in_frame_7_1 ));
    Odrv4 I__12384 (
            .O(N__54866),
            .I(\c0.data_in_frame_7_1 ));
    InMux I__12383 (
            .O(N__54859),
            .I(N__54856));
    LocalMux I__12382 (
            .O(N__54856),
            .I(\c0.n6_adj_4273 ));
    InMux I__12381 (
            .O(N__54853),
            .I(N__54850));
    LocalMux I__12380 (
            .O(N__54850),
            .I(\c0.n22139 ));
    CascadeMux I__12379 (
            .O(N__54847),
            .I(N__54844));
    InMux I__12378 (
            .O(N__54844),
            .I(N__54841));
    LocalMux I__12377 (
            .O(N__54841),
            .I(N__54838));
    Span4Mux_h I__12376 (
            .O(N__54838),
            .I(N__54835));
    Odrv4 I__12375 (
            .O(N__54835),
            .I(\c0.n6_adj_4243 ));
    InMux I__12374 (
            .O(N__54832),
            .I(N__54829));
    LocalMux I__12373 (
            .O(N__54829),
            .I(N__54825));
    InMux I__12372 (
            .O(N__54828),
            .I(N__54822));
    Span4Mux_v I__12371 (
            .O(N__54825),
            .I(N__54819));
    LocalMux I__12370 (
            .O(N__54822),
            .I(N__54816));
    Span4Mux_h I__12369 (
            .O(N__54819),
            .I(N__54812));
    Span4Mux_v I__12368 (
            .O(N__54816),
            .I(N__54809));
    InMux I__12367 (
            .O(N__54815),
            .I(N__54806));
    Odrv4 I__12366 (
            .O(N__54812),
            .I(\c0.n13861 ));
    Odrv4 I__12365 (
            .O(N__54809),
            .I(\c0.n13861 ));
    LocalMux I__12364 (
            .O(N__54806),
            .I(\c0.n13861 ));
    CascadeMux I__12363 (
            .O(N__54799),
            .I(\c0.n5813_cascade_ ));
    InMux I__12362 (
            .O(N__54796),
            .I(N__54792));
    InMux I__12361 (
            .O(N__54795),
            .I(N__54789));
    LocalMux I__12360 (
            .O(N__54792),
            .I(N__54784));
    LocalMux I__12359 (
            .O(N__54789),
            .I(N__54784));
    Span4Mux_v I__12358 (
            .O(N__54784),
            .I(N__54781));
    Odrv4 I__12357 (
            .O(N__54781),
            .I(\c0.n21967 ));
    InMux I__12356 (
            .O(N__54778),
            .I(N__54773));
    InMux I__12355 (
            .O(N__54777),
            .I(N__54768));
    InMux I__12354 (
            .O(N__54776),
            .I(N__54768));
    LocalMux I__12353 (
            .O(N__54773),
            .I(N__54761));
    LocalMux I__12352 (
            .O(N__54768),
            .I(N__54761));
    InMux I__12351 (
            .O(N__54767),
            .I(N__54756));
    InMux I__12350 (
            .O(N__54766),
            .I(N__54756));
    Odrv12 I__12349 (
            .O(N__54761),
            .I(\c0.n13237 ));
    LocalMux I__12348 (
            .O(N__54756),
            .I(\c0.n13237 ));
    InMux I__12347 (
            .O(N__54751),
            .I(N__54748));
    LocalMux I__12346 (
            .O(N__54748),
            .I(N__54743));
    InMux I__12345 (
            .O(N__54747),
            .I(N__54740));
    InMux I__12344 (
            .O(N__54746),
            .I(N__54737));
    Span4Mux_h I__12343 (
            .O(N__54743),
            .I(N__54734));
    LocalMux I__12342 (
            .O(N__54740),
            .I(N__54731));
    LocalMux I__12341 (
            .O(N__54737),
            .I(N__54726));
    Span4Mux_v I__12340 (
            .O(N__54734),
            .I(N__54726));
    Span4Mux_v I__12339 (
            .O(N__54731),
            .I(N__54723));
    Odrv4 I__12338 (
            .O(N__54726),
            .I(\c0.data_in_frame_7_6 ));
    Odrv4 I__12337 (
            .O(N__54723),
            .I(\c0.data_in_frame_7_6 ));
    InMux I__12336 (
            .O(N__54718),
            .I(N__54715));
    LocalMux I__12335 (
            .O(N__54715),
            .I(N__54711));
    InMux I__12334 (
            .O(N__54714),
            .I(N__54706));
    Span4Mux_h I__12333 (
            .O(N__54711),
            .I(N__54703));
    InMux I__12332 (
            .O(N__54710),
            .I(N__54700));
    InMux I__12331 (
            .O(N__54709),
            .I(N__54697));
    LocalMux I__12330 (
            .O(N__54706),
            .I(\c0.data_in_frame_10_0 ));
    Odrv4 I__12329 (
            .O(N__54703),
            .I(\c0.data_in_frame_10_0 ));
    LocalMux I__12328 (
            .O(N__54700),
            .I(\c0.data_in_frame_10_0 ));
    LocalMux I__12327 (
            .O(N__54697),
            .I(\c0.data_in_frame_10_0 ));
    CascadeMux I__12326 (
            .O(N__54688),
            .I(\c0.n10_adj_4245_cascade_ ));
    InMux I__12325 (
            .O(N__54685),
            .I(N__54679));
    InMux I__12324 (
            .O(N__54684),
            .I(N__54676));
    InMux I__12323 (
            .O(N__54683),
            .I(N__54673));
    InMux I__12322 (
            .O(N__54682),
            .I(N__54670));
    LocalMux I__12321 (
            .O(N__54679),
            .I(N__54667));
    LocalMux I__12320 (
            .O(N__54676),
            .I(N__54664));
    LocalMux I__12319 (
            .O(N__54673),
            .I(N__54660));
    LocalMux I__12318 (
            .O(N__54670),
            .I(N__54657));
    Span4Mux_h I__12317 (
            .O(N__54667),
            .I(N__54654));
    Span4Mux_v I__12316 (
            .O(N__54664),
            .I(N__54651));
    InMux I__12315 (
            .O(N__54663),
            .I(N__54648));
    Span4Mux_h I__12314 (
            .O(N__54660),
            .I(N__54643));
    Span4Mux_v I__12313 (
            .O(N__54657),
            .I(N__54643));
    Odrv4 I__12312 (
            .O(N__54654),
            .I(\c0.n13099 ));
    Odrv4 I__12311 (
            .O(N__54651),
            .I(\c0.n13099 ));
    LocalMux I__12310 (
            .O(N__54648),
            .I(\c0.n13099 ));
    Odrv4 I__12309 (
            .O(N__54643),
            .I(\c0.n13099 ));
    InMux I__12308 (
            .O(N__54634),
            .I(N__54630));
    CascadeMux I__12307 (
            .O(N__54633),
            .I(N__54627));
    LocalMux I__12306 (
            .O(N__54630),
            .I(N__54623));
    InMux I__12305 (
            .O(N__54627),
            .I(N__54618));
    InMux I__12304 (
            .O(N__54626),
            .I(N__54618));
    Odrv4 I__12303 (
            .O(N__54623),
            .I(\c0.data_in_frame_9_1 ));
    LocalMux I__12302 (
            .O(N__54618),
            .I(\c0.data_in_frame_9_1 ));
    InMux I__12301 (
            .O(N__54613),
            .I(N__54610));
    LocalMux I__12300 (
            .O(N__54610),
            .I(N__54607));
    Span4Mux_v I__12299 (
            .O(N__54607),
            .I(N__54604));
    Odrv4 I__12298 (
            .O(N__54604),
            .I(\c0.n14037 ));
    InMux I__12297 (
            .O(N__54601),
            .I(N__54595));
    InMux I__12296 (
            .O(N__54600),
            .I(N__54595));
    LocalMux I__12295 (
            .O(N__54595),
            .I(\c0.n22233 ));
    CascadeMux I__12294 (
            .O(N__54592),
            .I(N__54589));
    InMux I__12293 (
            .O(N__54589),
            .I(N__54584));
    InMux I__12292 (
            .O(N__54588),
            .I(N__54581));
    InMux I__12291 (
            .O(N__54587),
            .I(N__54578));
    LocalMux I__12290 (
            .O(N__54584),
            .I(\c0.data_in_frame_11_3 ));
    LocalMux I__12289 (
            .O(N__54581),
            .I(\c0.data_in_frame_11_3 ));
    LocalMux I__12288 (
            .O(N__54578),
            .I(\c0.data_in_frame_11_3 ));
    InMux I__12287 (
            .O(N__54571),
            .I(N__54568));
    LocalMux I__12286 (
            .O(N__54568),
            .I(\c0.n10_adj_4274 ));
    InMux I__12285 (
            .O(N__54565),
            .I(N__54562));
    LocalMux I__12284 (
            .O(N__54562),
            .I(N__54558));
    InMux I__12283 (
            .O(N__54561),
            .I(N__54555));
    Span4Mux_h I__12282 (
            .O(N__54558),
            .I(N__54552));
    LocalMux I__12281 (
            .O(N__54555),
            .I(N__54549));
    Odrv4 I__12280 (
            .O(N__54552),
            .I(\c0.n22108 ));
    Odrv4 I__12279 (
            .O(N__54549),
            .I(\c0.n22108 ));
    CascadeMux I__12278 (
            .O(N__54544),
            .I(\c0.n4_adj_4240_cascade_ ));
    InMux I__12277 (
            .O(N__54541),
            .I(N__54538));
    LocalMux I__12276 (
            .O(N__54538),
            .I(N__54535));
    Odrv4 I__12275 (
            .O(N__54535),
            .I(\c0.n22060 ));
    CascadeMux I__12274 (
            .O(N__54532),
            .I(\c0.n6_adj_4244_cascade_ ));
    InMux I__12273 (
            .O(N__54529),
            .I(N__54525));
    InMux I__12272 (
            .O(N__54528),
            .I(N__54522));
    LocalMux I__12271 (
            .O(N__54525),
            .I(N__54519));
    LocalMux I__12270 (
            .O(N__54522),
            .I(\c0.n21097 ));
    Odrv4 I__12269 (
            .O(N__54519),
            .I(\c0.n21097 ));
    CascadeMux I__12268 (
            .O(N__54514),
            .I(\c0.n20240_cascade_ ));
    InMux I__12267 (
            .O(N__54511),
            .I(N__54508));
    LocalMux I__12266 (
            .O(N__54508),
            .I(N__54504));
    CascadeMux I__12265 (
            .O(N__54507),
            .I(N__54501));
    Span4Mux_h I__12264 (
            .O(N__54504),
            .I(N__54497));
    InMux I__12263 (
            .O(N__54501),
            .I(N__54494));
    InMux I__12262 (
            .O(N__54500),
            .I(N__54491));
    Span4Mux_v I__12261 (
            .O(N__54497),
            .I(N__54488));
    LocalMux I__12260 (
            .O(N__54494),
            .I(\c0.data_in_frame_15_0 ));
    LocalMux I__12259 (
            .O(N__54491),
            .I(\c0.data_in_frame_15_0 ));
    Odrv4 I__12258 (
            .O(N__54488),
            .I(\c0.data_in_frame_15_0 ));
    CascadeMux I__12257 (
            .O(N__54481),
            .I(\c0.n22385_cascade_ ));
    CascadeMux I__12256 (
            .O(N__54478),
            .I(N__54474));
    InMux I__12255 (
            .O(N__54477),
            .I(N__54471));
    InMux I__12254 (
            .O(N__54474),
            .I(N__54468));
    LocalMux I__12253 (
            .O(N__54471),
            .I(N__54464));
    LocalMux I__12252 (
            .O(N__54468),
            .I(N__54461));
    InMux I__12251 (
            .O(N__54467),
            .I(N__54458));
    Span4Mux_v I__12250 (
            .O(N__54464),
            .I(N__54453));
    Span4Mux_h I__12249 (
            .O(N__54461),
            .I(N__54453));
    LocalMux I__12248 (
            .O(N__54458),
            .I(data_in_frame_14_5));
    Odrv4 I__12247 (
            .O(N__54453),
            .I(data_in_frame_14_5));
    InMux I__12246 (
            .O(N__54448),
            .I(N__54444));
    InMux I__12245 (
            .O(N__54447),
            .I(N__54441));
    LocalMux I__12244 (
            .O(N__54444),
            .I(data_in_frame_14_3));
    LocalMux I__12243 (
            .O(N__54441),
            .I(data_in_frame_14_3));
    CascadeMux I__12242 (
            .O(N__54436),
            .I(N__54433));
    InMux I__12241 (
            .O(N__54433),
            .I(N__54429));
    InMux I__12240 (
            .O(N__54432),
            .I(N__54426));
    LocalMux I__12239 (
            .O(N__54429),
            .I(\c0.data_in_frame_4_0 ));
    LocalMux I__12238 (
            .O(N__54426),
            .I(\c0.data_in_frame_4_0 ));
    InMux I__12237 (
            .O(N__54421),
            .I(N__54417));
    InMux I__12236 (
            .O(N__54420),
            .I(N__54414));
    LocalMux I__12235 (
            .O(N__54417),
            .I(N__54411));
    LocalMux I__12234 (
            .O(N__54414),
            .I(N__54408));
    Span4Mux_v I__12233 (
            .O(N__54411),
            .I(N__54404));
    Span4Mux_v I__12232 (
            .O(N__54408),
            .I(N__54401));
    CascadeMux I__12231 (
            .O(N__54407),
            .I(N__54396));
    Span4Mux_v I__12230 (
            .O(N__54404),
            .I(N__54390));
    Span4Mux_h I__12229 (
            .O(N__54401),
            .I(N__54390));
    InMux I__12228 (
            .O(N__54400),
            .I(N__54387));
    InMux I__12227 (
            .O(N__54399),
            .I(N__54384));
    InMux I__12226 (
            .O(N__54396),
            .I(N__54379));
    InMux I__12225 (
            .O(N__54395),
            .I(N__54379));
    Sp12to4 I__12224 (
            .O(N__54390),
            .I(N__54374));
    LocalMux I__12223 (
            .O(N__54387),
            .I(N__54374));
    LocalMux I__12222 (
            .O(N__54384),
            .I(data_in_frame_1_4));
    LocalMux I__12221 (
            .O(N__54379),
            .I(data_in_frame_1_4));
    Odrv12 I__12220 (
            .O(N__54374),
            .I(data_in_frame_1_4));
    InMux I__12219 (
            .O(N__54367),
            .I(N__54364));
    LocalMux I__12218 (
            .O(N__54364),
            .I(N__54360));
    InMux I__12217 (
            .O(N__54363),
            .I(N__54357));
    Span4Mux_v I__12216 (
            .O(N__54360),
            .I(N__54352));
    LocalMux I__12215 (
            .O(N__54357),
            .I(N__54352));
    Span4Mux_h I__12214 (
            .O(N__54352),
            .I(N__54349));
    Odrv4 I__12213 (
            .O(N__54349),
            .I(\c0.n21797 ));
    CascadeMux I__12212 (
            .O(N__54346),
            .I(r_SM_Main_2_N_3681_2_cascade_));
    CascadeMux I__12211 (
            .O(N__54343),
            .I(N__54340));
    InMux I__12210 (
            .O(N__54340),
            .I(N__54337));
    LocalMux I__12209 (
            .O(N__54337),
            .I(N__54334));
    Span12Mux_h I__12208 (
            .O(N__54334),
            .I(N__54331));
    Span12Mux_v I__12207 (
            .O(N__54331),
            .I(N__54328));
    Span12Mux_h I__12206 (
            .O(N__54328),
            .I(N__54325));
    Odrv12 I__12205 (
            .O(N__54325),
            .I(n14283));
    InMux I__12204 (
            .O(N__54322),
            .I(N__54316));
    InMux I__12203 (
            .O(N__54321),
            .I(N__54313));
    InMux I__12202 (
            .O(N__54320),
            .I(N__54308));
    InMux I__12201 (
            .O(N__54319),
            .I(N__54308));
    LocalMux I__12200 (
            .O(N__54316),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__12199 (
            .O(N__54313),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__12198 (
            .O(N__54308),
            .I(\c0.rx.r_Clock_Count_4 ));
    InMux I__12197 (
            .O(N__54301),
            .I(N__54297));
    InMux I__12196 (
            .O(N__54300),
            .I(N__54294));
    LocalMux I__12195 (
            .O(N__54297),
            .I(\c0.rx.n18655 ));
    LocalMux I__12194 (
            .O(N__54294),
            .I(\c0.rx.n18655 ));
    CascadeMux I__12193 (
            .O(N__54289),
            .I(N__54286));
    InMux I__12192 (
            .O(N__54286),
            .I(N__54280));
    InMux I__12191 (
            .O(N__54285),
            .I(N__54277));
    InMux I__12190 (
            .O(N__54284),
            .I(N__54274));
    InMux I__12189 (
            .O(N__54283),
            .I(N__54271));
    LocalMux I__12188 (
            .O(N__54280),
            .I(\c0.rx.r_Clock_Count_0 ));
    LocalMux I__12187 (
            .O(N__54277),
            .I(\c0.rx.r_Clock_Count_0 ));
    LocalMux I__12186 (
            .O(N__54274),
            .I(\c0.rx.r_Clock_Count_0 ));
    LocalMux I__12185 (
            .O(N__54271),
            .I(\c0.rx.r_Clock_Count_0 ));
    InMux I__12184 (
            .O(N__54262),
            .I(N__54258));
    InMux I__12183 (
            .O(N__54261),
            .I(N__54255));
    LocalMux I__12182 (
            .O(N__54258),
            .I(\c0.rx.n80 ));
    LocalMux I__12181 (
            .O(N__54255),
            .I(\c0.rx.n80 ));
    SRMux I__12180 (
            .O(N__54250),
            .I(N__54247));
    LocalMux I__12179 (
            .O(N__54247),
            .I(N__54244));
    Span4Mux_h I__12178 (
            .O(N__54244),
            .I(N__54241));
    Span4Mux_h I__12177 (
            .O(N__54241),
            .I(N__54238));
    Span4Mux_v I__12176 (
            .O(N__54238),
            .I(N__54235));
    Odrv4 I__12175 (
            .O(N__54235),
            .I(\c0.rx.n21783 ));
    InMux I__12174 (
            .O(N__54232),
            .I(N__54229));
    LocalMux I__12173 (
            .O(N__54229),
            .I(N__54226));
    Span4Mux_v I__12172 (
            .O(N__54226),
            .I(N__54223));
    Sp12to4 I__12171 (
            .O(N__54223),
            .I(N__54220));
    Span12Mux_h I__12170 (
            .O(N__54220),
            .I(N__54217));
    Odrv12 I__12169 (
            .O(N__54217),
            .I(\c0.rx.r_Rx_Data_R ));
    InMux I__12168 (
            .O(N__54214),
            .I(N__54210));
    CascadeMux I__12167 (
            .O(N__54213),
            .I(N__54207));
    LocalMux I__12166 (
            .O(N__54210),
            .I(N__54204));
    InMux I__12165 (
            .O(N__54207),
            .I(N__54201));
    Span4Mux_v I__12164 (
            .O(N__54204),
            .I(N__54198));
    LocalMux I__12163 (
            .O(N__54201),
            .I(\c0.data_in_frame_12_6 ));
    Odrv4 I__12162 (
            .O(N__54198),
            .I(\c0.data_in_frame_12_6 ));
    InMux I__12161 (
            .O(N__54193),
            .I(N__54190));
    LocalMux I__12160 (
            .O(N__54190),
            .I(N__54185));
    InMux I__12159 (
            .O(N__54189),
            .I(N__54180));
    InMux I__12158 (
            .O(N__54188),
            .I(N__54180));
    Odrv4 I__12157 (
            .O(N__54185),
            .I(\c0.data_in_frame_15_3 ));
    LocalMux I__12156 (
            .O(N__54180),
            .I(\c0.data_in_frame_15_3 ));
    InMux I__12155 (
            .O(N__54175),
            .I(N__54171));
    InMux I__12154 (
            .O(N__54174),
            .I(N__54168));
    LocalMux I__12153 (
            .O(N__54171),
            .I(N__54165));
    LocalMux I__12152 (
            .O(N__54168),
            .I(N__54161));
    Span4Mux_v I__12151 (
            .O(N__54165),
            .I(N__54158));
    InMux I__12150 (
            .O(N__54164),
            .I(N__54155));
    Odrv4 I__12149 (
            .O(N__54161),
            .I(\c0.n20927 ));
    Odrv4 I__12148 (
            .O(N__54158),
            .I(\c0.n20927 ));
    LocalMux I__12147 (
            .O(N__54155),
            .I(\c0.n20927 ));
    InMux I__12146 (
            .O(N__54148),
            .I(N__54145));
    LocalMux I__12145 (
            .O(N__54145),
            .I(N__54142));
    Odrv12 I__12144 (
            .O(N__54142),
            .I(\c0.n22119 ));
    CascadeMux I__12143 (
            .O(N__54139),
            .I(\c0.n21099_cascade_ ));
    InMux I__12142 (
            .O(N__54136),
            .I(N__54132));
    InMux I__12141 (
            .O(N__54135),
            .I(N__54127));
    LocalMux I__12140 (
            .O(N__54132),
            .I(N__54124));
    InMux I__12139 (
            .O(N__54131),
            .I(N__54119));
    InMux I__12138 (
            .O(N__54130),
            .I(N__54119));
    LocalMux I__12137 (
            .O(N__54127),
            .I(\c0.n21160 ));
    Odrv4 I__12136 (
            .O(N__54124),
            .I(\c0.n21160 ));
    LocalMux I__12135 (
            .O(N__54119),
            .I(\c0.n21160 ));
    InMux I__12134 (
            .O(N__54112),
            .I(N__54108));
    InMux I__12133 (
            .O(N__54111),
            .I(N__54105));
    LocalMux I__12132 (
            .O(N__54108),
            .I(N__54100));
    LocalMux I__12131 (
            .O(N__54105),
            .I(N__54100));
    Odrv4 I__12130 (
            .O(N__54100),
            .I(\c0.data_in_frame_29_6 ));
    InMux I__12129 (
            .O(N__54097),
            .I(N__54094));
    LocalMux I__12128 (
            .O(N__54094),
            .I(N__54090));
    InMux I__12127 (
            .O(N__54093),
            .I(N__54087));
    Span4Mux_h I__12126 (
            .O(N__54090),
            .I(N__54084));
    LocalMux I__12125 (
            .O(N__54087),
            .I(\c0.n63_adj_4293 ));
    Odrv4 I__12124 (
            .O(N__54084),
            .I(\c0.n63_adj_4293 ));
    CascadeMux I__12123 (
            .O(N__54079),
            .I(\c0.n22148_cascade_ ));
    InMux I__12122 (
            .O(N__54076),
            .I(N__54073));
    LocalMux I__12121 (
            .O(N__54073),
            .I(\c0.n21233 ));
    InMux I__12120 (
            .O(N__54070),
            .I(N__54067));
    LocalMux I__12119 (
            .O(N__54067),
            .I(N__54064));
    Span4Mux_h I__12118 (
            .O(N__54064),
            .I(N__54061));
    Odrv4 I__12117 (
            .O(N__54061),
            .I(\c0.n26_adj_4294 ));
    CascadeMux I__12116 (
            .O(N__54058),
            .I(\c0.rx.n12862_cascade_ ));
    InMux I__12115 (
            .O(N__54055),
            .I(N__54051));
    InMux I__12114 (
            .O(N__54054),
            .I(N__54048));
    LocalMux I__12113 (
            .O(N__54051),
            .I(\c0.rx.r_Clock_Count_7 ));
    LocalMux I__12112 (
            .O(N__54048),
            .I(\c0.rx.r_Clock_Count_7 ));
    InMux I__12111 (
            .O(N__54043),
            .I(N__54039));
    InMux I__12110 (
            .O(N__54042),
            .I(N__54036));
    LocalMux I__12109 (
            .O(N__54039),
            .I(\c0.rx.r_Clock_Count_5 ));
    LocalMux I__12108 (
            .O(N__54036),
            .I(\c0.rx.r_Clock_Count_5 ));
    InMux I__12107 (
            .O(N__54031),
            .I(N__54027));
    InMux I__12106 (
            .O(N__54030),
            .I(N__54024));
    LocalMux I__12105 (
            .O(N__54027),
            .I(\c0.rx.r_Clock_Count_6 ));
    LocalMux I__12104 (
            .O(N__54024),
            .I(\c0.rx.r_Clock_Count_6 ));
    CascadeMux I__12103 (
            .O(N__54019),
            .I(\c0.rx.n80_cascade_ ));
    InMux I__12102 (
            .O(N__54016),
            .I(N__54012));
    InMux I__12101 (
            .O(N__54015),
            .I(N__54009));
    LocalMux I__12100 (
            .O(N__54012),
            .I(N__54004));
    LocalMux I__12099 (
            .O(N__54009),
            .I(N__54001));
    InMux I__12098 (
            .O(N__54008),
            .I(N__53998));
    InMux I__12097 (
            .O(N__54007),
            .I(N__53995));
    Odrv4 I__12096 (
            .O(N__54004),
            .I(\c0.n13761 ));
    Odrv4 I__12095 (
            .O(N__54001),
            .I(\c0.n13761 ));
    LocalMux I__12094 (
            .O(N__53998),
            .I(\c0.n13761 ));
    LocalMux I__12093 (
            .O(N__53995),
            .I(\c0.n13761 ));
    InMux I__12092 (
            .O(N__53986),
            .I(N__53983));
    LocalMux I__12091 (
            .O(N__53983),
            .I(\c0.n22145 ));
    InMux I__12090 (
            .O(N__53980),
            .I(N__53976));
    InMux I__12089 (
            .O(N__53979),
            .I(N__53973));
    LocalMux I__12088 (
            .O(N__53976),
            .I(\c0.n21949 ));
    LocalMux I__12087 (
            .O(N__53973),
            .I(\c0.n21949 ));
    CascadeMux I__12086 (
            .O(N__53968),
            .I(\c0.n22145_cascade_ ));
    InMux I__12085 (
            .O(N__53965),
            .I(N__53962));
    LocalMux I__12084 (
            .O(N__53962),
            .I(\c0.n10_adj_4297 ));
    CascadeMux I__12083 (
            .O(N__53959),
            .I(\c0.n23335_cascade_ ));
    CascadeMux I__12082 (
            .O(N__53956),
            .I(N__53953));
    InMux I__12081 (
            .O(N__53953),
            .I(N__53950));
    LocalMux I__12080 (
            .O(N__53950),
            .I(N__53947));
    Span4Mux_v I__12079 (
            .O(N__53947),
            .I(N__53944));
    Odrv4 I__12078 (
            .O(N__53944),
            .I(\c0.n21_adj_4300 ));
    CascadeMux I__12077 (
            .O(N__53941),
            .I(N__53937));
    CascadeMux I__12076 (
            .O(N__53940),
            .I(N__53934));
    InMux I__12075 (
            .O(N__53937),
            .I(N__53931));
    InMux I__12074 (
            .O(N__53934),
            .I(N__53928));
    LocalMux I__12073 (
            .O(N__53931),
            .I(N__53925));
    LocalMux I__12072 (
            .O(N__53928),
            .I(\c0.data_in_frame_29_3 ));
    Odrv4 I__12071 (
            .O(N__53925),
            .I(\c0.data_in_frame_29_3 ));
    CascadeMux I__12070 (
            .O(N__53920),
            .I(N__53917));
    InMux I__12069 (
            .O(N__53917),
            .I(N__53913));
    InMux I__12068 (
            .O(N__53916),
            .I(N__53910));
    LocalMux I__12067 (
            .O(N__53913),
            .I(\c0.data_in_frame_28_0 ));
    LocalMux I__12066 (
            .O(N__53910),
            .I(\c0.data_in_frame_28_0 ));
    InMux I__12065 (
            .O(N__53905),
            .I(N__53902));
    LocalMux I__12064 (
            .O(N__53902),
            .I(N__53898));
    InMux I__12063 (
            .O(N__53901),
            .I(N__53895));
    Span4Mux_v I__12062 (
            .O(N__53898),
            .I(N__53892));
    LocalMux I__12061 (
            .O(N__53895),
            .I(N__53889));
    Span4Mux_h I__12060 (
            .O(N__53892),
            .I(N__53886));
    Span4Mux_h I__12059 (
            .O(N__53889),
            .I(N__53883));
    Span4Mux_v I__12058 (
            .O(N__53886),
            .I(N__53880));
    Span4Mux_v I__12057 (
            .O(N__53883),
            .I(N__53877));
    Span4Mux_v I__12056 (
            .O(N__53880),
            .I(N__53874));
    Span4Mux_v I__12055 (
            .O(N__53877),
            .I(N__53871));
    Odrv4 I__12054 (
            .O(N__53874),
            .I(\c0.n6404 ));
    Odrv4 I__12053 (
            .O(N__53871),
            .I(\c0.n6404 ));
    InMux I__12052 (
            .O(N__53866),
            .I(N__53863));
    LocalMux I__12051 (
            .O(N__53863),
            .I(N__53859));
    InMux I__12050 (
            .O(N__53862),
            .I(N__53856));
    Span12Mux_v I__12049 (
            .O(N__53859),
            .I(N__53851));
    LocalMux I__12048 (
            .O(N__53856),
            .I(N__53851));
    Odrv12 I__12047 (
            .O(N__53851),
            .I(\c0.n21834 ));
    InMux I__12046 (
            .O(N__53848),
            .I(N__53845));
    LocalMux I__12045 (
            .O(N__53845),
            .I(N__53842));
    Odrv4 I__12044 (
            .O(N__53842),
            .I(\c0.n22040 ));
    CascadeMux I__12043 (
            .O(N__53839),
            .I(\c0.n22040_cascade_ ));
    InMux I__12042 (
            .O(N__53836),
            .I(N__53833));
    LocalMux I__12041 (
            .O(N__53833),
            .I(N__53830));
    Odrv4 I__12040 (
            .O(N__53830),
            .I(\c0.n21208 ));
    InMux I__12039 (
            .O(N__53827),
            .I(N__53824));
    LocalMux I__12038 (
            .O(N__53824),
            .I(\c0.n21099 ));
    CascadeMux I__12037 (
            .O(N__53821),
            .I(\c0.n6_adj_4219_cascade_ ));
    CascadeMux I__12036 (
            .O(N__53818),
            .I(N__53814));
    InMux I__12035 (
            .O(N__53817),
            .I(N__53811));
    InMux I__12034 (
            .O(N__53814),
            .I(N__53806));
    LocalMux I__12033 (
            .O(N__53811),
            .I(N__53803));
    InMux I__12032 (
            .O(N__53810),
            .I(N__53800));
    InMux I__12031 (
            .O(N__53809),
            .I(N__53797));
    LocalMux I__12030 (
            .O(N__53806),
            .I(\c0.data_in_frame_21_2 ));
    Odrv4 I__12029 (
            .O(N__53803),
            .I(\c0.data_in_frame_21_2 ));
    LocalMux I__12028 (
            .O(N__53800),
            .I(\c0.data_in_frame_21_2 ));
    LocalMux I__12027 (
            .O(N__53797),
            .I(\c0.data_in_frame_21_2 ));
    InMux I__12026 (
            .O(N__53788),
            .I(N__53783));
    InMux I__12025 (
            .O(N__53787),
            .I(N__53780));
    InMux I__12024 (
            .O(N__53786),
            .I(N__53777));
    LocalMux I__12023 (
            .O(N__53783),
            .I(\c0.n22197 ));
    LocalMux I__12022 (
            .O(N__53780),
            .I(\c0.n22197 ));
    LocalMux I__12021 (
            .O(N__53777),
            .I(\c0.n22197 ));
    CascadeMux I__12020 (
            .O(N__53770),
            .I(\c0.n21949_cascade_ ));
    InMux I__12019 (
            .O(N__53767),
            .I(N__53763));
    CascadeMux I__12018 (
            .O(N__53766),
            .I(N__53759));
    LocalMux I__12017 (
            .O(N__53763),
            .I(N__53756));
    InMux I__12016 (
            .O(N__53762),
            .I(N__53751));
    InMux I__12015 (
            .O(N__53759),
            .I(N__53751));
    Odrv4 I__12014 (
            .O(N__53756),
            .I(\c0.n20137 ));
    LocalMux I__12013 (
            .O(N__53751),
            .I(\c0.n20137 ));
    CascadeMux I__12012 (
            .O(N__53746),
            .I(\c0.n22157_cascade_ ));
    InMux I__12011 (
            .O(N__53743),
            .I(N__53740));
    LocalMux I__12010 (
            .O(N__53740),
            .I(N__53737));
    Span4Mux_h I__12009 (
            .O(N__53737),
            .I(N__53734));
    Odrv4 I__12008 (
            .O(N__53734),
            .I(\c0.n20846 ));
    CascadeMux I__12007 (
            .O(N__53731),
            .I(\c0.n20846_cascade_ ));
    InMux I__12006 (
            .O(N__53728),
            .I(N__53724));
    CascadeMux I__12005 (
            .O(N__53727),
            .I(N__53721));
    LocalMux I__12004 (
            .O(N__53724),
            .I(N__53716));
    InMux I__12003 (
            .O(N__53721),
            .I(N__53713));
    InMux I__12002 (
            .O(N__53720),
            .I(N__53710));
    InMux I__12001 (
            .O(N__53719),
            .I(N__53707));
    Sp12to4 I__12000 (
            .O(N__53716),
            .I(N__53700));
    LocalMux I__11999 (
            .O(N__53713),
            .I(N__53700));
    LocalMux I__11998 (
            .O(N__53710),
            .I(N__53700));
    LocalMux I__11997 (
            .O(N__53707),
            .I(\c0.data_in_frame_25_4 ));
    Odrv12 I__11996 (
            .O(N__53700),
            .I(\c0.data_in_frame_25_4 ));
    InMux I__11995 (
            .O(N__53695),
            .I(N__53691));
    CascadeMux I__11994 (
            .O(N__53694),
            .I(N__53686));
    LocalMux I__11993 (
            .O(N__53691),
            .I(N__53683));
    InMux I__11992 (
            .O(N__53690),
            .I(N__53678));
    InMux I__11991 (
            .O(N__53689),
            .I(N__53678));
    InMux I__11990 (
            .O(N__53686),
            .I(N__53675));
    Span4Mux_h I__11989 (
            .O(N__53683),
            .I(N__53672));
    LocalMux I__11988 (
            .O(N__53678),
            .I(N__53669));
    LocalMux I__11987 (
            .O(N__53675),
            .I(N__53664));
    Span4Mux_v I__11986 (
            .O(N__53672),
            .I(N__53664));
    Span4Mux_h I__11985 (
            .O(N__53669),
            .I(N__53661));
    Odrv4 I__11984 (
            .O(N__53664),
            .I(\c0.data_in_frame_25_2 ));
    Odrv4 I__11983 (
            .O(N__53661),
            .I(\c0.data_in_frame_25_2 ));
    InMux I__11982 (
            .O(N__53656),
            .I(N__53651));
    CascadeMux I__11981 (
            .O(N__53655),
            .I(N__53647));
    InMux I__11980 (
            .O(N__53654),
            .I(N__53644));
    LocalMux I__11979 (
            .O(N__53651),
            .I(N__53641));
    InMux I__11978 (
            .O(N__53650),
            .I(N__53636));
    InMux I__11977 (
            .O(N__53647),
            .I(N__53636));
    LocalMux I__11976 (
            .O(N__53644),
            .I(N__53633));
    Span4Mux_v I__11975 (
            .O(N__53641),
            .I(N__53630));
    LocalMux I__11974 (
            .O(N__53636),
            .I(N__53627));
    Span4Mux_h I__11973 (
            .O(N__53633),
            .I(N__53623));
    Span4Mux_h I__11972 (
            .O(N__53630),
            .I(N__53618));
    Span4Mux_h I__11971 (
            .O(N__53627),
            .I(N__53618));
    InMux I__11970 (
            .O(N__53626),
            .I(N__53615));
    Span4Mux_v I__11969 (
            .O(N__53623),
            .I(N__53612));
    Span4Mux_v I__11968 (
            .O(N__53618),
            .I(N__53609));
    LocalMux I__11967 (
            .O(N__53615),
            .I(\c0.data_in_frame_25_3 ));
    Odrv4 I__11966 (
            .O(N__53612),
            .I(\c0.data_in_frame_25_3 ));
    Odrv4 I__11965 (
            .O(N__53609),
            .I(\c0.data_in_frame_25_3 ));
    InMux I__11964 (
            .O(N__53602),
            .I(N__53595));
    InMux I__11963 (
            .O(N__53601),
            .I(N__53590));
    InMux I__11962 (
            .O(N__53600),
            .I(N__53590));
    InMux I__11961 (
            .O(N__53599),
            .I(N__53587));
    CascadeMux I__11960 (
            .O(N__53598),
            .I(N__53584));
    LocalMux I__11959 (
            .O(N__53595),
            .I(N__53581));
    LocalMux I__11958 (
            .O(N__53590),
            .I(N__53576));
    LocalMux I__11957 (
            .O(N__53587),
            .I(N__53576));
    InMux I__11956 (
            .O(N__53584),
            .I(N__53573));
    Span4Mux_h I__11955 (
            .O(N__53581),
            .I(N__53570));
    Span4Mux_h I__11954 (
            .O(N__53576),
            .I(N__53567));
    LocalMux I__11953 (
            .O(N__53573),
            .I(\c0.data_in_frame_25_5 ));
    Odrv4 I__11952 (
            .O(N__53570),
            .I(\c0.data_in_frame_25_5 ));
    Odrv4 I__11951 (
            .O(N__53567),
            .I(\c0.data_in_frame_25_5 ));
    InMux I__11950 (
            .O(N__53560),
            .I(N__53557));
    LocalMux I__11949 (
            .O(N__53557),
            .I(N__53554));
    Span4Mux_h I__11948 (
            .O(N__53554),
            .I(N__53551));
    Odrv4 I__11947 (
            .O(N__53551),
            .I(\c0.n22370 ));
    InMux I__11946 (
            .O(N__53548),
            .I(N__53545));
    LocalMux I__11945 (
            .O(N__53545),
            .I(\c0.n12_adj_4491 ));
    InMux I__11944 (
            .O(N__53542),
            .I(N__53539));
    LocalMux I__11943 (
            .O(N__53539),
            .I(\c0.n23009 ));
    CascadeMux I__11942 (
            .O(N__53536),
            .I(\c0.n22370_cascade_ ));
    CascadeMux I__11941 (
            .O(N__53533),
            .I(N__53529));
    InMux I__11940 (
            .O(N__53532),
            .I(N__53524));
    InMux I__11939 (
            .O(N__53529),
            .I(N__53524));
    LocalMux I__11938 (
            .O(N__53524),
            .I(N__53521));
    Odrv4 I__11937 (
            .O(N__53521),
            .I(\c0.n23356 ));
    SRMux I__11936 (
            .O(N__53518),
            .I(N__53515));
    LocalMux I__11935 (
            .O(N__53515),
            .I(N__53512));
    Span4Mux_h I__11934 (
            .O(N__53512),
            .I(N__53509));
    Span4Mux_h I__11933 (
            .O(N__53509),
            .I(N__53506));
    Odrv4 I__11932 (
            .O(N__53506),
            .I(\c0.n21366 ));
    InMux I__11931 (
            .O(N__53503),
            .I(N__53499));
    InMux I__11930 (
            .O(N__53502),
            .I(N__53496));
    LocalMux I__11929 (
            .O(N__53499),
            .I(N__53493));
    LocalMux I__11928 (
            .O(N__53496),
            .I(N__53490));
    Span4Mux_h I__11927 (
            .O(N__53493),
            .I(N__53487));
    Span4Mux_v I__11926 (
            .O(N__53490),
            .I(N__53482));
    Span4Mux_v I__11925 (
            .O(N__53487),
            .I(N__53482));
    Span4Mux_h I__11924 (
            .O(N__53482),
            .I(N__53479));
    Odrv4 I__11923 (
            .O(N__53479),
            .I(\c0.n21855 ));
    CascadeMux I__11922 (
            .O(N__53476),
            .I(N__53472));
    InMux I__11921 (
            .O(N__53475),
            .I(N__53469));
    InMux I__11920 (
            .O(N__53472),
            .I(N__53466));
    LocalMux I__11919 (
            .O(N__53469),
            .I(N__53461));
    LocalMux I__11918 (
            .O(N__53466),
            .I(N__53458));
    InMux I__11917 (
            .O(N__53465),
            .I(N__53452));
    InMux I__11916 (
            .O(N__53464),
            .I(N__53452));
    Span4Mux_h I__11915 (
            .O(N__53461),
            .I(N__53449));
    Span4Mux_h I__11914 (
            .O(N__53458),
            .I(N__53445));
    InMux I__11913 (
            .O(N__53457),
            .I(N__53442));
    LocalMux I__11912 (
            .O(N__53452),
            .I(N__53437));
    Span4Mux_h I__11911 (
            .O(N__53449),
            .I(N__53437));
    InMux I__11910 (
            .O(N__53448),
            .I(N__53433));
    Span4Mux_v I__11909 (
            .O(N__53445),
            .I(N__53426));
    LocalMux I__11908 (
            .O(N__53442),
            .I(N__53426));
    Span4Mux_v I__11907 (
            .O(N__53437),
            .I(N__53426));
    InMux I__11906 (
            .O(N__53436),
            .I(N__53423));
    LocalMux I__11905 (
            .O(N__53433),
            .I(encoder0_position_2));
    Odrv4 I__11904 (
            .O(N__53426),
            .I(encoder0_position_2));
    LocalMux I__11903 (
            .O(N__53423),
            .I(encoder0_position_2));
    InMux I__11902 (
            .O(N__53416),
            .I(N__53413));
    LocalMux I__11901 (
            .O(N__53413),
            .I(N__53410));
    Span4Mux_h I__11900 (
            .O(N__53410),
            .I(N__53406));
    InMux I__11899 (
            .O(N__53409),
            .I(N__53403));
    Span4Mux_h I__11898 (
            .O(N__53406),
            .I(N__53400));
    LocalMux I__11897 (
            .O(N__53403),
            .I(N__53397));
    Odrv4 I__11896 (
            .O(N__53400),
            .I(\c0.n22248 ));
    Odrv4 I__11895 (
            .O(N__53397),
            .I(\c0.n22248 ));
    InMux I__11894 (
            .O(N__53392),
            .I(N__53389));
    LocalMux I__11893 (
            .O(N__53389),
            .I(N__53383));
    InMux I__11892 (
            .O(N__53388),
            .I(N__53380));
    InMux I__11891 (
            .O(N__53387),
            .I(N__53375));
    InMux I__11890 (
            .O(N__53386),
            .I(N__53375));
    Span4Mux_h I__11889 (
            .O(N__53383),
            .I(N__53372));
    LocalMux I__11888 (
            .O(N__53380),
            .I(N__53369));
    LocalMux I__11887 (
            .O(N__53375),
            .I(N__53365));
    Span4Mux_v I__11886 (
            .O(N__53372),
            .I(N__53360));
    Span4Mux_h I__11885 (
            .O(N__53369),
            .I(N__53360));
    InMux I__11884 (
            .O(N__53368),
            .I(N__53357));
    Span4Mux_h I__11883 (
            .O(N__53365),
            .I(N__53354));
    Span4Mux_h I__11882 (
            .O(N__53360),
            .I(N__53351));
    LocalMux I__11881 (
            .O(N__53357),
            .I(N__53346));
    Sp12to4 I__11880 (
            .O(N__53354),
            .I(N__53346));
    Span4Mux_v I__11879 (
            .O(N__53351),
            .I(N__53343));
    Span12Mux_v I__11878 (
            .O(N__53346),
            .I(N__53340));
    Odrv4 I__11877 (
            .O(N__53343),
            .I(\c0.n13379 ));
    Odrv12 I__11876 (
            .O(N__53340),
            .I(\c0.n13379 ));
    CascadeMux I__11875 (
            .O(N__53335),
            .I(N__53332));
    InMux I__11874 (
            .O(N__53332),
            .I(N__53329));
    LocalMux I__11873 (
            .O(N__53329),
            .I(N__53325));
    InMux I__11872 (
            .O(N__53328),
            .I(N__53322));
    Span4Mux_v I__11871 (
            .O(N__53325),
            .I(N__53318));
    LocalMux I__11870 (
            .O(N__53322),
            .I(N__53315));
    InMux I__11869 (
            .O(N__53321),
            .I(N__53312));
    Span4Mux_h I__11868 (
            .O(N__53318),
            .I(N__53307));
    Span4Mux_v I__11867 (
            .O(N__53315),
            .I(N__53307));
    LocalMux I__11866 (
            .O(N__53312),
            .I(\c0.data_in_frame_20_7 ));
    Odrv4 I__11865 (
            .O(N__53307),
            .I(\c0.data_in_frame_20_7 ));
    CascadeMux I__11864 (
            .O(N__53302),
            .I(\c0.n28_cascade_ ));
    CascadeMux I__11863 (
            .O(N__53299),
            .I(\c0.n23640_cascade_ ));
    CascadeMux I__11862 (
            .O(N__53296),
            .I(\c0.n22305_cascade_ ));
    InMux I__11861 (
            .O(N__53293),
            .I(N__53287));
    InMux I__11860 (
            .O(N__53292),
            .I(N__53287));
    LocalMux I__11859 (
            .O(N__53287),
            .I(N__53283));
    InMux I__11858 (
            .O(N__53286),
            .I(N__53280));
    Span4Mux_v I__11857 (
            .O(N__53283),
            .I(N__53274));
    LocalMux I__11856 (
            .O(N__53280),
            .I(N__53274));
    CascadeMux I__11855 (
            .O(N__53279),
            .I(N__53271));
    Span4Mux_h I__11854 (
            .O(N__53274),
            .I(N__53268));
    InMux I__11853 (
            .O(N__53271),
            .I(N__53265));
    Span4Mux_h I__11852 (
            .O(N__53268),
            .I(N__53262));
    LocalMux I__11851 (
            .O(N__53265),
            .I(\c0.data_in_frame_21_1 ));
    Odrv4 I__11850 (
            .O(N__53262),
            .I(\c0.data_in_frame_21_1 ));
    InMux I__11849 (
            .O(N__53257),
            .I(N__53251));
    InMux I__11848 (
            .O(N__53256),
            .I(N__53251));
    LocalMux I__11847 (
            .O(N__53251),
            .I(\c0.n23640 ));
    InMux I__11846 (
            .O(N__53248),
            .I(N__53245));
    LocalMux I__11845 (
            .O(N__53245),
            .I(\c0.n22305 ));
    InMux I__11844 (
            .O(N__53242),
            .I(N__53238));
    InMux I__11843 (
            .O(N__53241),
            .I(N__53235));
    LocalMux I__11842 (
            .O(N__53238),
            .I(N__53232));
    LocalMux I__11841 (
            .O(N__53235),
            .I(\c0.data_in_frame_20_1 ));
    Odrv4 I__11840 (
            .O(N__53232),
            .I(\c0.data_in_frame_20_1 ));
    CascadeMux I__11839 (
            .O(N__53227),
            .I(\c0.n6_adj_4226_cascade_ ));
    CascadeMux I__11838 (
            .O(N__53224),
            .I(\c0.n23615_cascade_ ));
    CascadeMux I__11837 (
            .O(N__53221),
            .I(\c0.n22100_cascade_ ));
    InMux I__11836 (
            .O(N__53218),
            .I(N__53214));
    InMux I__11835 (
            .O(N__53217),
            .I(N__53211));
    LocalMux I__11834 (
            .O(N__53214),
            .I(\c0.n22081 ));
    LocalMux I__11833 (
            .O(N__53211),
            .I(\c0.n22081 ));
    CascadeMux I__11832 (
            .O(N__53206),
            .I(N__53203));
    InMux I__11831 (
            .O(N__53203),
            .I(N__53200));
    LocalMux I__11830 (
            .O(N__53200),
            .I(\c0.n6_adj_4224 ));
    InMux I__11829 (
            .O(N__53197),
            .I(N__53190));
    InMux I__11828 (
            .O(N__53196),
            .I(N__53185));
    InMux I__11827 (
            .O(N__53195),
            .I(N__53182));
    InMux I__11826 (
            .O(N__53194),
            .I(N__53178));
    InMux I__11825 (
            .O(N__53193),
            .I(N__53171));
    LocalMux I__11824 (
            .O(N__53190),
            .I(N__53165));
    InMux I__11823 (
            .O(N__53189),
            .I(N__53162));
    InMux I__11822 (
            .O(N__53188),
            .I(N__53159));
    LocalMux I__11821 (
            .O(N__53185),
            .I(N__53156));
    LocalMux I__11820 (
            .O(N__53182),
            .I(N__53153));
    InMux I__11819 (
            .O(N__53181),
            .I(N__53150));
    LocalMux I__11818 (
            .O(N__53178),
            .I(N__53147));
    InMux I__11817 (
            .O(N__53177),
            .I(N__53144));
    InMux I__11816 (
            .O(N__53176),
            .I(N__53141));
    InMux I__11815 (
            .O(N__53175),
            .I(N__53138));
    CascadeMux I__11814 (
            .O(N__53174),
            .I(N__53132));
    LocalMux I__11813 (
            .O(N__53171),
            .I(N__53125));
    InMux I__11812 (
            .O(N__53170),
            .I(N__53120));
    InMux I__11811 (
            .O(N__53169),
            .I(N__53120));
    CascadeMux I__11810 (
            .O(N__53168),
            .I(N__53117));
    Span4Mux_v I__11809 (
            .O(N__53165),
            .I(N__53110));
    LocalMux I__11808 (
            .O(N__53162),
            .I(N__53110));
    LocalMux I__11807 (
            .O(N__53159),
            .I(N__53105));
    Span4Mux_v I__11806 (
            .O(N__53156),
            .I(N__53105));
    Span4Mux_v I__11805 (
            .O(N__53153),
            .I(N__53098));
    LocalMux I__11804 (
            .O(N__53150),
            .I(N__53098));
    Span4Mux_v I__11803 (
            .O(N__53147),
            .I(N__53098));
    LocalMux I__11802 (
            .O(N__53144),
            .I(N__53093));
    LocalMux I__11801 (
            .O(N__53141),
            .I(N__53093));
    LocalMux I__11800 (
            .O(N__53138),
            .I(N__53090));
    InMux I__11799 (
            .O(N__53137),
            .I(N__53087));
    InMux I__11798 (
            .O(N__53136),
            .I(N__53084));
    InMux I__11797 (
            .O(N__53135),
            .I(N__53077));
    InMux I__11796 (
            .O(N__53132),
            .I(N__53077));
    InMux I__11795 (
            .O(N__53131),
            .I(N__53077));
    InMux I__11794 (
            .O(N__53130),
            .I(N__53070));
    InMux I__11793 (
            .O(N__53129),
            .I(N__53070));
    InMux I__11792 (
            .O(N__53128),
            .I(N__53070));
    Span4Mux_v I__11791 (
            .O(N__53125),
            .I(N__53065));
    LocalMux I__11790 (
            .O(N__53120),
            .I(N__53065));
    InMux I__11789 (
            .O(N__53117),
            .I(N__53058));
    InMux I__11788 (
            .O(N__53116),
            .I(N__53058));
    InMux I__11787 (
            .O(N__53115),
            .I(N__53058));
    Span4Mux_h I__11786 (
            .O(N__53110),
            .I(N__53053));
    Span4Mux_h I__11785 (
            .O(N__53105),
            .I(N__53053));
    Span4Mux_h I__11784 (
            .O(N__53098),
            .I(N__53046));
    Span4Mux_v I__11783 (
            .O(N__53093),
            .I(N__53046));
    Span4Mux_h I__11782 (
            .O(N__53090),
            .I(N__53046));
    LocalMux I__11781 (
            .O(N__53087),
            .I(\c0.n21737 ));
    LocalMux I__11780 (
            .O(N__53084),
            .I(\c0.n21737 ));
    LocalMux I__11779 (
            .O(N__53077),
            .I(\c0.n21737 ));
    LocalMux I__11778 (
            .O(N__53070),
            .I(\c0.n21737 ));
    Odrv4 I__11777 (
            .O(N__53065),
            .I(\c0.n21737 ));
    LocalMux I__11776 (
            .O(N__53058),
            .I(\c0.n21737 ));
    Odrv4 I__11775 (
            .O(N__53053),
            .I(\c0.n21737 ));
    Odrv4 I__11774 (
            .O(N__53046),
            .I(\c0.n21737 ));
    InMux I__11773 (
            .O(N__53029),
            .I(N__53023));
    InMux I__11772 (
            .O(N__53028),
            .I(N__53016));
    InMux I__11771 (
            .O(N__53027),
            .I(N__53013));
    InMux I__11770 (
            .O(N__53026),
            .I(N__53006));
    LocalMux I__11769 (
            .O(N__53023),
            .I(N__53003));
    InMux I__11768 (
            .O(N__53022),
            .I(N__53000));
    InMux I__11767 (
            .O(N__53021),
            .I(N__52993));
    InMux I__11766 (
            .O(N__53020),
            .I(N__52993));
    InMux I__11765 (
            .O(N__53019),
            .I(N__52993));
    LocalMux I__11764 (
            .O(N__53016),
            .I(N__52988));
    LocalMux I__11763 (
            .O(N__53013),
            .I(N__52988));
    InMux I__11762 (
            .O(N__53012),
            .I(N__52985));
    InMux I__11761 (
            .O(N__53011),
            .I(N__52982));
    InMux I__11760 (
            .O(N__53010),
            .I(N__52978));
    InMux I__11759 (
            .O(N__53009),
            .I(N__52975));
    LocalMux I__11758 (
            .O(N__53006),
            .I(N__52967));
    Span4Mux_h I__11757 (
            .O(N__53003),
            .I(N__52964));
    LocalMux I__11756 (
            .O(N__53000),
            .I(N__52961));
    LocalMux I__11755 (
            .O(N__52993),
            .I(N__52958));
    Span4Mux_v I__11754 (
            .O(N__52988),
            .I(N__52951));
    LocalMux I__11753 (
            .O(N__52985),
            .I(N__52951));
    LocalMux I__11752 (
            .O(N__52982),
            .I(N__52951));
    InMux I__11751 (
            .O(N__52981),
            .I(N__52948));
    LocalMux I__11750 (
            .O(N__52978),
            .I(N__52942));
    LocalMux I__11749 (
            .O(N__52975),
            .I(N__52942));
    InMux I__11748 (
            .O(N__52974),
            .I(N__52939));
    InMux I__11747 (
            .O(N__52973),
            .I(N__52934));
    InMux I__11746 (
            .O(N__52972),
            .I(N__52934));
    InMux I__11745 (
            .O(N__52971),
            .I(N__52929));
    InMux I__11744 (
            .O(N__52970),
            .I(N__52929));
    Span4Mux_h I__11743 (
            .O(N__52967),
            .I(N__52924));
    Span4Mux_h I__11742 (
            .O(N__52964),
            .I(N__52924));
    Span4Mux_v I__11741 (
            .O(N__52961),
            .I(N__52919));
    Span4Mux_h I__11740 (
            .O(N__52958),
            .I(N__52919));
    Span4Mux_v I__11739 (
            .O(N__52951),
            .I(N__52914));
    LocalMux I__11738 (
            .O(N__52948),
            .I(N__52914));
    InMux I__11737 (
            .O(N__52947),
            .I(N__52911));
    Span4Mux_v I__11736 (
            .O(N__52942),
            .I(N__52902));
    LocalMux I__11735 (
            .O(N__52939),
            .I(N__52902));
    LocalMux I__11734 (
            .O(N__52934),
            .I(N__52902));
    LocalMux I__11733 (
            .O(N__52929),
            .I(N__52902));
    Odrv4 I__11732 (
            .O(N__52924),
            .I(\c0.n6_adj_4353 ));
    Odrv4 I__11731 (
            .O(N__52919),
            .I(\c0.n6_adj_4353 ));
    Odrv4 I__11730 (
            .O(N__52914),
            .I(\c0.n6_adj_4353 ));
    LocalMux I__11729 (
            .O(N__52911),
            .I(\c0.n6_adj_4353 ));
    Odrv4 I__11728 (
            .O(N__52902),
            .I(\c0.n6_adj_4353 ));
    InMux I__11727 (
            .O(N__52891),
            .I(N__52881));
    InMux I__11726 (
            .O(N__52890),
            .I(N__52878));
    InMux I__11725 (
            .O(N__52889),
            .I(N__52875));
    InMux I__11724 (
            .O(N__52888),
            .I(N__52864));
    InMux I__11723 (
            .O(N__52887),
            .I(N__52861));
    InMux I__11722 (
            .O(N__52886),
            .I(N__52855));
    InMux I__11721 (
            .O(N__52885),
            .I(N__52852));
    InMux I__11720 (
            .O(N__52884),
            .I(N__52849));
    LocalMux I__11719 (
            .O(N__52881),
            .I(N__52840));
    LocalMux I__11718 (
            .O(N__52878),
            .I(N__52837));
    LocalMux I__11717 (
            .O(N__52875),
            .I(N__52834));
    InMux I__11716 (
            .O(N__52874),
            .I(N__52831));
    InMux I__11715 (
            .O(N__52873),
            .I(N__52828));
    InMux I__11714 (
            .O(N__52872),
            .I(N__52825));
    InMux I__11713 (
            .O(N__52871),
            .I(N__52822));
    InMux I__11712 (
            .O(N__52870),
            .I(N__52819));
    InMux I__11711 (
            .O(N__52869),
            .I(N__52816));
    InMux I__11710 (
            .O(N__52868),
            .I(N__52812));
    InMux I__11709 (
            .O(N__52867),
            .I(N__52809));
    LocalMux I__11708 (
            .O(N__52864),
            .I(N__52804));
    LocalMux I__11707 (
            .O(N__52861),
            .I(N__52804));
    InMux I__11706 (
            .O(N__52860),
            .I(N__52801));
    InMux I__11705 (
            .O(N__52859),
            .I(N__52798));
    InMux I__11704 (
            .O(N__52858),
            .I(N__52795));
    LocalMux I__11703 (
            .O(N__52855),
            .I(N__52792));
    LocalMux I__11702 (
            .O(N__52852),
            .I(N__52787));
    LocalMux I__11701 (
            .O(N__52849),
            .I(N__52787));
    InMux I__11700 (
            .O(N__52848),
            .I(N__52784));
    InMux I__11699 (
            .O(N__52847),
            .I(N__52781));
    InMux I__11698 (
            .O(N__52846),
            .I(N__52778));
    InMux I__11697 (
            .O(N__52845),
            .I(N__52775));
    InMux I__11696 (
            .O(N__52844),
            .I(N__52772));
    InMux I__11695 (
            .O(N__52843),
            .I(N__52769));
    Span4Mux_h I__11694 (
            .O(N__52840),
            .I(N__52764));
    Span4Mux_v I__11693 (
            .O(N__52837),
            .I(N__52764));
    Span4Mux_v I__11692 (
            .O(N__52834),
            .I(N__52749));
    LocalMux I__11691 (
            .O(N__52831),
            .I(N__52749));
    LocalMux I__11690 (
            .O(N__52828),
            .I(N__52749));
    LocalMux I__11689 (
            .O(N__52825),
            .I(N__52749));
    LocalMux I__11688 (
            .O(N__52822),
            .I(N__52749));
    LocalMux I__11687 (
            .O(N__52819),
            .I(N__52749));
    LocalMux I__11686 (
            .O(N__52816),
            .I(N__52749));
    InMux I__11685 (
            .O(N__52815),
            .I(N__52746));
    LocalMux I__11684 (
            .O(N__52812),
            .I(N__52741));
    LocalMux I__11683 (
            .O(N__52809),
            .I(N__52738));
    Span4Mux_v I__11682 (
            .O(N__52804),
            .I(N__52731));
    LocalMux I__11681 (
            .O(N__52801),
            .I(N__52731));
    LocalMux I__11680 (
            .O(N__52798),
            .I(N__52731));
    LocalMux I__11679 (
            .O(N__52795),
            .I(N__52728));
    Span4Mux_v I__11678 (
            .O(N__52792),
            .I(N__52725));
    Span4Mux_h I__11677 (
            .O(N__52787),
            .I(N__52710));
    LocalMux I__11676 (
            .O(N__52784),
            .I(N__52710));
    LocalMux I__11675 (
            .O(N__52781),
            .I(N__52710));
    LocalMux I__11674 (
            .O(N__52778),
            .I(N__52710));
    LocalMux I__11673 (
            .O(N__52775),
            .I(N__52710));
    LocalMux I__11672 (
            .O(N__52772),
            .I(N__52710));
    LocalMux I__11671 (
            .O(N__52769),
            .I(N__52710));
    Span4Mux_h I__11670 (
            .O(N__52764),
            .I(N__52703));
    Span4Mux_v I__11669 (
            .O(N__52749),
            .I(N__52703));
    LocalMux I__11668 (
            .O(N__52746),
            .I(N__52703));
    InMux I__11667 (
            .O(N__52745),
            .I(N__52700));
    InMux I__11666 (
            .O(N__52744),
            .I(N__52697));
    Span12Mux_h I__11665 (
            .O(N__52741),
            .I(N__52694));
    Span4Mux_h I__11664 (
            .O(N__52738),
            .I(N__52691));
    Span4Mux_v I__11663 (
            .O(N__52731),
            .I(N__52686));
    Span4Mux_h I__11662 (
            .O(N__52728),
            .I(N__52686));
    Span4Mux_v I__11661 (
            .O(N__52725),
            .I(N__52679));
    Span4Mux_v I__11660 (
            .O(N__52710),
            .I(N__52679));
    Span4Mux_h I__11659 (
            .O(N__52703),
            .I(N__52679));
    LocalMux I__11658 (
            .O(N__52700),
            .I(N__52674));
    LocalMux I__11657 (
            .O(N__52697),
            .I(N__52674));
    Odrv12 I__11656 (
            .O(N__52694),
            .I(\c0.n5_adj_4342 ));
    Odrv4 I__11655 (
            .O(N__52691),
            .I(\c0.n5_adj_4342 ));
    Odrv4 I__11654 (
            .O(N__52686),
            .I(\c0.n5_adj_4342 ));
    Odrv4 I__11653 (
            .O(N__52679),
            .I(\c0.n5_adj_4342 ));
    Odrv12 I__11652 (
            .O(N__52674),
            .I(\c0.n5_adj_4342 ));
    CascadeMux I__11651 (
            .O(N__52663),
            .I(N__52660));
    InMux I__11650 (
            .O(N__52660),
            .I(N__52654));
    InMux I__11649 (
            .O(N__52659),
            .I(N__52654));
    LocalMux I__11648 (
            .O(N__52654),
            .I(N__52651));
    Span4Mux_h I__11647 (
            .O(N__52651),
            .I(N__52646));
    InMux I__11646 (
            .O(N__52650),
            .I(N__52641));
    InMux I__11645 (
            .O(N__52649),
            .I(N__52641));
    Span4Mux_v I__11644 (
            .O(N__52646),
            .I(N__52638));
    LocalMux I__11643 (
            .O(N__52641),
            .I(\c0.FRAME_MATCHER_state_20 ));
    Odrv4 I__11642 (
            .O(N__52638),
            .I(\c0.FRAME_MATCHER_state_20 ));
    InMux I__11641 (
            .O(N__52633),
            .I(N__52630));
    LocalMux I__11640 (
            .O(N__52630),
            .I(N__52626));
    InMux I__11639 (
            .O(N__52629),
            .I(N__52623));
    Span4Mux_v I__11638 (
            .O(N__52626),
            .I(N__52618));
    LocalMux I__11637 (
            .O(N__52623),
            .I(N__52618));
    Span4Mux_h I__11636 (
            .O(N__52618),
            .I(N__52615));
    Odrv4 I__11635 (
            .O(N__52615),
            .I(\c0.n13190 ));
    CascadeMux I__11634 (
            .O(N__52612),
            .I(\c0.n18_adj_4222_cascade_ ));
    InMux I__11633 (
            .O(N__52609),
            .I(N__52605));
    InMux I__11632 (
            .O(N__52608),
            .I(N__52602));
    LocalMux I__11631 (
            .O(N__52605),
            .I(N__52597));
    LocalMux I__11630 (
            .O(N__52602),
            .I(N__52597));
    Span4Mux_v I__11629 (
            .O(N__52597),
            .I(N__52593));
    InMux I__11628 (
            .O(N__52596),
            .I(N__52590));
    Odrv4 I__11627 (
            .O(N__52593),
            .I(\c0.n22270 ));
    LocalMux I__11626 (
            .O(N__52590),
            .I(\c0.n22270 ));
    InMux I__11625 (
            .O(N__52585),
            .I(N__52582));
    LocalMux I__11624 (
            .O(N__52582),
            .I(N__52579));
    Odrv12 I__11623 (
            .O(N__52579),
            .I(\c0.n6_adj_4221 ));
    InMux I__11622 (
            .O(N__52576),
            .I(N__52573));
    LocalMux I__11621 (
            .O(N__52573),
            .I(N__52570));
    Span4Mux_h I__11620 (
            .O(N__52570),
            .I(N__52567));
    Odrv4 I__11619 (
            .O(N__52567),
            .I(\c0.n22308 ));
    CascadeMux I__11618 (
            .O(N__52564),
            .I(\c0.n22003_cascade_ ));
    InMux I__11617 (
            .O(N__52561),
            .I(N__52558));
    LocalMux I__11616 (
            .O(N__52558),
            .I(\c0.n5943 ));
    CascadeMux I__11615 (
            .O(N__52555),
            .I(\c0.n6221_cascade_ ));
    InMux I__11614 (
            .O(N__52552),
            .I(N__52549));
    LocalMux I__11613 (
            .O(N__52549),
            .I(\c0.n22003 ));
    InMux I__11612 (
            .O(N__52546),
            .I(N__52543));
    LocalMux I__11611 (
            .O(N__52543),
            .I(N__52540));
    Span4Mux_h I__11610 (
            .O(N__52540),
            .I(N__52536));
    InMux I__11609 (
            .O(N__52539),
            .I(N__52531));
    Span4Mux_v I__11608 (
            .O(N__52536),
            .I(N__52528));
    InMux I__11607 (
            .O(N__52535),
            .I(N__52525));
    InMux I__11606 (
            .O(N__52534),
            .I(N__52522));
    LocalMux I__11605 (
            .O(N__52531),
            .I(\c0.data_in_frame_10_2 ));
    Odrv4 I__11604 (
            .O(N__52528),
            .I(\c0.data_in_frame_10_2 ));
    LocalMux I__11603 (
            .O(N__52525),
            .I(\c0.data_in_frame_10_2 ));
    LocalMux I__11602 (
            .O(N__52522),
            .I(\c0.data_in_frame_10_2 ));
    CascadeMux I__11601 (
            .O(N__52513),
            .I(\c0.n20402_cascade_ ));
    InMux I__11600 (
            .O(N__52510),
            .I(N__52506));
    CascadeMux I__11599 (
            .O(N__52509),
            .I(N__52502));
    LocalMux I__11598 (
            .O(N__52506),
            .I(N__52499));
    InMux I__11597 (
            .O(N__52505),
            .I(N__52496));
    InMux I__11596 (
            .O(N__52502),
            .I(N__52493));
    Span4Mux_v I__11595 (
            .O(N__52499),
            .I(N__52490));
    LocalMux I__11594 (
            .O(N__52496),
            .I(N__52487));
    LocalMux I__11593 (
            .O(N__52493),
            .I(\c0.data_in_frame_9_6 ));
    Odrv4 I__11592 (
            .O(N__52490),
            .I(\c0.data_in_frame_9_6 ));
    Odrv4 I__11591 (
            .O(N__52487),
            .I(\c0.data_in_frame_9_6 ));
    CascadeMux I__11590 (
            .O(N__52480),
            .I(N__52477));
    InMux I__11589 (
            .O(N__52477),
            .I(N__52470));
    InMux I__11588 (
            .O(N__52476),
            .I(N__52470));
    InMux I__11587 (
            .O(N__52475),
            .I(N__52467));
    LocalMux I__11586 (
            .O(N__52470),
            .I(\c0.data_in_frame_9_4 ));
    LocalMux I__11585 (
            .O(N__52467),
            .I(\c0.data_in_frame_9_4 ));
    InMux I__11584 (
            .O(N__52462),
            .I(N__52456));
    InMux I__11583 (
            .O(N__52461),
            .I(N__52456));
    LocalMux I__11582 (
            .O(N__52456),
            .I(N__52453));
    Odrv4 I__11581 (
            .O(N__52453),
            .I(\c0.n21873 ));
    InMux I__11580 (
            .O(N__52450),
            .I(N__52447));
    LocalMux I__11579 (
            .O(N__52447),
            .I(N__52444));
    Span4Mux_v I__11578 (
            .O(N__52444),
            .I(N__52440));
    InMux I__11577 (
            .O(N__52443),
            .I(N__52437));
    Span4Mux_h I__11576 (
            .O(N__52440),
            .I(N__52432));
    LocalMux I__11575 (
            .O(N__52437),
            .I(N__52432));
    Span4Mux_h I__11574 (
            .O(N__52432),
            .I(N__52429));
    Odrv4 I__11573 (
            .O(N__52429),
            .I(\c0.n13287 ));
    InMux I__11572 (
            .O(N__52426),
            .I(N__52423));
    LocalMux I__11571 (
            .O(N__52423),
            .I(N__52420));
    Span4Mux_h I__11570 (
            .O(N__52420),
            .I(N__52417));
    Span4Mux_v I__11569 (
            .O(N__52417),
            .I(N__52414));
    Odrv4 I__11568 (
            .O(N__52414),
            .I(\c0.n22443 ));
    CascadeMux I__11567 (
            .O(N__52411),
            .I(\c0.n10_adj_4242_cascade_ ));
    InMux I__11566 (
            .O(N__52408),
            .I(N__52404));
    CascadeMux I__11565 (
            .O(N__52407),
            .I(N__52401));
    LocalMux I__11564 (
            .O(N__52404),
            .I(N__52398));
    InMux I__11563 (
            .O(N__52401),
            .I(N__52395));
    Span4Mux_h I__11562 (
            .O(N__52398),
            .I(N__52392));
    LocalMux I__11561 (
            .O(N__52395),
            .I(N__52386));
    Span4Mux_h I__11560 (
            .O(N__52392),
            .I(N__52386));
    InMux I__11559 (
            .O(N__52391),
            .I(N__52383));
    Odrv4 I__11558 (
            .O(N__52386),
            .I(\c0.data_in_frame_8_1 ));
    LocalMux I__11557 (
            .O(N__52383),
            .I(\c0.data_in_frame_8_1 ));
    InMux I__11556 (
            .O(N__52378),
            .I(N__52372));
    InMux I__11555 (
            .O(N__52377),
            .I(N__52367));
    InMux I__11554 (
            .O(N__52376),
            .I(N__52367));
    InMux I__11553 (
            .O(N__52375),
            .I(N__52364));
    LocalMux I__11552 (
            .O(N__52372),
            .I(N__52361));
    LocalMux I__11551 (
            .O(N__52367),
            .I(N__52358));
    LocalMux I__11550 (
            .O(N__52364),
            .I(\c0.data_in_frame_16_6 ));
    Odrv4 I__11549 (
            .O(N__52361),
            .I(\c0.data_in_frame_16_6 ));
    Odrv4 I__11548 (
            .O(N__52358),
            .I(\c0.data_in_frame_16_6 ));
    CascadeMux I__11547 (
            .O(N__52351),
            .I(\c0.n13786_cascade_ ));
    InMux I__11546 (
            .O(N__52348),
            .I(N__52345));
    LocalMux I__11545 (
            .O(N__52345),
            .I(N__52340));
    InMux I__11544 (
            .O(N__52344),
            .I(N__52335));
    InMux I__11543 (
            .O(N__52343),
            .I(N__52335));
    Odrv12 I__11542 (
            .O(N__52340),
            .I(\c0.n21170 ));
    LocalMux I__11541 (
            .O(N__52335),
            .I(\c0.n21170 ));
    InMux I__11540 (
            .O(N__52330),
            .I(N__52326));
    CascadeMux I__11539 (
            .O(N__52329),
            .I(N__52323));
    LocalMux I__11538 (
            .O(N__52326),
            .I(N__52320));
    InMux I__11537 (
            .O(N__52323),
            .I(N__52317));
    Span4Mux_h I__11536 (
            .O(N__52320),
            .I(N__52314));
    LocalMux I__11535 (
            .O(N__52317),
            .I(\c0.n13974 ));
    Odrv4 I__11534 (
            .O(N__52314),
            .I(\c0.n13974 ));
    InMux I__11533 (
            .O(N__52309),
            .I(N__52306));
    LocalMux I__11532 (
            .O(N__52306),
            .I(\c0.n22245 ));
    CascadeMux I__11531 (
            .O(N__52303),
            .I(N__52300));
    InMux I__11530 (
            .O(N__52300),
            .I(N__52297));
    LocalMux I__11529 (
            .O(N__52297),
            .I(N__52294));
    Odrv4 I__11528 (
            .O(N__52294),
            .I(\c0.n22379 ));
    CascadeMux I__11527 (
            .O(N__52291),
            .I(N__52288));
    InMux I__11526 (
            .O(N__52288),
            .I(N__52285));
    LocalMux I__11525 (
            .O(N__52285),
            .I(\c0.n38_adj_4260 ));
    InMux I__11524 (
            .O(N__52282),
            .I(N__52279));
    LocalMux I__11523 (
            .O(N__52279),
            .I(\c0.n6_adj_4256 ));
    InMux I__11522 (
            .O(N__52276),
            .I(N__52271));
    CascadeMux I__11521 (
            .O(N__52275),
            .I(N__52268));
    InMux I__11520 (
            .O(N__52274),
            .I(N__52265));
    LocalMux I__11519 (
            .O(N__52271),
            .I(N__52262));
    InMux I__11518 (
            .O(N__52268),
            .I(N__52259));
    LocalMux I__11517 (
            .O(N__52265),
            .I(N__52256));
    Span4Mux_v I__11516 (
            .O(N__52262),
            .I(N__52253));
    LocalMux I__11515 (
            .O(N__52259),
            .I(\c0.data_in_frame_7_3 ));
    Odrv4 I__11514 (
            .O(N__52256),
            .I(\c0.data_in_frame_7_3 ));
    Odrv4 I__11513 (
            .O(N__52253),
            .I(\c0.data_in_frame_7_3 ));
    CascadeMux I__11512 (
            .O(N__52246),
            .I(N__52243));
    InMux I__11511 (
            .O(N__52243),
            .I(N__52240));
    LocalMux I__11510 (
            .O(N__52240),
            .I(N__52237));
    Span4Mux_v I__11509 (
            .O(N__52237),
            .I(N__52234));
    Span4Mux_v I__11508 (
            .O(N__52234),
            .I(N__52230));
    InMux I__11507 (
            .O(N__52233),
            .I(N__52226));
    Span4Mux_h I__11506 (
            .O(N__52230),
            .I(N__52223));
    InMux I__11505 (
            .O(N__52229),
            .I(N__52220));
    LocalMux I__11504 (
            .O(N__52226),
            .I(N__52217));
    Odrv4 I__11503 (
            .O(N__52223),
            .I(\c0.n13488 ));
    LocalMux I__11502 (
            .O(N__52220),
            .I(\c0.n13488 ));
    Odrv4 I__11501 (
            .O(N__52217),
            .I(\c0.n13488 ));
    CascadeMux I__11500 (
            .O(N__52210),
            .I(\c0.n22139_cascade_ ));
    CascadeMux I__11499 (
            .O(N__52207),
            .I(N__52203));
    InMux I__11498 (
            .O(N__52206),
            .I(N__52199));
    InMux I__11497 (
            .O(N__52203),
            .I(N__52196));
    InMux I__11496 (
            .O(N__52202),
            .I(N__52193));
    LocalMux I__11495 (
            .O(N__52199),
            .I(N__52190));
    LocalMux I__11494 (
            .O(N__52196),
            .I(\c0.data_in_frame_9_0 ));
    LocalMux I__11493 (
            .O(N__52193),
            .I(\c0.data_in_frame_9_0 ));
    Odrv12 I__11492 (
            .O(N__52190),
            .I(\c0.data_in_frame_9_0 ));
    InMux I__11491 (
            .O(N__52183),
            .I(N__52180));
    LocalMux I__11490 (
            .O(N__52180),
            .I(N__52175));
    InMux I__11489 (
            .O(N__52179),
            .I(N__52172));
    InMux I__11488 (
            .O(N__52178),
            .I(N__52168));
    Span4Mux_v I__11487 (
            .O(N__52175),
            .I(N__52165));
    LocalMux I__11486 (
            .O(N__52172),
            .I(N__52162));
    InMux I__11485 (
            .O(N__52171),
            .I(N__52159));
    LocalMux I__11484 (
            .O(N__52168),
            .I(N__52156));
    Span4Mux_h I__11483 (
            .O(N__52165),
            .I(N__52149));
    Span4Mux_v I__11482 (
            .O(N__52162),
            .I(N__52149));
    LocalMux I__11481 (
            .O(N__52159),
            .I(N__52149));
    Odrv4 I__11480 (
            .O(N__52156),
            .I(\c0.n13605 ));
    Odrv4 I__11479 (
            .O(N__52149),
            .I(\c0.n13605 ));
    InMux I__11478 (
            .O(N__52144),
            .I(N__52138));
    InMux I__11477 (
            .O(N__52143),
            .I(N__52138));
    LocalMux I__11476 (
            .O(N__52138),
            .I(N__52135));
    Span4Mux_h I__11475 (
            .O(N__52135),
            .I(N__52129));
    InMux I__11474 (
            .O(N__52134),
            .I(N__52122));
    InMux I__11473 (
            .O(N__52133),
            .I(N__52122));
    InMux I__11472 (
            .O(N__52132),
            .I(N__52122));
    Span4Mux_v I__11471 (
            .O(N__52129),
            .I(N__52119));
    LocalMux I__11470 (
            .O(N__52122),
            .I(N__52116));
    Odrv4 I__11469 (
            .O(N__52119),
            .I(\c0.n13043 ));
    Odrv12 I__11468 (
            .O(N__52116),
            .I(\c0.n13043 ));
    InMux I__11467 (
            .O(N__52111),
            .I(N__52108));
    LocalMux I__11466 (
            .O(N__52108),
            .I(N__52102));
    InMux I__11465 (
            .O(N__52107),
            .I(N__52099));
    InMux I__11464 (
            .O(N__52106),
            .I(N__52095));
    InMux I__11463 (
            .O(N__52105),
            .I(N__52092));
    Span4Mux_v I__11462 (
            .O(N__52102),
            .I(N__52089));
    LocalMux I__11461 (
            .O(N__52099),
            .I(N__52086));
    InMux I__11460 (
            .O(N__52098),
            .I(N__52083));
    LocalMux I__11459 (
            .O(N__52095),
            .I(\c0.data_in_frame_8_6 ));
    LocalMux I__11458 (
            .O(N__52092),
            .I(\c0.data_in_frame_8_6 ));
    Odrv4 I__11457 (
            .O(N__52089),
            .I(\c0.data_in_frame_8_6 ));
    Odrv12 I__11456 (
            .O(N__52086),
            .I(\c0.data_in_frame_8_6 ));
    LocalMux I__11455 (
            .O(N__52083),
            .I(\c0.data_in_frame_8_6 ));
    CascadeMux I__11454 (
            .O(N__52072),
            .I(\c0.n21822_cascade_ ));
    InMux I__11453 (
            .O(N__52069),
            .I(N__52065));
    CascadeMux I__11452 (
            .O(N__52068),
            .I(N__52062));
    LocalMux I__11451 (
            .O(N__52065),
            .I(N__52059));
    InMux I__11450 (
            .O(N__52062),
            .I(N__52055));
    Span4Mux_h I__11449 (
            .O(N__52059),
            .I(N__52051));
    CascadeMux I__11448 (
            .O(N__52058),
            .I(N__52047));
    LocalMux I__11447 (
            .O(N__52055),
            .I(N__52044));
    InMux I__11446 (
            .O(N__52054),
            .I(N__52041));
    Sp12to4 I__11445 (
            .O(N__52051),
            .I(N__52038));
    InMux I__11444 (
            .O(N__52050),
            .I(N__52035));
    InMux I__11443 (
            .O(N__52047),
            .I(N__52031));
    Span4Mux_v I__11442 (
            .O(N__52044),
            .I(N__52028));
    LocalMux I__11441 (
            .O(N__52041),
            .I(N__52025));
    Span12Mux_v I__11440 (
            .O(N__52038),
            .I(N__52020));
    LocalMux I__11439 (
            .O(N__52035),
            .I(N__52020));
    InMux I__11438 (
            .O(N__52034),
            .I(N__52017));
    LocalMux I__11437 (
            .O(N__52031),
            .I(data_in_frame_1_2));
    Odrv4 I__11436 (
            .O(N__52028),
            .I(data_in_frame_1_2));
    Odrv4 I__11435 (
            .O(N__52025),
            .I(data_in_frame_1_2));
    Odrv12 I__11434 (
            .O(N__52020),
            .I(data_in_frame_1_2));
    LocalMux I__11433 (
            .O(N__52017),
            .I(data_in_frame_1_2));
    InMux I__11432 (
            .O(N__52006),
            .I(N__52003));
    LocalMux I__11431 (
            .O(N__52003),
            .I(\c0.n22334 ));
    CascadeMux I__11430 (
            .O(N__52000),
            .I(\c0.n22334_cascade_ ));
    InMux I__11429 (
            .O(N__51997),
            .I(N__51991));
    InMux I__11428 (
            .O(N__51996),
            .I(N__51991));
    LocalMux I__11427 (
            .O(N__51991),
            .I(N__51987));
    InMux I__11426 (
            .O(N__51990),
            .I(N__51984));
    Odrv4 I__11425 (
            .O(N__51987),
            .I(\c0.n22051 ));
    LocalMux I__11424 (
            .O(N__51984),
            .I(\c0.n22051 ));
    InMux I__11423 (
            .O(N__51979),
            .I(N__51975));
    InMux I__11422 (
            .O(N__51978),
            .I(N__51971));
    LocalMux I__11421 (
            .O(N__51975),
            .I(N__51967));
    InMux I__11420 (
            .O(N__51974),
            .I(N__51964));
    LocalMux I__11419 (
            .O(N__51971),
            .I(N__51961));
    InMux I__11418 (
            .O(N__51970),
            .I(N__51958));
    Span4Mux_h I__11417 (
            .O(N__51967),
            .I(N__51953));
    LocalMux I__11416 (
            .O(N__51964),
            .I(N__51953));
    Span4Mux_h I__11415 (
            .O(N__51961),
            .I(N__51950));
    LocalMux I__11414 (
            .O(N__51958),
            .I(\c0.n15_adj_4404 ));
    Odrv4 I__11413 (
            .O(N__51953),
            .I(\c0.n15_adj_4404 ));
    Odrv4 I__11412 (
            .O(N__51950),
            .I(\c0.n15_adj_4404 ));
    InMux I__11411 (
            .O(N__51943),
            .I(N__51939));
    CascadeMux I__11410 (
            .O(N__51942),
            .I(N__51935));
    LocalMux I__11409 (
            .O(N__51939),
            .I(N__51932));
    InMux I__11408 (
            .O(N__51938),
            .I(N__51927));
    InMux I__11407 (
            .O(N__51935),
            .I(N__51927));
    Span4Mux_v I__11406 (
            .O(N__51932),
            .I(N__51924));
    LocalMux I__11405 (
            .O(N__51927),
            .I(\c0.data_in_frame_8_0 ));
    Odrv4 I__11404 (
            .O(N__51924),
            .I(\c0.data_in_frame_8_0 ));
    CascadeMux I__11403 (
            .O(N__51919),
            .I(N__51915));
    CascadeMux I__11402 (
            .O(N__51918),
            .I(N__51911));
    InMux I__11401 (
            .O(N__51915),
            .I(N__51907));
    InMux I__11400 (
            .O(N__51914),
            .I(N__51904));
    InMux I__11399 (
            .O(N__51911),
            .I(N__51899));
    InMux I__11398 (
            .O(N__51910),
            .I(N__51899));
    LocalMux I__11397 (
            .O(N__51907),
            .I(\c0.data_in_frame_7_7 ));
    LocalMux I__11396 (
            .O(N__51904),
            .I(\c0.data_in_frame_7_7 ));
    LocalMux I__11395 (
            .O(N__51899),
            .I(\c0.data_in_frame_7_7 ));
    InMux I__11394 (
            .O(N__51892),
            .I(N__51889));
    LocalMux I__11393 (
            .O(N__51889),
            .I(\c0.n6_adj_4259 ));
    InMux I__11392 (
            .O(N__51886),
            .I(N__51883));
    LocalMux I__11391 (
            .O(N__51883),
            .I(N__51880));
    Odrv4 I__11390 (
            .O(N__51880),
            .I(\c0.n39_adj_4263 ));
    InMux I__11389 (
            .O(N__51877),
            .I(N__51874));
    LocalMux I__11388 (
            .O(N__51874),
            .I(N__51871));
    Odrv4 I__11387 (
            .O(N__51871),
            .I(\c0.n40_adj_4261 ));
    CascadeMux I__11386 (
            .O(N__51868),
            .I(\c0.n22060_cascade_ ));
    InMux I__11385 (
            .O(N__51865),
            .I(N__51862));
    LocalMux I__11384 (
            .O(N__51862),
            .I(\c0.n44_adj_4262 ));
    CascadeMux I__11383 (
            .O(N__51859),
            .I(\c0.n11_adj_4266_cascade_ ));
    InMux I__11382 (
            .O(N__51856),
            .I(N__51851));
    InMux I__11381 (
            .O(N__51855),
            .I(N__51846));
    InMux I__11380 (
            .O(N__51854),
            .I(N__51846));
    LocalMux I__11379 (
            .O(N__51851),
            .I(\c0.n13425 ));
    LocalMux I__11378 (
            .O(N__51846),
            .I(\c0.n13425 ));
    CascadeMux I__11377 (
            .O(N__51841),
            .I(\c0.n22842_cascade_ ));
    InMux I__11376 (
            .O(N__51838),
            .I(N__51833));
    InMux I__11375 (
            .O(N__51837),
            .I(N__51830));
    InMux I__11374 (
            .O(N__51836),
            .I(N__51827));
    LocalMux I__11373 (
            .O(N__51833),
            .I(\c0.data_in_frame_5_6 ));
    LocalMux I__11372 (
            .O(N__51830),
            .I(\c0.data_in_frame_5_6 ));
    LocalMux I__11371 (
            .O(N__51827),
            .I(\c0.data_in_frame_5_6 ));
    InMux I__11370 (
            .O(N__51820),
            .I(N__51816));
    InMux I__11369 (
            .O(N__51819),
            .I(N__51813));
    LocalMux I__11368 (
            .O(N__51816),
            .I(N__51810));
    LocalMux I__11367 (
            .O(N__51813),
            .I(\c0.n22283 ));
    Odrv12 I__11366 (
            .O(N__51810),
            .I(\c0.n22283 ));
    CascadeMux I__11365 (
            .O(N__51805),
            .I(\c0.n13488_cascade_ ));
    InMux I__11364 (
            .O(N__51802),
            .I(N__51797));
    InMux I__11363 (
            .O(N__51801),
            .I(N__51794));
    InMux I__11362 (
            .O(N__51800),
            .I(N__51791));
    LocalMux I__11361 (
            .O(N__51797),
            .I(N__51788));
    LocalMux I__11360 (
            .O(N__51794),
            .I(N__51785));
    LocalMux I__11359 (
            .O(N__51791),
            .I(\c0.n13180 ));
    Odrv12 I__11358 (
            .O(N__51788),
            .I(\c0.n13180 ));
    Odrv12 I__11357 (
            .O(N__51785),
            .I(\c0.n13180 ));
    InMux I__11356 (
            .O(N__51778),
            .I(N__51768));
    InMux I__11355 (
            .O(N__51777),
            .I(N__51768));
    InMux I__11354 (
            .O(N__51776),
            .I(N__51765));
    InMux I__11353 (
            .O(N__51775),
            .I(N__51762));
    InMux I__11352 (
            .O(N__51774),
            .I(N__51759));
    CascadeMux I__11351 (
            .O(N__51773),
            .I(N__51756));
    LocalMux I__11350 (
            .O(N__51768),
            .I(N__51750));
    LocalMux I__11349 (
            .O(N__51765),
            .I(N__51747));
    LocalMux I__11348 (
            .O(N__51762),
            .I(N__51744));
    LocalMux I__11347 (
            .O(N__51759),
            .I(N__51741));
    InMux I__11346 (
            .O(N__51756),
            .I(N__51738));
    InMux I__11345 (
            .O(N__51755),
            .I(N__51733));
    InMux I__11344 (
            .O(N__51754),
            .I(N__51733));
    InMux I__11343 (
            .O(N__51753),
            .I(N__51730));
    Span4Mux_h I__11342 (
            .O(N__51750),
            .I(N__51721));
    Span4Mux_v I__11341 (
            .O(N__51747),
            .I(N__51721));
    Span4Mux_h I__11340 (
            .O(N__51744),
            .I(N__51721));
    Span4Mux_v I__11339 (
            .O(N__51741),
            .I(N__51721));
    LocalMux I__11338 (
            .O(N__51738),
            .I(\c0.data_in_frame_0_5 ));
    LocalMux I__11337 (
            .O(N__51733),
            .I(\c0.data_in_frame_0_5 ));
    LocalMux I__11336 (
            .O(N__51730),
            .I(\c0.data_in_frame_0_5 ));
    Odrv4 I__11335 (
            .O(N__51721),
            .I(\c0.data_in_frame_0_5 ));
    InMux I__11334 (
            .O(N__51712),
            .I(N__51707));
    InMux I__11333 (
            .O(N__51711),
            .I(N__51704));
    InMux I__11332 (
            .O(N__51710),
            .I(N__51701));
    LocalMux I__11331 (
            .O(N__51707),
            .I(N__51697));
    LocalMux I__11330 (
            .O(N__51704),
            .I(N__51694));
    LocalMux I__11329 (
            .O(N__51701),
            .I(N__51691));
    InMux I__11328 (
            .O(N__51700),
            .I(N__51688));
    Span4Mux_h I__11327 (
            .O(N__51697),
            .I(N__51680));
    Span4Mux_v I__11326 (
            .O(N__51694),
            .I(N__51673));
    Span4Mux_h I__11325 (
            .O(N__51691),
            .I(N__51673));
    LocalMux I__11324 (
            .O(N__51688),
            .I(N__51673));
    InMux I__11323 (
            .O(N__51687),
            .I(N__51670));
    InMux I__11322 (
            .O(N__51686),
            .I(N__51665));
    InMux I__11321 (
            .O(N__51685),
            .I(N__51665));
    InMux I__11320 (
            .O(N__51684),
            .I(N__51660));
    InMux I__11319 (
            .O(N__51683),
            .I(N__51660));
    Odrv4 I__11318 (
            .O(N__51680),
            .I(\c0.data_in_frame_0_6 ));
    Odrv4 I__11317 (
            .O(N__51673),
            .I(\c0.data_in_frame_0_6 ));
    LocalMux I__11316 (
            .O(N__51670),
            .I(\c0.data_in_frame_0_6 ));
    LocalMux I__11315 (
            .O(N__51665),
            .I(\c0.data_in_frame_0_6 ));
    LocalMux I__11314 (
            .O(N__51660),
            .I(\c0.data_in_frame_0_6 ));
    CascadeMux I__11313 (
            .O(N__51649),
            .I(N__51646));
    InMux I__11312 (
            .O(N__51646),
            .I(N__51643));
    LocalMux I__11311 (
            .O(N__51643),
            .I(N__51640));
    Span4Mux_h I__11310 (
            .O(N__51640),
            .I(N__51637));
    Span4Mux_v I__11309 (
            .O(N__51637),
            .I(N__51634));
    Odrv4 I__11308 (
            .O(N__51634),
            .I(\c0.n23827 ));
    InMux I__11307 (
            .O(N__51631),
            .I(N__51627));
    CascadeMux I__11306 (
            .O(N__51630),
            .I(N__51624));
    LocalMux I__11305 (
            .O(N__51627),
            .I(N__51619));
    InMux I__11304 (
            .O(N__51624),
            .I(N__51616));
    InMux I__11303 (
            .O(N__51623),
            .I(N__51613));
    InMux I__11302 (
            .O(N__51622),
            .I(N__51610));
    Sp12to4 I__11301 (
            .O(N__51619),
            .I(N__51607));
    LocalMux I__11300 (
            .O(N__51616),
            .I(\c0.data_in_frame_5_3 ));
    LocalMux I__11299 (
            .O(N__51613),
            .I(\c0.data_in_frame_5_3 ));
    LocalMux I__11298 (
            .O(N__51610),
            .I(\c0.data_in_frame_5_3 ));
    Odrv12 I__11297 (
            .O(N__51607),
            .I(\c0.data_in_frame_5_3 ));
    CascadeMux I__11296 (
            .O(N__51598),
            .I(N__51593));
    CascadeMux I__11295 (
            .O(N__51597),
            .I(N__51589));
    InMux I__11294 (
            .O(N__51596),
            .I(N__51586));
    InMux I__11293 (
            .O(N__51593),
            .I(N__51581));
    InMux I__11292 (
            .O(N__51592),
            .I(N__51581));
    InMux I__11291 (
            .O(N__51589),
            .I(N__51578));
    LocalMux I__11290 (
            .O(N__51586),
            .I(\c0.data_in_frame_7_5 ));
    LocalMux I__11289 (
            .O(N__51581),
            .I(\c0.data_in_frame_7_5 ));
    LocalMux I__11288 (
            .O(N__51578),
            .I(\c0.data_in_frame_7_5 ));
    InMux I__11287 (
            .O(N__51571),
            .I(N__51568));
    LocalMux I__11286 (
            .O(N__51568),
            .I(N__51563));
    InMux I__11285 (
            .O(N__51567),
            .I(N__51560));
    InMux I__11284 (
            .O(N__51566),
            .I(N__51557));
    Odrv4 I__11283 (
            .O(N__51563),
            .I(\c0.n12484 ));
    LocalMux I__11282 (
            .O(N__51560),
            .I(\c0.n12484 ));
    LocalMux I__11281 (
            .O(N__51557),
            .I(\c0.n12484 ));
    CascadeMux I__11280 (
            .O(N__51550),
            .I(\c0.n20368_cascade_ ));
    CascadeMux I__11279 (
            .O(N__51547),
            .I(N__51544));
    InMux I__11278 (
            .O(N__51544),
            .I(N__51540));
    InMux I__11277 (
            .O(N__51543),
            .I(N__51537));
    LocalMux I__11276 (
            .O(N__51540),
            .I(N__51534));
    LocalMux I__11275 (
            .O(N__51537),
            .I(N__51531));
    Odrv4 I__11274 (
            .O(N__51534),
            .I(\c0.data_in_frame_10_1 ));
    Odrv4 I__11273 (
            .O(N__51531),
            .I(\c0.data_in_frame_10_1 ));
    CascadeMux I__11272 (
            .O(N__51526),
            .I(\c0.n22133_cascade_ ));
    InMux I__11271 (
            .O(N__51523),
            .I(N__51520));
    LocalMux I__11270 (
            .O(N__51520),
            .I(\c0.n21925 ));
    CascadeMux I__11269 (
            .O(N__51517),
            .I(\c0.n20927_cascade_ ));
    InMux I__11268 (
            .O(N__51514),
            .I(N__51511));
    LocalMux I__11267 (
            .O(N__51511),
            .I(\c0.n22133 ));
    InMux I__11266 (
            .O(N__51508),
            .I(N__51505));
    LocalMux I__11265 (
            .O(N__51505),
            .I(\c0.n36 ));
    InMux I__11264 (
            .O(N__51502),
            .I(\c0.rx.n19539 ));
    CEMux I__11263 (
            .O(N__51499),
            .I(N__51496));
    LocalMux I__11262 (
            .O(N__51496),
            .I(N__51493));
    Span4Mux_h I__11261 (
            .O(N__51493),
            .I(N__51490));
    Span4Mux_h I__11260 (
            .O(N__51490),
            .I(N__51487));
    Odrv4 I__11259 (
            .O(N__51487),
            .I(\c0.rx.n14391 ));
    SRMux I__11258 (
            .O(N__51484),
            .I(N__51481));
    LocalMux I__11257 (
            .O(N__51481),
            .I(N__51478));
    Odrv12 I__11256 (
            .O(N__51478),
            .I(\c0.rx.n17411 ));
    InMux I__11255 (
            .O(N__51475),
            .I(N__51467));
    InMux I__11254 (
            .O(N__51474),
            .I(N__51458));
    InMux I__11253 (
            .O(N__51473),
            .I(N__51458));
    InMux I__11252 (
            .O(N__51472),
            .I(N__51455));
    InMux I__11251 (
            .O(N__51471),
            .I(N__51452));
    InMux I__11250 (
            .O(N__51470),
            .I(N__51445));
    LocalMux I__11249 (
            .O(N__51467),
            .I(N__51440));
    InMux I__11248 (
            .O(N__51466),
            .I(N__51437));
    InMux I__11247 (
            .O(N__51465),
            .I(N__51426));
    InMux I__11246 (
            .O(N__51464),
            .I(N__51426));
    InMux I__11245 (
            .O(N__51463),
            .I(N__51426));
    LocalMux I__11244 (
            .O(N__51458),
            .I(N__51423));
    LocalMux I__11243 (
            .O(N__51455),
            .I(N__51420));
    LocalMux I__11242 (
            .O(N__51452),
            .I(N__51417));
    InMux I__11241 (
            .O(N__51451),
            .I(N__51414));
    InMux I__11240 (
            .O(N__51450),
            .I(N__51404));
    InMux I__11239 (
            .O(N__51449),
            .I(N__51404));
    InMux I__11238 (
            .O(N__51448),
            .I(N__51399));
    LocalMux I__11237 (
            .O(N__51445),
            .I(N__51395));
    InMux I__11236 (
            .O(N__51444),
            .I(N__51390));
    InMux I__11235 (
            .O(N__51443),
            .I(N__51390));
    Span4Mux_h I__11234 (
            .O(N__51440),
            .I(N__51383));
    LocalMux I__11233 (
            .O(N__51437),
            .I(N__51383));
    InMux I__11232 (
            .O(N__51436),
            .I(N__51380));
    InMux I__11231 (
            .O(N__51435),
            .I(N__51373));
    InMux I__11230 (
            .O(N__51434),
            .I(N__51373));
    InMux I__11229 (
            .O(N__51433),
            .I(N__51373));
    LocalMux I__11228 (
            .O(N__51426),
            .I(N__51368));
    Span4Mux_v I__11227 (
            .O(N__51423),
            .I(N__51363));
    Span4Mux_h I__11226 (
            .O(N__51420),
            .I(N__51356));
    Span4Mux_v I__11225 (
            .O(N__51417),
            .I(N__51356));
    LocalMux I__11224 (
            .O(N__51414),
            .I(N__51356));
    InMux I__11223 (
            .O(N__51413),
            .I(N__51351));
    InMux I__11222 (
            .O(N__51412),
            .I(N__51351));
    InMux I__11221 (
            .O(N__51411),
            .I(N__51348));
    InMux I__11220 (
            .O(N__51410),
            .I(N__51343));
    InMux I__11219 (
            .O(N__51409),
            .I(N__51343));
    LocalMux I__11218 (
            .O(N__51404),
            .I(N__51340));
    InMux I__11217 (
            .O(N__51403),
            .I(N__51335));
    InMux I__11216 (
            .O(N__51402),
            .I(N__51335));
    LocalMux I__11215 (
            .O(N__51399),
            .I(N__51332));
    InMux I__11214 (
            .O(N__51398),
            .I(N__51329));
    Span4Mux_h I__11213 (
            .O(N__51395),
            .I(N__51326));
    LocalMux I__11212 (
            .O(N__51390),
            .I(N__51323));
    InMux I__11211 (
            .O(N__51389),
            .I(N__51317));
    InMux I__11210 (
            .O(N__51388),
            .I(N__51317));
    Span4Mux_v I__11209 (
            .O(N__51383),
            .I(N__51312));
    LocalMux I__11208 (
            .O(N__51380),
            .I(N__51312));
    LocalMux I__11207 (
            .O(N__51373),
            .I(N__51309));
    InMux I__11206 (
            .O(N__51372),
            .I(N__51304));
    InMux I__11205 (
            .O(N__51371),
            .I(N__51304));
    Span4Mux_h I__11204 (
            .O(N__51368),
            .I(N__51301));
    InMux I__11203 (
            .O(N__51367),
            .I(N__51296));
    InMux I__11202 (
            .O(N__51366),
            .I(N__51296));
    Sp12to4 I__11201 (
            .O(N__51363),
            .I(N__51293));
    Span4Mux_h I__11200 (
            .O(N__51356),
            .I(N__51290));
    LocalMux I__11199 (
            .O(N__51351),
            .I(N__51287));
    LocalMux I__11198 (
            .O(N__51348),
            .I(N__51282));
    LocalMux I__11197 (
            .O(N__51343),
            .I(N__51282));
    Span4Mux_v I__11196 (
            .O(N__51340),
            .I(N__51277));
    LocalMux I__11195 (
            .O(N__51335),
            .I(N__51277));
    Span4Mux_v I__11194 (
            .O(N__51332),
            .I(N__51272));
    LocalMux I__11193 (
            .O(N__51329),
            .I(N__51272));
    Span4Mux_h I__11192 (
            .O(N__51326),
            .I(N__51267));
    Span4Mux_h I__11191 (
            .O(N__51323),
            .I(N__51267));
    InMux I__11190 (
            .O(N__51322),
            .I(N__51264));
    LocalMux I__11189 (
            .O(N__51317),
            .I(N__51257));
    Span4Mux_v I__11188 (
            .O(N__51312),
            .I(N__51257));
    Span4Mux_v I__11187 (
            .O(N__51309),
            .I(N__51257));
    LocalMux I__11186 (
            .O(N__51304),
            .I(N__51250));
    Span4Mux_h I__11185 (
            .O(N__51301),
            .I(N__51250));
    LocalMux I__11184 (
            .O(N__51296),
            .I(N__51250));
    Span12Mux_h I__11183 (
            .O(N__51293),
            .I(N__51247));
    Sp12to4 I__11182 (
            .O(N__51290),
            .I(N__51244));
    Span4Mux_v I__11181 (
            .O(N__51287),
            .I(N__51239));
    Span4Mux_v I__11180 (
            .O(N__51282),
            .I(N__51239));
    Span4Mux_h I__11179 (
            .O(N__51277),
            .I(N__51236));
    Span4Mux_h I__11178 (
            .O(N__51272),
            .I(N__51231));
    Span4Mux_v I__11177 (
            .O(N__51267),
            .I(N__51231));
    LocalMux I__11176 (
            .O(N__51264),
            .I(N__51224));
    Span4Mux_h I__11175 (
            .O(N__51257),
            .I(N__51224));
    Span4Mux_v I__11174 (
            .O(N__51250),
            .I(N__51224));
    Span12Mux_v I__11173 (
            .O(N__51247),
            .I(N__51221));
    Span12Mux_s10_v I__11172 (
            .O(N__51244),
            .I(N__51218));
    Odrv4 I__11171 (
            .O(N__51239),
            .I(\c0.data_out_frame_29_7_N_1483_0 ));
    Odrv4 I__11170 (
            .O(N__51236),
            .I(\c0.data_out_frame_29_7_N_1483_0 ));
    Odrv4 I__11169 (
            .O(N__51231),
            .I(\c0.data_out_frame_29_7_N_1483_0 ));
    Odrv4 I__11168 (
            .O(N__51224),
            .I(\c0.data_out_frame_29_7_N_1483_0 ));
    Odrv12 I__11167 (
            .O(N__51221),
            .I(\c0.data_out_frame_29_7_N_1483_0 ));
    Odrv12 I__11166 (
            .O(N__51218),
            .I(\c0.data_out_frame_29_7_N_1483_0 ));
    InMux I__11165 (
            .O(N__51205),
            .I(N__51200));
    InMux I__11164 (
            .O(N__51204),
            .I(N__51197));
    InMux I__11163 (
            .O(N__51203),
            .I(N__51194));
    LocalMux I__11162 (
            .O(N__51200),
            .I(N__51182));
    LocalMux I__11161 (
            .O(N__51197),
            .I(N__51182));
    LocalMux I__11160 (
            .O(N__51194),
            .I(N__51182));
    InMux I__11159 (
            .O(N__51193),
            .I(N__51179));
    InMux I__11158 (
            .O(N__51192),
            .I(N__51176));
    InMux I__11157 (
            .O(N__51191),
            .I(N__51169));
    InMux I__11156 (
            .O(N__51190),
            .I(N__51166));
    InMux I__11155 (
            .O(N__51189),
            .I(N__51163));
    Span4Mux_v I__11154 (
            .O(N__51182),
            .I(N__51151));
    LocalMux I__11153 (
            .O(N__51179),
            .I(N__51151));
    LocalMux I__11152 (
            .O(N__51176),
            .I(N__51151));
    InMux I__11151 (
            .O(N__51175),
            .I(N__51148));
    InMux I__11150 (
            .O(N__51174),
            .I(N__51145));
    InMux I__11149 (
            .O(N__51173),
            .I(N__51142));
    InMux I__11148 (
            .O(N__51172),
            .I(N__51139));
    LocalMux I__11147 (
            .O(N__51169),
            .I(N__51132));
    LocalMux I__11146 (
            .O(N__51166),
            .I(N__51132));
    LocalMux I__11145 (
            .O(N__51163),
            .I(N__51132));
    InMux I__11144 (
            .O(N__51162),
            .I(N__51127));
    InMux I__11143 (
            .O(N__51161),
            .I(N__51124));
    InMux I__11142 (
            .O(N__51160),
            .I(N__51119));
    InMux I__11141 (
            .O(N__51159),
            .I(N__51114));
    InMux I__11140 (
            .O(N__51158),
            .I(N__51114));
    Span4Mux_v I__11139 (
            .O(N__51151),
            .I(N__51104));
    LocalMux I__11138 (
            .O(N__51148),
            .I(N__51104));
    LocalMux I__11137 (
            .O(N__51145),
            .I(N__51104));
    LocalMux I__11136 (
            .O(N__51142),
            .I(N__51101));
    LocalMux I__11135 (
            .O(N__51139),
            .I(N__51093));
    Span4Mux_h I__11134 (
            .O(N__51132),
            .I(N__51090));
    InMux I__11133 (
            .O(N__51131),
            .I(N__51082));
    InMux I__11132 (
            .O(N__51130),
            .I(N__51079));
    LocalMux I__11131 (
            .O(N__51127),
            .I(N__51074));
    LocalMux I__11130 (
            .O(N__51124),
            .I(N__51074));
    InMux I__11129 (
            .O(N__51123),
            .I(N__51071));
    InMux I__11128 (
            .O(N__51122),
            .I(N__51061));
    LocalMux I__11127 (
            .O(N__51119),
            .I(N__51056));
    LocalMux I__11126 (
            .O(N__51114),
            .I(N__51056));
    InMux I__11125 (
            .O(N__51113),
            .I(N__51049));
    InMux I__11124 (
            .O(N__51112),
            .I(N__51046));
    CascadeMux I__11123 (
            .O(N__51111),
            .I(N__51043));
    Span4Mux_v I__11122 (
            .O(N__51104),
            .I(N__51036));
    Span4Mux_s1_v I__11121 (
            .O(N__51101),
            .I(N__51036));
    InMux I__11120 (
            .O(N__51100),
            .I(N__51033));
    InMux I__11119 (
            .O(N__51099),
            .I(N__51030));
    InMux I__11118 (
            .O(N__51098),
            .I(N__51027));
    InMux I__11117 (
            .O(N__51097),
            .I(N__51024));
    InMux I__11116 (
            .O(N__51096),
            .I(N__51021));
    Span4Mux_h I__11115 (
            .O(N__51093),
            .I(N__51016));
    Span4Mux_v I__11114 (
            .O(N__51090),
            .I(N__51016));
    CascadeMux I__11113 (
            .O(N__51089),
            .I(N__51013));
    InMux I__11112 (
            .O(N__51088),
            .I(N__51007));
    InMux I__11111 (
            .O(N__51087),
            .I(N__51004));
    InMux I__11110 (
            .O(N__51086),
            .I(N__51001));
    InMux I__11109 (
            .O(N__51085),
            .I(N__50998));
    LocalMux I__11108 (
            .O(N__51082),
            .I(N__50995));
    LocalMux I__11107 (
            .O(N__51079),
            .I(N__50988));
    Span4Mux_s2_v I__11106 (
            .O(N__51074),
            .I(N__50988));
    LocalMux I__11105 (
            .O(N__51071),
            .I(N__50988));
    CascadeMux I__11104 (
            .O(N__51070),
            .I(N__50984));
    InMux I__11103 (
            .O(N__51069),
            .I(N__50981));
    InMux I__11102 (
            .O(N__51068),
            .I(N__50975));
    InMux I__11101 (
            .O(N__51067),
            .I(N__50975));
    CascadeMux I__11100 (
            .O(N__51066),
            .I(N__50970));
    CascadeMux I__11099 (
            .O(N__51065),
            .I(N__50966));
    InMux I__11098 (
            .O(N__51064),
            .I(N__50963));
    LocalMux I__11097 (
            .O(N__51061),
            .I(N__50956));
    Span4Mux_h I__11096 (
            .O(N__51056),
            .I(N__50956));
    InMux I__11095 (
            .O(N__51055),
            .I(N__50951));
    InMux I__11094 (
            .O(N__51054),
            .I(N__50948));
    InMux I__11093 (
            .O(N__51053),
            .I(N__50945));
    InMux I__11092 (
            .O(N__51052),
            .I(N__50942));
    LocalMux I__11091 (
            .O(N__51049),
            .I(N__50937));
    LocalMux I__11090 (
            .O(N__51046),
            .I(N__50937));
    InMux I__11089 (
            .O(N__51043),
            .I(N__50930));
    InMux I__11088 (
            .O(N__51042),
            .I(N__50930));
    InMux I__11087 (
            .O(N__51041),
            .I(N__50930));
    Sp12to4 I__11086 (
            .O(N__51036),
            .I(N__50924));
    LocalMux I__11085 (
            .O(N__51033),
            .I(N__50924));
    LocalMux I__11084 (
            .O(N__51030),
            .I(N__50919));
    LocalMux I__11083 (
            .O(N__51027),
            .I(N__50919));
    LocalMux I__11082 (
            .O(N__51024),
            .I(N__50914));
    LocalMux I__11081 (
            .O(N__51021),
            .I(N__50914));
    Span4Mux_v I__11080 (
            .O(N__51016),
            .I(N__50911));
    InMux I__11079 (
            .O(N__51013),
            .I(N__50904));
    InMux I__11078 (
            .O(N__51012),
            .I(N__50904));
    InMux I__11077 (
            .O(N__51011),
            .I(N__50904));
    InMux I__11076 (
            .O(N__51010),
            .I(N__50901));
    LocalMux I__11075 (
            .O(N__51007),
            .I(N__50888));
    LocalMux I__11074 (
            .O(N__51004),
            .I(N__50888));
    LocalMux I__11073 (
            .O(N__51001),
            .I(N__50888));
    LocalMux I__11072 (
            .O(N__50998),
            .I(N__50888));
    Span4Mux_v I__11071 (
            .O(N__50995),
            .I(N__50888));
    Span4Mux_v I__11070 (
            .O(N__50988),
            .I(N__50888));
    InMux I__11069 (
            .O(N__50987),
            .I(N__50883));
    InMux I__11068 (
            .O(N__50984),
            .I(N__50883));
    LocalMux I__11067 (
            .O(N__50981),
            .I(N__50880));
    InMux I__11066 (
            .O(N__50980),
            .I(N__50877));
    LocalMux I__11065 (
            .O(N__50975),
            .I(N__50874));
    InMux I__11064 (
            .O(N__50974),
            .I(N__50871));
    InMux I__11063 (
            .O(N__50973),
            .I(N__50866));
    InMux I__11062 (
            .O(N__50970),
            .I(N__50866));
    InMux I__11061 (
            .O(N__50969),
            .I(N__50861));
    InMux I__11060 (
            .O(N__50966),
            .I(N__50861));
    LocalMux I__11059 (
            .O(N__50963),
            .I(N__50858));
    InMux I__11058 (
            .O(N__50962),
            .I(N__50853));
    InMux I__11057 (
            .O(N__50961),
            .I(N__50853));
    Sp12to4 I__11056 (
            .O(N__50956),
            .I(N__50850));
    InMux I__11055 (
            .O(N__50955),
            .I(N__50846));
    InMux I__11054 (
            .O(N__50954),
            .I(N__50843));
    LocalMux I__11053 (
            .O(N__50951),
            .I(N__50830));
    LocalMux I__11052 (
            .O(N__50948),
            .I(N__50830));
    LocalMux I__11051 (
            .O(N__50945),
            .I(N__50830));
    LocalMux I__11050 (
            .O(N__50942),
            .I(N__50830));
    Span4Mux_v I__11049 (
            .O(N__50937),
            .I(N__50830));
    LocalMux I__11048 (
            .O(N__50930),
            .I(N__50830));
    InMux I__11047 (
            .O(N__50929),
            .I(N__50827));
    Span12Mux_h I__11046 (
            .O(N__50924),
            .I(N__50823));
    Span4Mux_h I__11045 (
            .O(N__50919),
            .I(N__50820));
    Span4Mux_h I__11044 (
            .O(N__50914),
            .I(N__50813));
    Span4Mux_v I__11043 (
            .O(N__50911),
            .I(N__50813));
    LocalMux I__11042 (
            .O(N__50904),
            .I(N__50813));
    LocalMux I__11041 (
            .O(N__50901),
            .I(N__50810));
    Span4Mux_v I__11040 (
            .O(N__50888),
            .I(N__50803));
    LocalMux I__11039 (
            .O(N__50883),
            .I(N__50803));
    Span4Mux_h I__11038 (
            .O(N__50880),
            .I(N__50803));
    LocalMux I__11037 (
            .O(N__50877),
            .I(N__50791));
    Sp12to4 I__11036 (
            .O(N__50874),
            .I(N__50791));
    LocalMux I__11035 (
            .O(N__50871),
            .I(N__50791));
    LocalMux I__11034 (
            .O(N__50866),
            .I(N__50791));
    LocalMux I__11033 (
            .O(N__50861),
            .I(N__50791));
    Span12Mux_h I__11032 (
            .O(N__50858),
            .I(N__50784));
    LocalMux I__11031 (
            .O(N__50853),
            .I(N__50784));
    Span12Mux_s7_v I__11030 (
            .O(N__50850),
            .I(N__50784));
    CascadeMux I__11029 (
            .O(N__50849),
            .I(N__50781));
    LocalMux I__11028 (
            .O(N__50846),
            .I(N__50768));
    LocalMux I__11027 (
            .O(N__50843),
            .I(N__50768));
    Span4Mux_v I__11026 (
            .O(N__50830),
            .I(N__50768));
    LocalMux I__11025 (
            .O(N__50827),
            .I(N__50768));
    InMux I__11024 (
            .O(N__50826),
            .I(N__50765));
    Span12Mux_v I__11023 (
            .O(N__50823),
            .I(N__50762));
    Span4Mux_v I__11022 (
            .O(N__50820),
            .I(N__50757));
    Span4Mux_v I__11021 (
            .O(N__50813),
            .I(N__50757));
    Span4Mux_h I__11020 (
            .O(N__50810),
            .I(N__50752));
    Span4Mux_h I__11019 (
            .O(N__50803),
            .I(N__50752));
    InMux I__11018 (
            .O(N__50802),
            .I(N__50749));
    Span12Mux_v I__11017 (
            .O(N__50791),
            .I(N__50744));
    Span12Mux_v I__11016 (
            .O(N__50784),
            .I(N__50744));
    InMux I__11015 (
            .O(N__50781),
            .I(N__50739));
    InMux I__11014 (
            .O(N__50780),
            .I(N__50739));
    InMux I__11013 (
            .O(N__50779),
            .I(N__50732));
    InMux I__11012 (
            .O(N__50778),
            .I(N__50732));
    InMux I__11011 (
            .O(N__50777),
            .I(N__50732));
    Span4Mux_h I__11010 (
            .O(N__50768),
            .I(N__50729));
    LocalMux I__11009 (
            .O(N__50765),
            .I(\c0.n1220 ));
    Odrv12 I__11008 (
            .O(N__50762),
            .I(\c0.n1220 ));
    Odrv4 I__11007 (
            .O(N__50757),
            .I(\c0.n1220 ));
    Odrv4 I__11006 (
            .O(N__50752),
            .I(\c0.n1220 ));
    LocalMux I__11005 (
            .O(N__50749),
            .I(\c0.n1220 ));
    Odrv12 I__11004 (
            .O(N__50744),
            .I(\c0.n1220 ));
    LocalMux I__11003 (
            .O(N__50739),
            .I(\c0.n1220 ));
    LocalMux I__11002 (
            .O(N__50732),
            .I(\c0.n1220 ));
    Odrv4 I__11001 (
            .O(N__50729),
            .I(\c0.n1220 ));
    InMux I__11000 (
            .O(N__50710),
            .I(N__50706));
    CascadeMux I__10999 (
            .O(N__50709),
            .I(N__50703));
    LocalMux I__10998 (
            .O(N__50706),
            .I(N__50700));
    InMux I__10997 (
            .O(N__50703),
            .I(N__50696));
    Span4Mux_v I__10996 (
            .O(N__50700),
            .I(N__50693));
    InMux I__10995 (
            .O(N__50699),
            .I(N__50690));
    LocalMux I__10994 (
            .O(N__50696),
            .I(N__50685));
    Span4Mux_v I__10993 (
            .O(N__50693),
            .I(N__50685));
    LocalMux I__10992 (
            .O(N__50690),
            .I(\c0.FRAME_MATCHER_i_28 ));
    Odrv4 I__10991 (
            .O(N__50685),
            .I(\c0.FRAME_MATCHER_i_28 ));
    InMux I__10990 (
            .O(N__50680),
            .I(N__50675));
    CascadeMux I__10989 (
            .O(N__50679),
            .I(N__50670));
    InMux I__10988 (
            .O(N__50678),
            .I(N__50655));
    LocalMux I__10987 (
            .O(N__50675),
            .I(N__50652));
    InMux I__10986 (
            .O(N__50674),
            .I(N__50643));
    InMux I__10985 (
            .O(N__50673),
            .I(N__50640));
    InMux I__10984 (
            .O(N__50670),
            .I(N__50637));
    InMux I__10983 (
            .O(N__50669),
            .I(N__50632));
    InMux I__10982 (
            .O(N__50668),
            .I(N__50632));
    InMux I__10981 (
            .O(N__50667),
            .I(N__50629));
    InMux I__10980 (
            .O(N__50666),
            .I(N__50622));
    InMux I__10979 (
            .O(N__50665),
            .I(N__50622));
    InMux I__10978 (
            .O(N__50664),
            .I(N__50622));
    InMux I__10977 (
            .O(N__50663),
            .I(N__50617));
    InMux I__10976 (
            .O(N__50662),
            .I(N__50612));
    InMux I__10975 (
            .O(N__50661),
            .I(N__50612));
    InMux I__10974 (
            .O(N__50660),
            .I(N__50606));
    InMux I__10973 (
            .O(N__50659),
            .I(N__50601));
    InMux I__10972 (
            .O(N__50658),
            .I(N__50601));
    LocalMux I__10971 (
            .O(N__50655),
            .I(N__50596));
    Span4Mux_v I__10970 (
            .O(N__50652),
            .I(N__50596));
    InMux I__10969 (
            .O(N__50651),
            .I(N__50591));
    InMux I__10968 (
            .O(N__50650),
            .I(N__50588));
    InMux I__10967 (
            .O(N__50649),
            .I(N__50583));
    InMux I__10966 (
            .O(N__50648),
            .I(N__50583));
    InMux I__10965 (
            .O(N__50647),
            .I(N__50578));
    InMux I__10964 (
            .O(N__50646),
            .I(N__50578));
    LocalMux I__10963 (
            .O(N__50643),
            .I(N__50567));
    LocalMux I__10962 (
            .O(N__50640),
            .I(N__50567));
    LocalMux I__10961 (
            .O(N__50637),
            .I(N__50567));
    LocalMux I__10960 (
            .O(N__50632),
            .I(N__50567));
    LocalMux I__10959 (
            .O(N__50629),
            .I(N__50567));
    LocalMux I__10958 (
            .O(N__50622),
            .I(N__50564));
    InMux I__10957 (
            .O(N__50621),
            .I(N__50561));
    InMux I__10956 (
            .O(N__50620),
            .I(N__50558));
    LocalMux I__10955 (
            .O(N__50617),
            .I(N__50553));
    LocalMux I__10954 (
            .O(N__50612),
            .I(N__50553));
    InMux I__10953 (
            .O(N__50611),
            .I(N__50546));
    InMux I__10952 (
            .O(N__50610),
            .I(N__50546));
    InMux I__10951 (
            .O(N__50609),
            .I(N__50546));
    LocalMux I__10950 (
            .O(N__50606),
            .I(N__50541));
    LocalMux I__10949 (
            .O(N__50601),
            .I(N__50541));
    Span4Mux_h I__10948 (
            .O(N__50596),
            .I(N__50538));
    InMux I__10947 (
            .O(N__50595),
            .I(N__50532));
    InMux I__10946 (
            .O(N__50594),
            .I(N__50532));
    LocalMux I__10945 (
            .O(N__50591),
            .I(N__50527));
    LocalMux I__10944 (
            .O(N__50588),
            .I(N__50527));
    LocalMux I__10943 (
            .O(N__50583),
            .I(N__50520));
    LocalMux I__10942 (
            .O(N__50578),
            .I(N__50520));
    Span4Mux_v I__10941 (
            .O(N__50567),
            .I(N__50520));
    Span4Mux_h I__10940 (
            .O(N__50564),
            .I(N__50517));
    LocalMux I__10939 (
            .O(N__50561),
            .I(N__50512));
    LocalMux I__10938 (
            .O(N__50558),
            .I(N__50512));
    Span12Mux_s7_v I__10937 (
            .O(N__50553),
            .I(N__50507));
    LocalMux I__10936 (
            .O(N__50546),
            .I(N__50507));
    Span4Mux_h I__10935 (
            .O(N__50541),
            .I(N__50504));
    Span4Mux_v I__10934 (
            .O(N__50538),
            .I(N__50501));
    InMux I__10933 (
            .O(N__50537),
            .I(N__50495));
    LocalMux I__10932 (
            .O(N__50532),
            .I(N__50486));
    Span4Mux_v I__10931 (
            .O(N__50527),
            .I(N__50486));
    Span4Mux_v I__10930 (
            .O(N__50520),
            .I(N__50486));
    Span4Mux_v I__10929 (
            .O(N__50517),
            .I(N__50486));
    Span12Mux_v I__10928 (
            .O(N__50512),
            .I(N__50481));
    Span12Mux_v I__10927 (
            .O(N__50507),
            .I(N__50481));
    Span4Mux_v I__10926 (
            .O(N__50504),
            .I(N__50478));
    Sp12to4 I__10925 (
            .O(N__50501),
            .I(N__50475));
    InMux I__10924 (
            .O(N__50500),
            .I(N__50468));
    InMux I__10923 (
            .O(N__50499),
            .I(N__50468));
    InMux I__10922 (
            .O(N__50498),
            .I(N__50468));
    LocalMux I__10921 (
            .O(N__50495),
            .I(\c0.n31_adj_4271 ));
    Odrv4 I__10920 (
            .O(N__50486),
            .I(\c0.n31_adj_4271 ));
    Odrv12 I__10919 (
            .O(N__50481),
            .I(\c0.n31_adj_4271 ));
    Odrv4 I__10918 (
            .O(N__50478),
            .I(\c0.n31_adj_4271 ));
    Odrv12 I__10917 (
            .O(N__50475),
            .I(\c0.n31_adj_4271 ));
    LocalMux I__10916 (
            .O(N__50468),
            .I(\c0.n31_adj_4271 ));
    SRMux I__10915 (
            .O(N__50455),
            .I(N__50452));
    LocalMux I__10914 (
            .O(N__50452),
            .I(N__50449));
    Span4Mux_h I__10913 (
            .O(N__50449),
            .I(N__50446));
    Odrv4 I__10912 (
            .O(N__50446),
            .I(\c0.n3_adj_4430 ));
    InMux I__10911 (
            .O(N__50443),
            .I(N__50440));
    LocalMux I__10910 (
            .O(N__50440),
            .I(N__50435));
    InMux I__10909 (
            .O(N__50439),
            .I(N__50432));
    InMux I__10908 (
            .O(N__50438),
            .I(N__50429));
    Span4Mux_v I__10907 (
            .O(N__50435),
            .I(N__50426));
    LocalMux I__10906 (
            .O(N__50432),
            .I(N__50423));
    LocalMux I__10905 (
            .O(N__50429),
            .I(\c0.data_in_frame_7_4 ));
    Odrv4 I__10904 (
            .O(N__50426),
            .I(\c0.data_in_frame_7_4 ));
    Odrv12 I__10903 (
            .O(N__50423),
            .I(\c0.data_in_frame_7_4 ));
    CascadeMux I__10902 (
            .O(N__50416),
            .I(\c0.n13555_cascade_ ));
    InMux I__10901 (
            .O(N__50413),
            .I(N__50410));
    LocalMux I__10900 (
            .O(N__50410),
            .I(N__50407));
    Span4Mux_h I__10899 (
            .O(N__50407),
            .I(N__50404));
    Span4Mux_v I__10898 (
            .O(N__50404),
            .I(N__50400));
    InMux I__10897 (
            .O(N__50403),
            .I(N__50397));
    Odrv4 I__10896 (
            .O(N__50400),
            .I(\c0.n13555 ));
    LocalMux I__10895 (
            .O(N__50397),
            .I(\c0.n13555 ));
    CascadeMux I__10894 (
            .O(N__50392),
            .I(\c0.n22043_cascade_ ));
    InMux I__10893 (
            .O(N__50389),
            .I(N__50385));
    InMux I__10892 (
            .O(N__50388),
            .I(N__50382));
    LocalMux I__10891 (
            .O(N__50385),
            .I(N__50378));
    LocalMux I__10890 (
            .O(N__50382),
            .I(N__50375));
    InMux I__10889 (
            .O(N__50381),
            .I(N__50372));
    Span4Mux_h I__10888 (
            .O(N__50378),
            .I(N__50369));
    Span4Mux_v I__10887 (
            .O(N__50375),
            .I(N__50365));
    LocalMux I__10886 (
            .O(N__50372),
            .I(N__50360));
    Span4Mux_v I__10885 (
            .O(N__50369),
            .I(N__50360));
    InMux I__10884 (
            .O(N__50368),
            .I(N__50357));
    Odrv4 I__10883 (
            .O(N__50365),
            .I(\c0.data_in_frame_2_6 ));
    Odrv4 I__10882 (
            .O(N__50360),
            .I(\c0.data_in_frame_2_6 ));
    LocalMux I__10881 (
            .O(N__50357),
            .I(\c0.data_in_frame_2_6 ));
    InMux I__10880 (
            .O(N__50350),
            .I(N__50346));
    InMux I__10879 (
            .O(N__50349),
            .I(N__50342));
    LocalMux I__10878 (
            .O(N__50346),
            .I(N__50336));
    InMux I__10877 (
            .O(N__50345),
            .I(N__50333));
    LocalMux I__10876 (
            .O(N__50342),
            .I(N__50330));
    InMux I__10875 (
            .O(N__50341),
            .I(N__50325));
    InMux I__10874 (
            .O(N__50340),
            .I(N__50325));
    InMux I__10873 (
            .O(N__50339),
            .I(N__50322));
    Span4Mux_h I__10872 (
            .O(N__50336),
            .I(N__50318));
    LocalMux I__10871 (
            .O(N__50333),
            .I(N__50315));
    Span4Mux_v I__10870 (
            .O(N__50330),
            .I(N__50308));
    LocalMux I__10869 (
            .O(N__50325),
            .I(N__50308));
    LocalMux I__10868 (
            .O(N__50322),
            .I(N__50308));
    InMux I__10867 (
            .O(N__50321),
            .I(N__50303));
    Span4Mux_v I__10866 (
            .O(N__50318),
            .I(N__50300));
    Span4Mux_v I__10865 (
            .O(N__50315),
            .I(N__50295));
    Span4Mux_h I__10864 (
            .O(N__50308),
            .I(N__50295));
    InMux I__10863 (
            .O(N__50307),
            .I(N__50290));
    InMux I__10862 (
            .O(N__50306),
            .I(N__50290));
    LocalMux I__10861 (
            .O(N__50303),
            .I(\c0.data_in_frame_0_4 ));
    Odrv4 I__10860 (
            .O(N__50300),
            .I(\c0.data_in_frame_0_4 ));
    Odrv4 I__10859 (
            .O(N__50295),
            .I(\c0.data_in_frame_0_4 ));
    LocalMux I__10858 (
            .O(N__50290),
            .I(\c0.data_in_frame_0_4 ));
    CascadeMux I__10857 (
            .O(N__50281),
            .I(N__50278));
    InMux I__10856 (
            .O(N__50278),
            .I(N__50275));
    LocalMux I__10855 (
            .O(N__50275),
            .I(N__50272));
    Odrv12 I__10854 (
            .O(N__50272),
            .I(\c0.n10_adj_4363 ));
    CascadeMux I__10853 (
            .O(N__50269),
            .I(\c0.rx.n22573_cascade_ ));
    CascadeMux I__10852 (
            .O(N__50266),
            .I(\c0.rx.n12_cascade_ ));
    InMux I__10851 (
            .O(N__50263),
            .I(bfn_20_24_0_));
    InMux I__10850 (
            .O(N__50260),
            .I(N__50256));
    InMux I__10849 (
            .O(N__50259),
            .I(N__50253));
    LocalMux I__10848 (
            .O(N__50256),
            .I(\c0.rx.r_Clock_Count_1 ));
    LocalMux I__10847 (
            .O(N__50253),
            .I(\c0.rx.r_Clock_Count_1 ));
    InMux I__10846 (
            .O(N__50248),
            .I(\c0.rx.n19533 ));
    InMux I__10845 (
            .O(N__50245),
            .I(N__50241));
    InMux I__10844 (
            .O(N__50244),
            .I(N__50238));
    LocalMux I__10843 (
            .O(N__50241),
            .I(\c0.rx.r_Clock_Count_2 ));
    LocalMux I__10842 (
            .O(N__50238),
            .I(\c0.rx.r_Clock_Count_2 ));
    InMux I__10841 (
            .O(N__50233),
            .I(\c0.rx.n19534 ));
    InMux I__10840 (
            .O(N__50230),
            .I(N__50226));
    InMux I__10839 (
            .O(N__50229),
            .I(N__50223));
    LocalMux I__10838 (
            .O(N__50226),
            .I(\c0.rx.r_Clock_Count_3 ));
    LocalMux I__10837 (
            .O(N__50223),
            .I(\c0.rx.r_Clock_Count_3 ));
    InMux I__10836 (
            .O(N__50218),
            .I(\c0.rx.n19535 ));
    InMux I__10835 (
            .O(N__50215),
            .I(\c0.rx.n19536 ));
    InMux I__10834 (
            .O(N__50212),
            .I(\c0.rx.n19537 ));
    InMux I__10833 (
            .O(N__50209),
            .I(\c0.rx.n19538 ));
    InMux I__10832 (
            .O(N__50206),
            .I(N__50201));
    InMux I__10831 (
            .O(N__50205),
            .I(N__50198));
    InMux I__10830 (
            .O(N__50204),
            .I(N__50195));
    LocalMux I__10829 (
            .O(N__50201),
            .I(N__50192));
    LocalMux I__10828 (
            .O(N__50198),
            .I(N__50186));
    LocalMux I__10827 (
            .O(N__50195),
            .I(N__50186));
    Span4Mux_h I__10826 (
            .O(N__50192),
            .I(N__50183));
    InMux I__10825 (
            .O(N__50191),
            .I(N__50180));
    Span4Mux_h I__10824 (
            .O(N__50186),
            .I(N__50177));
    Span4Mux_v I__10823 (
            .O(N__50183),
            .I(N__50174));
    LocalMux I__10822 (
            .O(N__50180),
            .I(\c0.data_in_frame_27_1 ));
    Odrv4 I__10821 (
            .O(N__50177),
            .I(\c0.data_in_frame_27_1 ));
    Odrv4 I__10820 (
            .O(N__50174),
            .I(\c0.data_in_frame_27_1 ));
    CascadeMux I__10819 (
            .O(N__50167),
            .I(N__50164));
    InMux I__10818 (
            .O(N__50164),
            .I(N__50161));
    LocalMux I__10817 (
            .O(N__50161),
            .I(N__50158));
    Span4Mux_v I__10816 (
            .O(N__50158),
            .I(N__50154));
    InMux I__10815 (
            .O(N__50157),
            .I(N__50151));
    Span4Mux_v I__10814 (
            .O(N__50154),
            .I(N__50148));
    LocalMux I__10813 (
            .O(N__50151),
            .I(N__50145));
    Span4Mux_v I__10812 (
            .O(N__50148),
            .I(N__50142));
    Span4Mux_v I__10811 (
            .O(N__50145),
            .I(N__50139));
    Span4Mux_v I__10810 (
            .O(N__50142),
            .I(N__50135));
    Span4Mux_v I__10809 (
            .O(N__50139),
            .I(N__50132));
    InMux I__10808 (
            .O(N__50138),
            .I(N__50129));
    Odrv4 I__10807 (
            .O(N__50135),
            .I(\c0.FRAME_MATCHER_i_10 ));
    Odrv4 I__10806 (
            .O(N__50132),
            .I(\c0.FRAME_MATCHER_i_10 ));
    LocalMux I__10805 (
            .O(N__50129),
            .I(\c0.FRAME_MATCHER_i_10 ));
    SRMux I__10804 (
            .O(N__50122),
            .I(N__50119));
    LocalMux I__10803 (
            .O(N__50119),
            .I(N__50116));
    Span4Mux_v I__10802 (
            .O(N__50116),
            .I(N__50113));
    Sp12to4 I__10801 (
            .O(N__50113),
            .I(N__50110));
    Odrv12 I__10800 (
            .O(N__50110),
            .I(\c0.n3_adj_4460 ));
    InMux I__10799 (
            .O(N__50107),
            .I(N__50103));
    InMux I__10798 (
            .O(N__50106),
            .I(N__50100));
    LocalMux I__10797 (
            .O(N__50103),
            .I(N__50097));
    LocalMux I__10796 (
            .O(N__50100),
            .I(N__50094));
    Span4Mux_v I__10795 (
            .O(N__50097),
            .I(N__50091));
    Span12Mux_h I__10794 (
            .O(N__50094),
            .I(N__50088));
    Span4Mux_v I__10793 (
            .O(N__50091),
            .I(N__50085));
    Odrv12 I__10792 (
            .O(N__50088),
            .I(n18678));
    Odrv4 I__10791 (
            .O(N__50085),
            .I(n18678));
    CascadeMux I__10790 (
            .O(N__50080),
            .I(\c0.rx.n18655_cascade_ ));
    CascadeMux I__10789 (
            .O(N__50077),
            .I(\c0.rx.n21704_cascade_ ));
    InMux I__10788 (
            .O(N__50074),
            .I(N__50065));
    InMux I__10787 (
            .O(N__50073),
            .I(N__50065));
    InMux I__10786 (
            .O(N__50072),
            .I(N__50065));
    LocalMux I__10785 (
            .O(N__50065),
            .I(\c0.data_in_frame_23_4 ));
    CascadeMux I__10784 (
            .O(N__50062),
            .I(\c0.n10_adj_4287_cascade_ ));
    InMux I__10783 (
            .O(N__50059),
            .I(N__50056));
    LocalMux I__10782 (
            .O(N__50056),
            .I(N__50053));
    Span4Mux_h I__10781 (
            .O(N__50053),
            .I(N__50050));
    Odrv4 I__10780 (
            .O(N__50050),
            .I(\c0.n22_adj_4298 ));
    InMux I__10779 (
            .O(N__50047),
            .I(N__50044));
    LocalMux I__10778 (
            .O(N__50044),
            .I(N__50041));
    Odrv4 I__10777 (
            .O(N__50041),
            .I(\c0.n13266 ));
    InMux I__10776 (
            .O(N__50038),
            .I(N__50035));
    LocalMux I__10775 (
            .O(N__50035),
            .I(N__50031));
    InMux I__10774 (
            .O(N__50034),
            .I(N__50028));
    Span4Mux_h I__10773 (
            .O(N__50031),
            .I(N__50025));
    LocalMux I__10772 (
            .O(N__50028),
            .I(\c0.data_in_frame_29_7 ));
    Odrv4 I__10771 (
            .O(N__50025),
            .I(\c0.data_in_frame_29_7 ));
    CascadeMux I__10770 (
            .O(N__50020),
            .I(\c0.n21233_cascade_ ));
    InMux I__10769 (
            .O(N__50017),
            .I(N__50014));
    LocalMux I__10768 (
            .O(N__50014),
            .I(\c0.n23506 ));
    CascadeMux I__10767 (
            .O(N__50011),
            .I(N__50007));
    CascadeMux I__10766 (
            .O(N__50010),
            .I(N__50004));
    InMux I__10765 (
            .O(N__50007),
            .I(N__50001));
    InMux I__10764 (
            .O(N__50004),
            .I(N__49998));
    LocalMux I__10763 (
            .O(N__50001),
            .I(N__49993));
    LocalMux I__10762 (
            .O(N__49998),
            .I(N__49993));
    Span4Mux_h I__10761 (
            .O(N__49993),
            .I(N__49989));
    InMux I__10760 (
            .O(N__49992),
            .I(N__49986));
    Odrv4 I__10759 (
            .O(N__49989),
            .I(\c0.FRAME_MATCHER_i_20 ));
    LocalMux I__10758 (
            .O(N__49986),
            .I(\c0.FRAME_MATCHER_i_20 ));
    SRMux I__10757 (
            .O(N__49981),
            .I(N__49978));
    LocalMux I__10756 (
            .O(N__49978),
            .I(N__49975));
    Span4Mux_v I__10755 (
            .O(N__49975),
            .I(N__49972));
    Odrv4 I__10754 (
            .O(N__49972),
            .I(\c0.n3_adj_4442 ));
    CascadeMux I__10753 (
            .O(N__49969),
            .I(N__49966));
    InMux I__10752 (
            .O(N__49966),
            .I(N__49963));
    LocalMux I__10751 (
            .O(N__49963),
            .I(N__49959));
    CascadeMux I__10750 (
            .O(N__49962),
            .I(N__49956));
    Span4Mux_h I__10749 (
            .O(N__49959),
            .I(N__49953));
    InMux I__10748 (
            .O(N__49956),
            .I(N__49950));
    Span4Mux_h I__10747 (
            .O(N__49953),
            .I(N__49947));
    LocalMux I__10746 (
            .O(N__49950),
            .I(\c0.data_in_frame_28_1 ));
    Odrv4 I__10745 (
            .O(N__49947),
            .I(\c0.data_in_frame_28_1 ));
    CascadeMux I__10744 (
            .O(N__49942),
            .I(\c0.n21870_cascade_ ));
    CascadeMux I__10743 (
            .O(N__49939),
            .I(N__49936));
    InMux I__10742 (
            .O(N__49936),
            .I(N__49931));
    InMux I__10741 (
            .O(N__49935),
            .I(N__49926));
    InMux I__10740 (
            .O(N__49934),
            .I(N__49926));
    LocalMux I__10739 (
            .O(N__49931),
            .I(\c0.data_in_frame_21_3 ));
    LocalMux I__10738 (
            .O(N__49926),
            .I(\c0.data_in_frame_21_3 ));
    InMux I__10737 (
            .O(N__49921),
            .I(N__49916));
    InMux I__10736 (
            .O(N__49920),
            .I(N__49913));
    InMux I__10735 (
            .O(N__49919),
            .I(N__49910));
    LocalMux I__10734 (
            .O(N__49916),
            .I(N__49905));
    LocalMux I__10733 (
            .O(N__49913),
            .I(N__49905));
    LocalMux I__10732 (
            .O(N__49910),
            .I(\c0.data_in_frame_23_5 ));
    Odrv4 I__10731 (
            .O(N__49905),
            .I(\c0.data_in_frame_23_5 ));
    CascadeMux I__10730 (
            .O(N__49900),
            .I(\c0.n21858_cascade_ ));
    CascadeMux I__10729 (
            .O(N__49897),
            .I(N__49894));
    InMux I__10728 (
            .O(N__49894),
            .I(N__49891));
    LocalMux I__10727 (
            .O(N__49891),
            .I(N__49886));
    InMux I__10726 (
            .O(N__49890),
            .I(N__49883));
    InMux I__10725 (
            .O(N__49889),
            .I(N__49880));
    Odrv4 I__10724 (
            .O(N__49886),
            .I(\c0.FRAME_MATCHER_i_16 ));
    LocalMux I__10723 (
            .O(N__49883),
            .I(\c0.FRAME_MATCHER_i_16 ));
    LocalMux I__10722 (
            .O(N__49880),
            .I(\c0.FRAME_MATCHER_i_16 ));
    InMux I__10721 (
            .O(N__49873),
            .I(N__49870));
    LocalMux I__10720 (
            .O(N__49870),
            .I(N__49867));
    Span4Mux_v I__10719 (
            .O(N__49867),
            .I(N__49864));
    Odrv4 I__10718 (
            .O(N__49864),
            .I(\c0.n16_adj_4375 ));
    CascadeMux I__10717 (
            .O(N__49861),
            .I(N__49858));
    InMux I__10716 (
            .O(N__49858),
            .I(N__49852));
    InMux I__10715 (
            .O(N__49857),
            .I(N__49852));
    LocalMux I__10714 (
            .O(N__49852),
            .I(N__49848));
    InMux I__10713 (
            .O(N__49851),
            .I(N__49845));
    Span4Mux_v I__10712 (
            .O(N__49848),
            .I(N__49842));
    LocalMux I__10711 (
            .O(N__49845),
            .I(\c0.FRAME_MATCHER_i_13 ));
    Odrv4 I__10710 (
            .O(N__49842),
            .I(\c0.FRAME_MATCHER_i_13 ));
    SRMux I__10709 (
            .O(N__49837),
            .I(N__49834));
    LocalMux I__10708 (
            .O(N__49834),
            .I(N__49831));
    Span4Mux_h I__10707 (
            .O(N__49831),
            .I(N__49828));
    Span4Mux_h I__10706 (
            .O(N__49828),
            .I(N__49825));
    Odrv4 I__10705 (
            .O(N__49825),
            .I(\c0.n3_adj_4454 ));
    InMux I__10704 (
            .O(N__49822),
            .I(N__49818));
    InMux I__10703 (
            .O(N__49821),
            .I(N__49815));
    LocalMux I__10702 (
            .O(N__49818),
            .I(N__49811));
    LocalMux I__10701 (
            .O(N__49815),
            .I(N__49808));
    InMux I__10700 (
            .O(N__49814),
            .I(N__49805));
    Span4Mux_v I__10699 (
            .O(N__49811),
            .I(N__49802));
    Odrv4 I__10698 (
            .O(N__49808),
            .I(\c0.FRAME_MATCHER_i_15 ));
    LocalMux I__10697 (
            .O(N__49805),
            .I(\c0.FRAME_MATCHER_i_15 ));
    Odrv4 I__10696 (
            .O(N__49802),
            .I(\c0.FRAME_MATCHER_i_15 ));
    SRMux I__10695 (
            .O(N__49795),
            .I(N__49792));
    LocalMux I__10694 (
            .O(N__49792),
            .I(N__49789));
    Span4Mux_h I__10693 (
            .O(N__49789),
            .I(N__49786));
    Odrv4 I__10692 (
            .O(N__49786),
            .I(\c0.n3_adj_4452 ));
    InMux I__10691 (
            .O(N__49783),
            .I(N__49780));
    LocalMux I__10690 (
            .O(N__49780),
            .I(N__49776));
    InMux I__10689 (
            .O(N__49779),
            .I(N__49773));
    Span4Mux_v I__10688 (
            .O(N__49776),
            .I(N__49768));
    LocalMux I__10687 (
            .O(N__49773),
            .I(N__49768));
    Span4Mux_v I__10686 (
            .O(N__49768),
            .I(N__49765));
    Odrv4 I__10685 (
            .O(N__49765),
            .I(\c0.n13697 ));
    CascadeMux I__10684 (
            .O(N__49762),
            .I(\c0.n22440_cascade_ ));
    InMux I__10683 (
            .O(N__49759),
            .I(N__49756));
    LocalMux I__10682 (
            .O(N__49756),
            .I(N__49750));
    InMux I__10681 (
            .O(N__49755),
            .I(N__49745));
    InMux I__10680 (
            .O(N__49754),
            .I(N__49745));
    CascadeMux I__10679 (
            .O(N__49753),
            .I(N__49742));
    Span4Mux_v I__10678 (
            .O(N__49750),
            .I(N__49737));
    LocalMux I__10677 (
            .O(N__49745),
            .I(N__49737));
    InMux I__10676 (
            .O(N__49742),
            .I(N__49733));
    Span4Mux_v I__10675 (
            .O(N__49737),
            .I(N__49730));
    InMux I__10674 (
            .O(N__49736),
            .I(N__49727));
    LocalMux I__10673 (
            .O(N__49733),
            .I(\c0.data_in_frame_10_7 ));
    Odrv4 I__10672 (
            .O(N__49730),
            .I(\c0.data_in_frame_10_7 ));
    LocalMux I__10671 (
            .O(N__49727),
            .I(\c0.data_in_frame_10_7 ));
    CascadeMux I__10670 (
            .O(N__49720),
            .I(\c0.n10_adj_4229_cascade_ ));
    CascadeMux I__10669 (
            .O(N__49717),
            .I(\c0.n5943_cascade_ ));
    CascadeMux I__10668 (
            .O(N__49714),
            .I(\c0.n22081_cascade_ ));
    CascadeMux I__10667 (
            .O(N__49711),
            .I(\c0.n22349_cascade_ ));
    InMux I__10666 (
            .O(N__49708),
            .I(N__49704));
    InMux I__10665 (
            .O(N__49707),
            .I(N__49700));
    LocalMux I__10664 (
            .O(N__49704),
            .I(N__49697));
    InMux I__10663 (
            .O(N__49703),
            .I(N__49694));
    LocalMux I__10662 (
            .O(N__49700),
            .I(N__49688));
    Span4Mux_v I__10661 (
            .O(N__49697),
            .I(N__49683));
    LocalMux I__10660 (
            .O(N__49694),
            .I(N__49683));
    InMux I__10659 (
            .O(N__49693),
            .I(N__49680));
    InMux I__10658 (
            .O(N__49692),
            .I(N__49675));
    InMux I__10657 (
            .O(N__49691),
            .I(N__49675));
    Span4Mux_v I__10656 (
            .O(N__49688),
            .I(N__49669));
    Span4Mux_h I__10655 (
            .O(N__49683),
            .I(N__49669));
    LocalMux I__10654 (
            .O(N__49680),
            .I(N__49664));
    LocalMux I__10653 (
            .O(N__49675),
            .I(N__49664));
    InMux I__10652 (
            .O(N__49674),
            .I(N__49661));
    Odrv4 I__10651 (
            .O(N__49669),
            .I(n21744));
    Odrv12 I__10650 (
            .O(N__49664),
            .I(n21744));
    LocalMux I__10649 (
            .O(N__49661),
            .I(n21744));
    InMux I__10648 (
            .O(N__49654),
            .I(N__49651));
    LocalMux I__10647 (
            .O(N__49651),
            .I(N__49648));
    Span4Mux_h I__10646 (
            .O(N__49648),
            .I(N__49645));
    Odrv4 I__10645 (
            .O(N__49645),
            .I(\c0.n6_adj_4386 ));
    CascadeMux I__10644 (
            .O(N__49642),
            .I(N__49638));
    InMux I__10643 (
            .O(N__49641),
            .I(N__49635));
    InMux I__10642 (
            .O(N__49638),
            .I(N__49631));
    LocalMux I__10641 (
            .O(N__49635),
            .I(N__49628));
    InMux I__10640 (
            .O(N__49634),
            .I(N__49625));
    LocalMux I__10639 (
            .O(N__49631),
            .I(N__49622));
    Span4Mux_h I__10638 (
            .O(N__49628),
            .I(N__49619));
    LocalMux I__10637 (
            .O(N__49625),
            .I(N__49616));
    Odrv12 I__10636 (
            .O(N__49622),
            .I(\c0.data_in_frame_4_3 ));
    Odrv4 I__10635 (
            .O(N__49619),
            .I(\c0.data_in_frame_4_3 ));
    Odrv12 I__10634 (
            .O(N__49616),
            .I(\c0.data_in_frame_4_3 ));
    CascadeMux I__10633 (
            .O(N__49609),
            .I(N__49605));
    InMux I__10632 (
            .O(N__49608),
            .I(N__49600));
    InMux I__10631 (
            .O(N__49605),
            .I(N__49600));
    LocalMux I__10630 (
            .O(N__49600),
            .I(data_in_frame_6_4));
    InMux I__10629 (
            .O(N__49597),
            .I(N__49593));
    CascadeMux I__10628 (
            .O(N__49596),
            .I(N__49590));
    LocalMux I__10627 (
            .O(N__49593),
            .I(N__49586));
    InMux I__10626 (
            .O(N__49590),
            .I(N__49581));
    InMux I__10625 (
            .O(N__49589),
            .I(N__49581));
    Span4Mux_h I__10624 (
            .O(N__49586),
            .I(N__49578));
    LocalMux I__10623 (
            .O(N__49581),
            .I(N__49573));
    Span4Mux_v I__10622 (
            .O(N__49578),
            .I(N__49573));
    Odrv4 I__10621 (
            .O(N__49573),
            .I(\c0.data_in_frame_4_2 ));
    InMux I__10620 (
            .O(N__49570),
            .I(N__49566));
    InMux I__10619 (
            .O(N__49569),
            .I(N__49562));
    LocalMux I__10618 (
            .O(N__49566),
            .I(N__49558));
    InMux I__10617 (
            .O(N__49565),
            .I(N__49555));
    LocalMux I__10616 (
            .O(N__49562),
            .I(N__49545));
    InMux I__10615 (
            .O(N__49561),
            .I(N__49542));
    Span4Mux_h I__10614 (
            .O(N__49558),
            .I(N__49539));
    LocalMux I__10613 (
            .O(N__49555),
            .I(N__49536));
    InMux I__10612 (
            .O(N__49554),
            .I(N__49531));
    InMux I__10611 (
            .O(N__49553),
            .I(N__49531));
    CascadeMux I__10610 (
            .O(N__49552),
            .I(N__49528));
    CascadeMux I__10609 (
            .O(N__49551),
            .I(N__49525));
    InMux I__10608 (
            .O(N__49550),
            .I(N__49520));
    InMux I__10607 (
            .O(N__49549),
            .I(N__49520));
    InMux I__10606 (
            .O(N__49548),
            .I(N__49514));
    Span4Mux_v I__10605 (
            .O(N__49545),
            .I(N__49501));
    LocalMux I__10604 (
            .O(N__49542),
            .I(N__49501));
    Span4Mux_h I__10603 (
            .O(N__49539),
            .I(N__49501));
    Span4Mux_h I__10602 (
            .O(N__49536),
            .I(N__49501));
    LocalMux I__10601 (
            .O(N__49531),
            .I(N__49501));
    InMux I__10600 (
            .O(N__49528),
            .I(N__49496));
    InMux I__10599 (
            .O(N__49525),
            .I(N__49496));
    LocalMux I__10598 (
            .O(N__49520),
            .I(N__49493));
    InMux I__10597 (
            .O(N__49519),
            .I(N__49488));
    InMux I__10596 (
            .O(N__49518),
            .I(N__49488));
    InMux I__10595 (
            .O(N__49517),
            .I(N__49485));
    LocalMux I__10594 (
            .O(N__49514),
            .I(N__49482));
    InMux I__10593 (
            .O(N__49513),
            .I(N__49477));
    InMux I__10592 (
            .O(N__49512),
            .I(N__49477));
    Span4Mux_v I__10591 (
            .O(N__49501),
            .I(N__49457));
    LocalMux I__10590 (
            .O(N__49496),
            .I(N__49457));
    Span4Mux_h I__10589 (
            .O(N__49493),
            .I(N__49457));
    LocalMux I__10588 (
            .O(N__49488),
            .I(N__49457));
    LocalMux I__10587 (
            .O(N__49485),
            .I(N__49457));
    Span4Mux_h I__10586 (
            .O(N__49482),
            .I(N__49457));
    LocalMux I__10585 (
            .O(N__49477),
            .I(N__49457));
    InMux I__10584 (
            .O(N__49476),
            .I(N__49438));
    InMux I__10583 (
            .O(N__49475),
            .I(N__49438));
    InMux I__10582 (
            .O(N__49474),
            .I(N__49431));
    InMux I__10581 (
            .O(N__49473),
            .I(N__49431));
    InMux I__10580 (
            .O(N__49472),
            .I(N__49431));
    Span4Mux_v I__10579 (
            .O(N__49457),
            .I(N__49428));
    InMux I__10578 (
            .O(N__49456),
            .I(N__49416));
    InMux I__10577 (
            .O(N__49455),
            .I(N__49416));
    InMux I__10576 (
            .O(N__49454),
            .I(N__49416));
    InMux I__10575 (
            .O(N__49453),
            .I(N__49416));
    CascadeMux I__10574 (
            .O(N__49452),
            .I(N__49407));
    CascadeMux I__10573 (
            .O(N__49451),
            .I(N__49404));
    InMux I__10572 (
            .O(N__49450),
            .I(N__49397));
    InMux I__10571 (
            .O(N__49449),
            .I(N__49397));
    InMux I__10570 (
            .O(N__49448),
            .I(N__49394));
    InMux I__10569 (
            .O(N__49447),
            .I(N__49386));
    InMux I__10568 (
            .O(N__49446),
            .I(N__49386));
    InMux I__10567 (
            .O(N__49445),
            .I(N__49383));
    InMux I__10566 (
            .O(N__49444),
            .I(N__49374));
    InMux I__10565 (
            .O(N__49443),
            .I(N__49374));
    LocalMux I__10564 (
            .O(N__49438),
            .I(N__49371));
    LocalMux I__10563 (
            .O(N__49431),
            .I(N__49366));
    Span4Mux_h I__10562 (
            .O(N__49428),
            .I(N__49366));
    InMux I__10561 (
            .O(N__49427),
            .I(N__49359));
    InMux I__10560 (
            .O(N__49426),
            .I(N__49359));
    InMux I__10559 (
            .O(N__49425),
            .I(N__49359));
    LocalMux I__10558 (
            .O(N__49416),
            .I(N__49353));
    InMux I__10557 (
            .O(N__49415),
            .I(N__49348));
    InMux I__10556 (
            .O(N__49414),
            .I(N__49348));
    InMux I__10555 (
            .O(N__49413),
            .I(N__49345));
    InMux I__10554 (
            .O(N__49412),
            .I(N__49340));
    InMux I__10553 (
            .O(N__49411),
            .I(N__49340));
    InMux I__10552 (
            .O(N__49410),
            .I(N__49337));
    InMux I__10551 (
            .O(N__49407),
            .I(N__49326));
    InMux I__10550 (
            .O(N__49404),
            .I(N__49326));
    InMux I__10549 (
            .O(N__49403),
            .I(N__49323));
    InMux I__10548 (
            .O(N__49402),
            .I(N__49317));
    LocalMux I__10547 (
            .O(N__49397),
            .I(N__49314));
    LocalMux I__10546 (
            .O(N__49394),
            .I(N__49311));
    InMux I__10545 (
            .O(N__49393),
            .I(N__49304));
    InMux I__10544 (
            .O(N__49392),
            .I(N__49304));
    InMux I__10543 (
            .O(N__49391),
            .I(N__49304));
    LocalMux I__10542 (
            .O(N__49386),
            .I(N__49299));
    LocalMux I__10541 (
            .O(N__49383),
            .I(N__49299));
    InMux I__10540 (
            .O(N__49382),
            .I(N__49292));
    InMux I__10539 (
            .O(N__49381),
            .I(N__49292));
    InMux I__10538 (
            .O(N__49380),
            .I(N__49292));
    InMux I__10537 (
            .O(N__49379),
            .I(N__49289));
    LocalMux I__10536 (
            .O(N__49374),
            .I(N__49280));
    Span4Mux_h I__10535 (
            .O(N__49371),
            .I(N__49280));
    Span4Mux_h I__10534 (
            .O(N__49366),
            .I(N__49280));
    LocalMux I__10533 (
            .O(N__49359),
            .I(N__49280));
    InMux I__10532 (
            .O(N__49358),
            .I(N__49275));
    InMux I__10531 (
            .O(N__49357),
            .I(N__49275));
    InMux I__10530 (
            .O(N__49356),
            .I(N__49266));
    Span4Mux_h I__10529 (
            .O(N__49353),
            .I(N__49261));
    LocalMux I__10528 (
            .O(N__49348),
            .I(N__49261));
    LocalMux I__10527 (
            .O(N__49345),
            .I(N__49256));
    LocalMux I__10526 (
            .O(N__49340),
            .I(N__49256));
    LocalMux I__10525 (
            .O(N__49337),
            .I(N__49250));
    InMux I__10524 (
            .O(N__49336),
            .I(N__49243));
    InMux I__10523 (
            .O(N__49335),
            .I(N__49243));
    InMux I__10522 (
            .O(N__49334),
            .I(N__49243));
    InMux I__10521 (
            .O(N__49333),
            .I(N__49236));
    InMux I__10520 (
            .O(N__49332),
            .I(N__49236));
    InMux I__10519 (
            .O(N__49331),
            .I(N__49236));
    LocalMux I__10518 (
            .O(N__49326),
            .I(N__49231));
    LocalMux I__10517 (
            .O(N__49323),
            .I(N__49231));
    InMux I__10516 (
            .O(N__49322),
            .I(N__49228));
    InMux I__10515 (
            .O(N__49321),
            .I(N__49223));
    InMux I__10514 (
            .O(N__49320),
            .I(N__49223));
    LocalMux I__10513 (
            .O(N__49317),
            .I(N__49212));
    Span4Mux_h I__10512 (
            .O(N__49314),
            .I(N__49212));
    Span4Mux_h I__10511 (
            .O(N__49311),
            .I(N__49212));
    LocalMux I__10510 (
            .O(N__49304),
            .I(N__49212));
    Span4Mux_h I__10509 (
            .O(N__49299),
            .I(N__49212));
    LocalMux I__10508 (
            .O(N__49292),
            .I(N__49207));
    LocalMux I__10507 (
            .O(N__49289),
            .I(N__49207));
    Span4Mux_v I__10506 (
            .O(N__49280),
            .I(N__49204));
    LocalMux I__10505 (
            .O(N__49275),
            .I(N__49198));
    InMux I__10504 (
            .O(N__49274),
            .I(N__49193));
    InMux I__10503 (
            .O(N__49273),
            .I(N__49193));
    InMux I__10502 (
            .O(N__49272),
            .I(N__49190));
    InMux I__10501 (
            .O(N__49271),
            .I(N__49183));
    InMux I__10500 (
            .O(N__49270),
            .I(N__49183));
    InMux I__10499 (
            .O(N__49269),
            .I(N__49183));
    LocalMux I__10498 (
            .O(N__49266),
            .I(N__49180));
    Span4Mux_h I__10497 (
            .O(N__49261),
            .I(N__49176));
    Span4Mux_h I__10496 (
            .O(N__49256),
            .I(N__49173));
    InMux I__10495 (
            .O(N__49255),
            .I(N__49166));
    InMux I__10494 (
            .O(N__49254),
            .I(N__49166));
    InMux I__10493 (
            .O(N__49253),
            .I(N__49166));
    Span4Mux_h I__10492 (
            .O(N__49250),
            .I(N__49161));
    LocalMux I__10491 (
            .O(N__49243),
            .I(N__49161));
    LocalMux I__10490 (
            .O(N__49236),
            .I(N__49156));
    Span4Mux_v I__10489 (
            .O(N__49231),
            .I(N__49156));
    LocalMux I__10488 (
            .O(N__49228),
            .I(N__49153));
    LocalMux I__10487 (
            .O(N__49223),
            .I(N__49150));
    Span4Mux_v I__10486 (
            .O(N__49212),
            .I(N__49145));
    Span4Mux_h I__10485 (
            .O(N__49207),
            .I(N__49145));
    Sp12to4 I__10484 (
            .O(N__49204),
            .I(N__49141));
    InMux I__10483 (
            .O(N__49203),
            .I(N__49136));
    InMux I__10482 (
            .O(N__49202),
            .I(N__49136));
    InMux I__10481 (
            .O(N__49201),
            .I(N__49133));
    Span4Mux_v I__10480 (
            .O(N__49198),
            .I(N__49130));
    LocalMux I__10479 (
            .O(N__49193),
            .I(N__49125));
    LocalMux I__10478 (
            .O(N__49190),
            .I(N__49125));
    LocalMux I__10477 (
            .O(N__49183),
            .I(N__49122));
    Span4Mux_h I__10476 (
            .O(N__49180),
            .I(N__49119));
    InMux I__10475 (
            .O(N__49179),
            .I(N__49116));
    Sp12to4 I__10474 (
            .O(N__49176),
            .I(N__49111));
    Sp12to4 I__10473 (
            .O(N__49173),
            .I(N__49111));
    LocalMux I__10472 (
            .O(N__49166),
            .I(N__49104));
    Span4Mux_v I__10471 (
            .O(N__49161),
            .I(N__49104));
    Span4Mux_v I__10470 (
            .O(N__49156),
            .I(N__49104));
    Span4Mux_h I__10469 (
            .O(N__49153),
            .I(N__49097));
    Span4Mux_v I__10468 (
            .O(N__49150),
            .I(N__49097));
    Span4Mux_h I__10467 (
            .O(N__49145),
            .I(N__49097));
    InMux I__10466 (
            .O(N__49144),
            .I(N__49094));
    Span12Mux_h I__10465 (
            .O(N__49141),
            .I(N__49087));
    LocalMux I__10464 (
            .O(N__49136),
            .I(N__49087));
    LocalMux I__10463 (
            .O(N__49133),
            .I(N__49087));
    Span4Mux_h I__10462 (
            .O(N__49130),
            .I(N__49084));
    Span12Mux_h I__10461 (
            .O(N__49125),
            .I(N__49081));
    Span4Mux_h I__10460 (
            .O(N__49122),
            .I(N__49076));
    Span4Mux_v I__10459 (
            .O(N__49119),
            .I(N__49076));
    LocalMux I__10458 (
            .O(N__49116),
            .I(N__49071));
    Span12Mux_v I__10457 (
            .O(N__49111),
            .I(N__49071));
    Span4Mux_h I__10456 (
            .O(N__49104),
            .I(N__49066));
    Span4Mux_v I__10455 (
            .O(N__49097),
            .I(N__49066));
    LocalMux I__10454 (
            .O(N__49094),
            .I(N__49061));
    Span12Mux_v I__10453 (
            .O(N__49087),
            .I(N__49061));
    Odrv4 I__10452 (
            .O(N__49084),
            .I(FRAME_MATCHER_state_31_N_2976_2));
    Odrv12 I__10451 (
            .O(N__49081),
            .I(FRAME_MATCHER_state_31_N_2976_2));
    Odrv4 I__10450 (
            .O(N__49076),
            .I(FRAME_MATCHER_state_31_N_2976_2));
    Odrv12 I__10449 (
            .O(N__49071),
            .I(FRAME_MATCHER_state_31_N_2976_2));
    Odrv4 I__10448 (
            .O(N__49066),
            .I(FRAME_MATCHER_state_31_N_2976_2));
    Odrv12 I__10447 (
            .O(N__49061),
            .I(FRAME_MATCHER_state_31_N_2976_2));
    InMux I__10446 (
            .O(N__49048),
            .I(N__49041));
    CascadeMux I__10445 (
            .O(N__49047),
            .I(N__49037));
    InMux I__10444 (
            .O(N__49046),
            .I(N__49030));
    InMux I__10443 (
            .O(N__49045),
            .I(N__49030));
    InMux I__10442 (
            .O(N__49044),
            .I(N__49030));
    LocalMux I__10441 (
            .O(N__49041),
            .I(N__49027));
    InMux I__10440 (
            .O(N__49040),
            .I(N__49014));
    InMux I__10439 (
            .O(N__49037),
            .I(N__49009));
    LocalMux I__10438 (
            .O(N__49030),
            .I(N__48994));
    Span4Mux_v I__10437 (
            .O(N__49027),
            .I(N__48994));
    InMux I__10436 (
            .O(N__49026),
            .I(N__48987));
    InMux I__10435 (
            .O(N__49025),
            .I(N__48987));
    InMux I__10434 (
            .O(N__49024),
            .I(N__48987));
    InMux I__10433 (
            .O(N__49023),
            .I(N__48982));
    InMux I__10432 (
            .O(N__49022),
            .I(N__48982));
    InMux I__10431 (
            .O(N__49021),
            .I(N__48971));
    InMux I__10430 (
            .O(N__49020),
            .I(N__48965));
    InMux I__10429 (
            .O(N__49019),
            .I(N__48962));
    InMux I__10428 (
            .O(N__49018),
            .I(N__48957));
    InMux I__10427 (
            .O(N__49017),
            .I(N__48957));
    LocalMux I__10426 (
            .O(N__49014),
            .I(N__48954));
    InMux I__10425 (
            .O(N__49013),
            .I(N__48950));
    InMux I__10424 (
            .O(N__49012),
            .I(N__48940));
    LocalMux I__10423 (
            .O(N__49009),
            .I(N__48935));
    InMux I__10422 (
            .O(N__49008),
            .I(N__48928));
    InMux I__10421 (
            .O(N__49007),
            .I(N__48928));
    InMux I__10420 (
            .O(N__49006),
            .I(N__48923));
    InMux I__10419 (
            .O(N__49005),
            .I(N__48923));
    InMux I__10418 (
            .O(N__49004),
            .I(N__48916));
    InMux I__10417 (
            .O(N__49003),
            .I(N__48916));
    InMux I__10416 (
            .O(N__49002),
            .I(N__48916));
    InMux I__10415 (
            .O(N__49001),
            .I(N__48909));
    InMux I__10414 (
            .O(N__49000),
            .I(N__48909));
    InMux I__10413 (
            .O(N__48999),
            .I(N__48909));
    Span4Mux_v I__10412 (
            .O(N__48994),
            .I(N__48904));
    LocalMux I__10411 (
            .O(N__48987),
            .I(N__48904));
    LocalMux I__10410 (
            .O(N__48982),
            .I(N__48901));
    CascadeMux I__10409 (
            .O(N__48981),
            .I(N__48898));
    InMux I__10408 (
            .O(N__48980),
            .I(N__48892));
    InMux I__10407 (
            .O(N__48979),
            .I(N__48877));
    InMux I__10406 (
            .O(N__48978),
            .I(N__48877));
    InMux I__10405 (
            .O(N__48977),
            .I(N__48877));
    InMux I__10404 (
            .O(N__48976),
            .I(N__48877));
    InMux I__10403 (
            .O(N__48975),
            .I(N__48872));
    InMux I__10402 (
            .O(N__48974),
            .I(N__48872));
    LocalMux I__10401 (
            .O(N__48971),
            .I(N__48869));
    InMux I__10400 (
            .O(N__48970),
            .I(N__48864));
    InMux I__10399 (
            .O(N__48969),
            .I(N__48864));
    InMux I__10398 (
            .O(N__48968),
            .I(N__48861));
    LocalMux I__10397 (
            .O(N__48965),
            .I(N__48858));
    LocalMux I__10396 (
            .O(N__48962),
            .I(N__48851));
    LocalMux I__10395 (
            .O(N__48957),
            .I(N__48851));
    Span4Mux_h I__10394 (
            .O(N__48954),
            .I(N__48851));
    CascadeMux I__10393 (
            .O(N__48953),
            .I(N__48848));
    LocalMux I__10392 (
            .O(N__48950),
            .I(N__48841));
    InMux I__10391 (
            .O(N__48949),
            .I(N__48834));
    InMux I__10390 (
            .O(N__48948),
            .I(N__48834));
    InMux I__10389 (
            .O(N__48947),
            .I(N__48834));
    InMux I__10388 (
            .O(N__48946),
            .I(N__48830));
    InMux I__10387 (
            .O(N__48945),
            .I(N__48827));
    InMux I__10386 (
            .O(N__48944),
            .I(N__48822));
    InMux I__10385 (
            .O(N__48943),
            .I(N__48822));
    LocalMux I__10384 (
            .O(N__48940),
            .I(N__48819));
    InMux I__10383 (
            .O(N__48939),
            .I(N__48814));
    InMux I__10382 (
            .O(N__48938),
            .I(N__48814));
    Span4Mux_v I__10381 (
            .O(N__48935),
            .I(N__48811));
    InMux I__10380 (
            .O(N__48934),
            .I(N__48806));
    InMux I__10379 (
            .O(N__48933),
            .I(N__48806));
    LocalMux I__10378 (
            .O(N__48928),
            .I(N__48801));
    LocalMux I__10377 (
            .O(N__48923),
            .I(N__48801));
    LocalMux I__10376 (
            .O(N__48916),
            .I(N__48792));
    LocalMux I__10375 (
            .O(N__48909),
            .I(N__48792));
    Span4Mux_h I__10374 (
            .O(N__48904),
            .I(N__48792));
    Span4Mux_h I__10373 (
            .O(N__48901),
            .I(N__48792));
    InMux I__10372 (
            .O(N__48898),
            .I(N__48789));
    InMux I__10371 (
            .O(N__48897),
            .I(N__48783));
    InMux I__10370 (
            .O(N__48896),
            .I(N__48783));
    InMux I__10369 (
            .O(N__48895),
            .I(N__48780));
    LocalMux I__10368 (
            .O(N__48892),
            .I(N__48777));
    InMux I__10367 (
            .O(N__48891),
            .I(N__48770));
    InMux I__10366 (
            .O(N__48890),
            .I(N__48770));
    InMux I__10365 (
            .O(N__48889),
            .I(N__48770));
    InMux I__10364 (
            .O(N__48888),
            .I(N__48763));
    InMux I__10363 (
            .O(N__48887),
            .I(N__48763));
    InMux I__10362 (
            .O(N__48886),
            .I(N__48763));
    LocalMux I__10361 (
            .O(N__48877),
            .I(N__48754));
    LocalMux I__10360 (
            .O(N__48872),
            .I(N__48754));
    Span4Mux_h I__10359 (
            .O(N__48869),
            .I(N__48754));
    LocalMux I__10358 (
            .O(N__48864),
            .I(N__48754));
    LocalMux I__10357 (
            .O(N__48861),
            .I(N__48747));
    Span4Mux_h I__10356 (
            .O(N__48858),
            .I(N__48747));
    Span4Mux_v I__10355 (
            .O(N__48851),
            .I(N__48747));
    InMux I__10354 (
            .O(N__48848),
            .I(N__48744));
    InMux I__10353 (
            .O(N__48847),
            .I(N__48728));
    InMux I__10352 (
            .O(N__48846),
            .I(N__48728));
    InMux I__10351 (
            .O(N__48845),
            .I(N__48723));
    InMux I__10350 (
            .O(N__48844),
            .I(N__48723));
    Span4Mux_h I__10349 (
            .O(N__48841),
            .I(N__48720));
    LocalMux I__10348 (
            .O(N__48834),
            .I(N__48717));
    InMux I__10347 (
            .O(N__48833),
            .I(N__48714));
    LocalMux I__10346 (
            .O(N__48830),
            .I(N__48709));
    LocalMux I__10345 (
            .O(N__48827),
            .I(N__48709));
    LocalMux I__10344 (
            .O(N__48822),
            .I(N__48706));
    Span4Mux_h I__10343 (
            .O(N__48819),
            .I(N__48703));
    LocalMux I__10342 (
            .O(N__48814),
            .I(N__48698));
    Span4Mux_v I__10341 (
            .O(N__48811),
            .I(N__48698));
    LocalMux I__10340 (
            .O(N__48806),
            .I(N__48690));
    Span4Mux_h I__10339 (
            .O(N__48801),
            .I(N__48690));
    Span4Mux_v I__10338 (
            .O(N__48792),
            .I(N__48690));
    LocalMux I__10337 (
            .O(N__48789),
            .I(N__48687));
    InMux I__10336 (
            .O(N__48788),
            .I(N__48684));
    LocalMux I__10335 (
            .O(N__48783),
            .I(N__48681));
    LocalMux I__10334 (
            .O(N__48780),
            .I(N__48676));
    Span4Mux_v I__10333 (
            .O(N__48777),
            .I(N__48676));
    LocalMux I__10332 (
            .O(N__48770),
            .I(N__48667));
    LocalMux I__10331 (
            .O(N__48763),
            .I(N__48667));
    Span4Mux_v I__10330 (
            .O(N__48754),
            .I(N__48667));
    Span4Mux_v I__10329 (
            .O(N__48747),
            .I(N__48667));
    LocalMux I__10328 (
            .O(N__48744),
            .I(N__48664));
    InMux I__10327 (
            .O(N__48743),
            .I(N__48659));
    InMux I__10326 (
            .O(N__48742),
            .I(N__48659));
    InMux I__10325 (
            .O(N__48741),
            .I(N__48656));
    InMux I__10324 (
            .O(N__48740),
            .I(N__48647));
    InMux I__10323 (
            .O(N__48739),
            .I(N__48647));
    InMux I__10322 (
            .O(N__48738),
            .I(N__48647));
    InMux I__10321 (
            .O(N__48737),
            .I(N__48647));
    InMux I__10320 (
            .O(N__48736),
            .I(N__48642));
    InMux I__10319 (
            .O(N__48735),
            .I(N__48642));
    InMux I__10318 (
            .O(N__48734),
            .I(N__48637));
    InMux I__10317 (
            .O(N__48733),
            .I(N__48637));
    LocalMux I__10316 (
            .O(N__48728),
            .I(N__48632));
    LocalMux I__10315 (
            .O(N__48723),
            .I(N__48632));
    Span4Mux_v I__10314 (
            .O(N__48720),
            .I(N__48629));
    Span12Mux_s11_v I__10313 (
            .O(N__48717),
            .I(N__48626));
    LocalMux I__10312 (
            .O(N__48714),
            .I(N__48615));
    Span4Mux_h I__10311 (
            .O(N__48709),
            .I(N__48615));
    Span4Mux_h I__10310 (
            .O(N__48706),
            .I(N__48615));
    Span4Mux_h I__10309 (
            .O(N__48703),
            .I(N__48615));
    Span4Mux_h I__10308 (
            .O(N__48698),
            .I(N__48615));
    InMux I__10307 (
            .O(N__48697),
            .I(N__48612));
    Span4Mux_h I__10306 (
            .O(N__48690),
            .I(N__48605));
    Span4Mux_h I__10305 (
            .O(N__48687),
            .I(N__48605));
    LocalMux I__10304 (
            .O(N__48684),
            .I(N__48605));
    Span4Mux_h I__10303 (
            .O(N__48681),
            .I(N__48596));
    Span4Mux_v I__10302 (
            .O(N__48676),
            .I(N__48596));
    Span4Mux_h I__10301 (
            .O(N__48667),
            .I(N__48596));
    Span4Mux_h I__10300 (
            .O(N__48664),
            .I(N__48596));
    LocalMux I__10299 (
            .O(N__48659),
            .I(n22661));
    LocalMux I__10298 (
            .O(N__48656),
            .I(n22661));
    LocalMux I__10297 (
            .O(N__48647),
            .I(n22661));
    LocalMux I__10296 (
            .O(N__48642),
            .I(n22661));
    LocalMux I__10295 (
            .O(N__48637),
            .I(n22661));
    Odrv12 I__10294 (
            .O(N__48632),
            .I(n22661));
    Odrv4 I__10293 (
            .O(N__48629),
            .I(n22661));
    Odrv12 I__10292 (
            .O(N__48626),
            .I(n22661));
    Odrv4 I__10291 (
            .O(N__48615),
            .I(n22661));
    LocalMux I__10290 (
            .O(N__48612),
            .I(n22661));
    Odrv4 I__10289 (
            .O(N__48605),
            .I(n22661));
    Odrv4 I__10288 (
            .O(N__48596),
            .I(n22661));
    CascadeMux I__10287 (
            .O(N__48571),
            .I(N__48567));
    CascadeMux I__10286 (
            .O(N__48570),
            .I(N__48563));
    InMux I__10285 (
            .O(N__48567),
            .I(N__48559));
    CascadeMux I__10284 (
            .O(N__48566),
            .I(N__48554));
    InMux I__10283 (
            .O(N__48563),
            .I(N__48548));
    InMux I__10282 (
            .O(N__48562),
            .I(N__48545));
    LocalMux I__10281 (
            .O(N__48559),
            .I(N__48542));
    InMux I__10280 (
            .O(N__48558),
            .I(N__48537));
    InMux I__10279 (
            .O(N__48557),
            .I(N__48537));
    InMux I__10278 (
            .O(N__48554),
            .I(N__48534));
    InMux I__10277 (
            .O(N__48553),
            .I(N__48530));
    InMux I__10276 (
            .O(N__48552),
            .I(N__48527));
    InMux I__10275 (
            .O(N__48551),
            .I(N__48524));
    LocalMux I__10274 (
            .O(N__48548),
            .I(N__48519));
    LocalMux I__10273 (
            .O(N__48545),
            .I(N__48519));
    Span4Mux_h I__10272 (
            .O(N__48542),
            .I(N__48516));
    LocalMux I__10271 (
            .O(N__48537),
            .I(N__48511));
    LocalMux I__10270 (
            .O(N__48534),
            .I(N__48511));
    InMux I__10269 (
            .O(N__48533),
            .I(N__48508));
    LocalMux I__10268 (
            .O(N__48530),
            .I(N__48503));
    LocalMux I__10267 (
            .O(N__48527),
            .I(N__48503));
    LocalMux I__10266 (
            .O(N__48524),
            .I(N__48498));
    Span4Mux_h I__10265 (
            .O(N__48519),
            .I(N__48498));
    Span4Mux_h I__10264 (
            .O(N__48516),
            .I(N__48493));
    Span4Mux_h I__10263 (
            .O(N__48511),
            .I(N__48493));
    LocalMux I__10262 (
            .O(N__48508),
            .I(encoder0_position_30));
    Odrv4 I__10261 (
            .O(N__48503),
            .I(encoder0_position_30));
    Odrv4 I__10260 (
            .O(N__48498),
            .I(encoder0_position_30));
    Odrv4 I__10259 (
            .O(N__48493),
            .I(encoder0_position_30));
    InMux I__10258 (
            .O(N__48484),
            .I(N__48481));
    LocalMux I__10257 (
            .O(N__48481),
            .I(N__48477));
    InMux I__10256 (
            .O(N__48480),
            .I(N__48474));
    Span4Mux_h I__10255 (
            .O(N__48477),
            .I(N__48471));
    LocalMux I__10254 (
            .O(N__48474),
            .I(data_out_frame_6_6));
    Odrv4 I__10253 (
            .O(N__48471),
            .I(data_out_frame_6_6));
    CascadeMux I__10252 (
            .O(N__48466),
            .I(N__48463));
    InMux I__10251 (
            .O(N__48463),
            .I(N__48460));
    LocalMux I__10250 (
            .O(N__48460),
            .I(N__48457));
    Span4Mux_v I__10249 (
            .O(N__48457),
            .I(N__48454));
    Odrv4 I__10248 (
            .O(N__48454),
            .I(\c0.n6_adj_4241 ));
    InMux I__10247 (
            .O(N__48451),
            .I(N__48445));
    InMux I__10246 (
            .O(N__48450),
            .I(N__48442));
    InMux I__10245 (
            .O(N__48449),
            .I(N__48437));
    InMux I__10244 (
            .O(N__48448),
            .I(N__48437));
    LocalMux I__10243 (
            .O(N__48445),
            .I(N__48434));
    LocalMux I__10242 (
            .O(N__48442),
            .I(N__48431));
    LocalMux I__10241 (
            .O(N__48437),
            .I(N__48428));
    Span4Mux_h I__10240 (
            .O(N__48434),
            .I(N__48425));
    Span4Mux_v I__10239 (
            .O(N__48431),
            .I(N__48420));
    Span4Mux_h I__10238 (
            .O(N__48428),
            .I(N__48420));
    Odrv4 I__10237 (
            .O(N__48425),
            .I(\c0.n13086 ));
    Odrv4 I__10236 (
            .O(N__48420),
            .I(\c0.n13086 ));
    CascadeMux I__10235 (
            .O(N__48415),
            .I(N__48411));
    InMux I__10234 (
            .O(N__48414),
            .I(N__48405));
    InMux I__10233 (
            .O(N__48411),
            .I(N__48405));
    CascadeMux I__10232 (
            .O(N__48410),
            .I(N__48402));
    LocalMux I__10231 (
            .O(N__48405),
            .I(N__48398));
    InMux I__10230 (
            .O(N__48402),
            .I(N__48393));
    InMux I__10229 (
            .O(N__48401),
            .I(N__48393));
    Odrv12 I__10228 (
            .O(N__48398),
            .I(\c0.data_in_frame_8_5 ));
    LocalMux I__10227 (
            .O(N__48393),
            .I(\c0.data_in_frame_8_5 ));
    CascadeMux I__10226 (
            .O(N__48388),
            .I(\c0.n22415_cascade_ ));
    CascadeMux I__10225 (
            .O(N__48385),
            .I(N__48380));
    InMux I__10224 (
            .O(N__48384),
            .I(N__48375));
    InMux I__10223 (
            .O(N__48383),
            .I(N__48375));
    InMux I__10222 (
            .O(N__48380),
            .I(N__48372));
    LocalMux I__10221 (
            .O(N__48375),
            .I(N__48369));
    LocalMux I__10220 (
            .O(N__48372),
            .I(\c0.data_in_frame_10_5 ));
    Odrv4 I__10219 (
            .O(N__48369),
            .I(\c0.data_in_frame_10_5 ));
    InMux I__10218 (
            .O(N__48364),
            .I(N__48361));
    LocalMux I__10217 (
            .O(N__48361),
            .I(N__48358));
    Odrv12 I__10216 (
            .O(N__48358),
            .I(\c0.n35 ));
    CascadeMux I__10215 (
            .O(N__48355),
            .I(\c0.n13771_cascade_ ));
    InMux I__10214 (
            .O(N__48352),
            .I(N__48346));
    InMux I__10213 (
            .O(N__48351),
            .I(N__48346));
    LocalMux I__10212 (
            .O(N__48346),
            .I(\c0.n22239 ));
    CascadeMux I__10211 (
            .O(N__48343),
            .I(\c0.n4_cascade_ ));
    InMux I__10210 (
            .O(N__48340),
            .I(N__48337));
    LocalMux I__10209 (
            .O(N__48337),
            .I(\c0.n37 ));
    InMux I__10208 (
            .O(N__48334),
            .I(N__48331));
    LocalMux I__10207 (
            .O(N__48331),
            .I(N__48328));
    Span4Mux_h I__10206 (
            .O(N__48328),
            .I(N__48325));
    Odrv4 I__10205 (
            .O(N__48325),
            .I(\c0.n6_adj_4220 ));
    CascadeMux I__10204 (
            .O(N__48322),
            .I(N__48318));
    CascadeMux I__10203 (
            .O(N__48321),
            .I(N__48314));
    InMux I__10202 (
            .O(N__48318),
            .I(N__48311));
    CascadeMux I__10201 (
            .O(N__48317),
            .I(N__48308));
    InMux I__10200 (
            .O(N__48314),
            .I(N__48305));
    LocalMux I__10199 (
            .O(N__48311),
            .I(N__48302));
    InMux I__10198 (
            .O(N__48308),
            .I(N__48299));
    LocalMux I__10197 (
            .O(N__48305),
            .I(\c0.data_in_frame_8_3 ));
    Odrv12 I__10196 (
            .O(N__48302),
            .I(\c0.data_in_frame_8_3 ));
    LocalMux I__10195 (
            .O(N__48299),
            .I(\c0.data_in_frame_8_3 ));
    InMux I__10194 (
            .O(N__48292),
            .I(N__48289));
    LocalMux I__10193 (
            .O(N__48289),
            .I(\c0.n13652 ));
    InMux I__10192 (
            .O(N__48286),
            .I(N__48283));
    LocalMux I__10191 (
            .O(N__48283),
            .I(\c0.n13771 ));
    InMux I__10190 (
            .O(N__48280),
            .I(N__48274));
    InMux I__10189 (
            .O(N__48279),
            .I(N__48274));
    LocalMux I__10188 (
            .O(N__48274),
            .I(\c0.data_in_frame_10_3 ));
    CascadeMux I__10187 (
            .O(N__48271),
            .I(N__48268));
    InMux I__10186 (
            .O(N__48268),
            .I(N__48265));
    LocalMux I__10185 (
            .O(N__48265),
            .I(\c0.n21964 ));
    InMux I__10184 (
            .O(N__48262),
            .I(N__48259));
    LocalMux I__10183 (
            .O(N__48259),
            .I(N__48256));
    Span4Mux_h I__10182 (
            .O(N__48256),
            .I(N__48252));
    InMux I__10181 (
            .O(N__48255),
            .I(N__48249));
    Odrv4 I__10180 (
            .O(N__48252),
            .I(\c0.n22280 ));
    LocalMux I__10179 (
            .O(N__48249),
            .I(\c0.n22280 ));
    CascadeMux I__10178 (
            .O(N__48244),
            .I(\c0.n21964_cascade_ ));
    InMux I__10177 (
            .O(N__48241),
            .I(N__48237));
    InMux I__10176 (
            .O(N__48240),
            .I(N__48234));
    LocalMux I__10175 (
            .O(N__48237),
            .I(N__48229));
    LocalMux I__10174 (
            .O(N__48234),
            .I(N__48226));
    InMux I__10173 (
            .O(N__48233),
            .I(N__48221));
    InMux I__10172 (
            .O(N__48232),
            .I(N__48221));
    Span4Mux_h I__10171 (
            .O(N__48229),
            .I(N__48216));
    Span4Mux_h I__10170 (
            .O(N__48226),
            .I(N__48216));
    LocalMux I__10169 (
            .O(N__48221),
            .I(N__48213));
    Odrv4 I__10168 (
            .O(N__48216),
            .I(\c0.n14113 ));
    Odrv4 I__10167 (
            .O(N__48213),
            .I(\c0.n14113 ));
    CascadeMux I__10166 (
            .O(N__48208),
            .I(N__48205));
    InMux I__10165 (
            .O(N__48205),
            .I(N__48201));
    CascadeMux I__10164 (
            .O(N__48204),
            .I(N__48198));
    LocalMux I__10163 (
            .O(N__48201),
            .I(N__48193));
    InMux I__10162 (
            .O(N__48198),
            .I(N__48190));
    InMux I__10161 (
            .O(N__48197),
            .I(N__48185));
    InMux I__10160 (
            .O(N__48196),
            .I(N__48185));
    Span4Mux_h I__10159 (
            .O(N__48193),
            .I(N__48182));
    LocalMux I__10158 (
            .O(N__48190),
            .I(N__48177));
    LocalMux I__10157 (
            .O(N__48185),
            .I(N__48177));
    Odrv4 I__10156 (
            .O(N__48182),
            .I(\c0.data_in_frame_2_5 ));
    Odrv4 I__10155 (
            .O(N__48177),
            .I(\c0.data_in_frame_2_5 ));
    CascadeMux I__10154 (
            .O(N__48172),
            .I(N__48165));
    CascadeMux I__10153 (
            .O(N__48171),
            .I(N__48162));
    CascadeMux I__10152 (
            .O(N__48170),
            .I(N__48159));
    CascadeMux I__10151 (
            .O(N__48169),
            .I(N__48155));
    CascadeMux I__10150 (
            .O(N__48168),
            .I(N__48150));
    InMux I__10149 (
            .O(N__48165),
            .I(N__48145));
    InMux I__10148 (
            .O(N__48162),
            .I(N__48145));
    InMux I__10147 (
            .O(N__48159),
            .I(N__48140));
    InMux I__10146 (
            .O(N__48158),
            .I(N__48140));
    InMux I__10145 (
            .O(N__48155),
            .I(N__48134));
    InMux I__10144 (
            .O(N__48154),
            .I(N__48134));
    CascadeMux I__10143 (
            .O(N__48153),
            .I(N__48131));
    InMux I__10142 (
            .O(N__48150),
            .I(N__48128));
    LocalMux I__10141 (
            .O(N__48145),
            .I(N__48125));
    LocalMux I__10140 (
            .O(N__48140),
            .I(N__48122));
    InMux I__10139 (
            .O(N__48139),
            .I(N__48119));
    LocalMux I__10138 (
            .O(N__48134),
            .I(N__48116));
    InMux I__10137 (
            .O(N__48131),
            .I(N__48113));
    LocalMux I__10136 (
            .O(N__48128),
            .I(N__48108));
    Span4Mux_v I__10135 (
            .O(N__48125),
            .I(N__48108));
    Span4Mux_h I__10134 (
            .O(N__48122),
            .I(N__48101));
    LocalMux I__10133 (
            .O(N__48119),
            .I(N__48101));
    Span4Mux_v I__10132 (
            .O(N__48116),
            .I(N__48101));
    LocalMux I__10131 (
            .O(N__48113),
            .I(\c0.data_in_frame_0_3 ));
    Odrv4 I__10130 (
            .O(N__48108),
            .I(\c0.data_in_frame_0_3 ));
    Odrv4 I__10129 (
            .O(N__48101),
            .I(\c0.data_in_frame_0_3 ));
    CascadeMux I__10128 (
            .O(N__48094),
            .I(N__48091));
    InMux I__10127 (
            .O(N__48091),
            .I(N__48081));
    InMux I__10126 (
            .O(N__48090),
            .I(N__48081));
    InMux I__10125 (
            .O(N__48089),
            .I(N__48081));
    InMux I__10124 (
            .O(N__48088),
            .I(N__48078));
    LocalMux I__10123 (
            .O(N__48081),
            .I(N__48075));
    LocalMux I__10122 (
            .O(N__48078),
            .I(N__48072));
    Span4Mux_v I__10121 (
            .O(N__48075),
            .I(N__48069));
    Span4Mux_v I__10120 (
            .O(N__48072),
            .I(N__48066));
    Span4Mux_h I__10119 (
            .O(N__48069),
            .I(N__48063));
    Odrv4 I__10118 (
            .O(N__48066),
            .I(\c0.n13398 ));
    Odrv4 I__10117 (
            .O(N__48063),
            .I(\c0.n13398 ));
    InMux I__10116 (
            .O(N__48058),
            .I(N__48055));
    LocalMux I__10115 (
            .O(N__48055),
            .I(N__48052));
    Span4Mux_v I__10114 (
            .O(N__48052),
            .I(N__48049));
    Span4Mux_h I__10113 (
            .O(N__48049),
            .I(N__48043));
    InMux I__10112 (
            .O(N__48048),
            .I(N__48040));
    CascadeMux I__10111 (
            .O(N__48047),
            .I(N__48037));
    InMux I__10110 (
            .O(N__48046),
            .I(N__48034));
    Span4Mux_v I__10109 (
            .O(N__48043),
            .I(N__48029));
    LocalMux I__10108 (
            .O(N__48040),
            .I(N__48029));
    InMux I__10107 (
            .O(N__48037),
            .I(N__48023));
    LocalMux I__10106 (
            .O(N__48034),
            .I(N__48018));
    Span4Mux_h I__10105 (
            .O(N__48029),
            .I(N__48018));
    InMux I__10104 (
            .O(N__48028),
            .I(N__48015));
    InMux I__10103 (
            .O(N__48027),
            .I(N__48010));
    InMux I__10102 (
            .O(N__48026),
            .I(N__48010));
    LocalMux I__10101 (
            .O(N__48023),
            .I(data_in_frame_1_3));
    Odrv4 I__10100 (
            .O(N__48018),
            .I(data_in_frame_1_3));
    LocalMux I__10099 (
            .O(N__48015),
            .I(data_in_frame_1_3));
    LocalMux I__10098 (
            .O(N__48010),
            .I(data_in_frame_1_3));
    InMux I__10097 (
            .O(N__48001),
            .I(N__47998));
    LocalMux I__10096 (
            .O(N__47998),
            .I(N__47994));
    InMux I__10095 (
            .O(N__47997),
            .I(N__47989));
    Span4Mux_h I__10094 (
            .O(N__47994),
            .I(N__47986));
    InMux I__10093 (
            .O(N__47993),
            .I(N__47983));
    InMux I__10092 (
            .O(N__47992),
            .I(N__47980));
    LocalMux I__10091 (
            .O(N__47989),
            .I(\c0.data_in_frame_3_5 ));
    Odrv4 I__10090 (
            .O(N__47986),
            .I(\c0.data_in_frame_3_5 ));
    LocalMux I__10089 (
            .O(N__47983),
            .I(\c0.data_in_frame_3_5 ));
    LocalMux I__10088 (
            .O(N__47980),
            .I(\c0.data_in_frame_3_5 ));
    CascadeMux I__10087 (
            .O(N__47971),
            .I(\c0.n13398_cascade_ ));
    InMux I__10086 (
            .O(N__47968),
            .I(N__47962));
    InMux I__10085 (
            .O(N__47967),
            .I(N__47962));
    LocalMux I__10084 (
            .O(N__47962),
            .I(N__47959));
    Odrv4 I__10083 (
            .O(N__47959),
            .I(\c0.n13852 ));
    InMux I__10082 (
            .O(N__47956),
            .I(N__47953));
    LocalMux I__10081 (
            .O(N__47953),
            .I(N__47950));
    Span4Mux_h I__10080 (
            .O(N__47950),
            .I(N__47946));
    InMux I__10079 (
            .O(N__47949),
            .I(N__47943));
    Odrv4 I__10078 (
            .O(N__47946),
            .I(\c0.n21794 ));
    LocalMux I__10077 (
            .O(N__47943),
            .I(\c0.n21794 ));
    InMux I__10076 (
            .O(N__47938),
            .I(N__47934));
    CascadeMux I__10075 (
            .O(N__47937),
            .I(N__47931));
    LocalMux I__10074 (
            .O(N__47934),
            .I(N__47927));
    InMux I__10073 (
            .O(N__47931),
            .I(N__47924));
    InMux I__10072 (
            .O(N__47930),
            .I(N__47921));
    Span4Mux_h I__10071 (
            .O(N__47927),
            .I(N__47918));
    LocalMux I__10070 (
            .O(N__47924),
            .I(\c0.data_in_frame_8_2 ));
    LocalMux I__10069 (
            .O(N__47921),
            .I(\c0.data_in_frame_8_2 ));
    Odrv4 I__10068 (
            .O(N__47918),
            .I(\c0.data_in_frame_8_2 ));
    CascadeMux I__10067 (
            .O(N__47911),
            .I(\c0.n21794_cascade_ ));
    InMux I__10066 (
            .O(N__47908),
            .I(N__47903));
    CascadeMux I__10065 (
            .O(N__47907),
            .I(N__47898));
    InMux I__10064 (
            .O(N__47906),
            .I(N__47895));
    LocalMux I__10063 (
            .O(N__47903),
            .I(N__47892));
    InMux I__10062 (
            .O(N__47902),
            .I(N__47889));
    InMux I__10061 (
            .O(N__47901),
            .I(N__47884));
    InMux I__10060 (
            .O(N__47898),
            .I(N__47884));
    LocalMux I__10059 (
            .O(N__47895),
            .I(N__47880));
    Span4Mux_v I__10058 (
            .O(N__47892),
            .I(N__47877));
    LocalMux I__10057 (
            .O(N__47889),
            .I(N__47874));
    LocalMux I__10056 (
            .O(N__47884),
            .I(N__47871));
    InMux I__10055 (
            .O(N__47883),
            .I(N__47868));
    Sp12to4 I__10054 (
            .O(N__47880),
            .I(N__47865));
    Span4Mux_v I__10053 (
            .O(N__47877),
            .I(N__47860));
    Span4Mux_v I__10052 (
            .O(N__47874),
            .I(N__47860));
    Span4Mux_h I__10051 (
            .O(N__47871),
            .I(N__47857));
    LocalMux I__10050 (
            .O(N__47868),
            .I(\c0.data_in_frame_5_7 ));
    Odrv12 I__10049 (
            .O(N__47865),
            .I(\c0.data_in_frame_5_7 ));
    Odrv4 I__10048 (
            .O(N__47860),
            .I(\c0.data_in_frame_5_7 ));
    Odrv4 I__10047 (
            .O(N__47857),
            .I(\c0.data_in_frame_5_7 ));
    CascadeMux I__10046 (
            .O(N__47848),
            .I(\c0.n6_adj_4257_cascade_ ));
    InMux I__10045 (
            .O(N__47845),
            .I(N__47841));
    InMux I__10044 (
            .O(N__47844),
            .I(N__47838));
    LocalMux I__10043 (
            .O(N__47841),
            .I(N__47835));
    LocalMux I__10042 (
            .O(N__47838),
            .I(N__47830));
    Span4Mux_h I__10041 (
            .O(N__47835),
            .I(N__47830));
    Odrv4 I__10040 (
            .O(N__47830),
            .I(\c0.n21825 ));
    InMux I__10039 (
            .O(N__47827),
            .I(N__47824));
    LocalMux I__10038 (
            .O(N__47824),
            .I(N__47820));
    InMux I__10037 (
            .O(N__47823),
            .I(N__47817));
    Span4Mux_h I__10036 (
            .O(N__47820),
            .I(N__47814));
    LocalMux I__10035 (
            .O(N__47817),
            .I(\c0.data_in_frame_9_5 ));
    Odrv4 I__10034 (
            .O(N__47814),
            .I(\c0.data_in_frame_9_5 ));
    CascadeMux I__10033 (
            .O(N__47809),
            .I(\c0.n8_adj_4254_cascade_ ));
    InMux I__10032 (
            .O(N__47806),
            .I(N__47803));
    LocalMux I__10031 (
            .O(N__47803),
            .I(N__47799));
    InMux I__10030 (
            .O(N__47802),
            .I(N__47796));
    Span4Mux_h I__10029 (
            .O(N__47799),
            .I(N__47793));
    LocalMux I__10028 (
            .O(N__47796),
            .I(\c0.n4_adj_4255 ));
    Odrv4 I__10027 (
            .O(N__47793),
            .I(\c0.n4_adj_4255 ));
    CascadeMux I__10026 (
            .O(N__47788),
            .I(N__47784));
    CascadeMux I__10025 (
            .O(N__47787),
            .I(N__47781));
    InMux I__10024 (
            .O(N__47784),
            .I(N__47778));
    InMux I__10023 (
            .O(N__47781),
            .I(N__47775));
    LocalMux I__10022 (
            .O(N__47778),
            .I(N__47772));
    LocalMux I__10021 (
            .O(N__47775),
            .I(\c0.data_in_frame_5_5 ));
    Odrv4 I__10020 (
            .O(N__47772),
            .I(\c0.data_in_frame_5_5 ));
    CascadeMux I__10019 (
            .O(N__47767),
            .I(N__47763));
    InMux I__10018 (
            .O(N__47766),
            .I(N__47759));
    InMux I__10017 (
            .O(N__47763),
            .I(N__47755));
    InMux I__10016 (
            .O(N__47762),
            .I(N__47752));
    LocalMux I__10015 (
            .O(N__47759),
            .I(N__47749));
    InMux I__10014 (
            .O(N__47758),
            .I(N__47746));
    LocalMux I__10013 (
            .O(N__47755),
            .I(\c0.data_in_frame_3_1 ));
    LocalMux I__10012 (
            .O(N__47752),
            .I(\c0.data_in_frame_3_1 ));
    Odrv4 I__10011 (
            .O(N__47749),
            .I(\c0.data_in_frame_3_1 ));
    LocalMux I__10010 (
            .O(N__47746),
            .I(\c0.data_in_frame_3_1 ));
    InMux I__10009 (
            .O(N__47737),
            .I(N__47733));
    CascadeMux I__10008 (
            .O(N__47736),
            .I(N__47730));
    LocalMux I__10007 (
            .O(N__47733),
            .I(N__47727));
    InMux I__10006 (
            .O(N__47730),
            .I(N__47722));
    Span4Mux_h I__10005 (
            .O(N__47727),
            .I(N__47719));
    InMux I__10004 (
            .O(N__47726),
            .I(N__47714));
    InMux I__10003 (
            .O(N__47725),
            .I(N__47714));
    LocalMux I__10002 (
            .O(N__47722),
            .I(\c0.data_in_frame_3_2 ));
    Odrv4 I__10001 (
            .O(N__47719),
            .I(\c0.data_in_frame_3_2 ));
    LocalMux I__10000 (
            .O(N__47714),
            .I(\c0.data_in_frame_3_2 ));
    InMux I__9999 (
            .O(N__47707),
            .I(N__47704));
    LocalMux I__9998 (
            .O(N__47704),
            .I(\c0.n6_adj_4395 ));
    InMux I__9997 (
            .O(N__47701),
            .I(N__47697));
    InMux I__9996 (
            .O(N__47700),
            .I(N__47694));
    LocalMux I__9995 (
            .O(N__47697),
            .I(N__47690));
    LocalMux I__9994 (
            .O(N__47694),
            .I(N__47685));
    CascadeMux I__9993 (
            .O(N__47693),
            .I(N__47681));
    Span4Mux_h I__9992 (
            .O(N__47690),
            .I(N__47678));
    CascadeMux I__9991 (
            .O(N__47689),
            .I(N__47675));
    CascadeMux I__9990 (
            .O(N__47688),
            .I(N__47672));
    Span4Mux_v I__9989 (
            .O(N__47685),
            .I(N__47669));
    InMux I__9988 (
            .O(N__47684),
            .I(N__47664));
    InMux I__9987 (
            .O(N__47681),
            .I(N__47664));
    Span4Mux_v I__9986 (
            .O(N__47678),
            .I(N__47661));
    InMux I__9985 (
            .O(N__47675),
            .I(N__47656));
    InMux I__9984 (
            .O(N__47672),
            .I(N__47656));
    Span4Mux_v I__9983 (
            .O(N__47669),
            .I(N__47651));
    LocalMux I__9982 (
            .O(N__47664),
            .I(N__47651));
    Odrv4 I__9981 (
            .O(N__47661),
            .I(data_in_frame_1_1));
    LocalMux I__9980 (
            .O(N__47656),
            .I(data_in_frame_1_1));
    Odrv4 I__9979 (
            .O(N__47651),
            .I(data_in_frame_1_1));
    InMux I__9978 (
            .O(N__47644),
            .I(N__47641));
    LocalMux I__9977 (
            .O(N__47641),
            .I(N__47637));
    InMux I__9976 (
            .O(N__47640),
            .I(N__47634));
    Span4Mux_v I__9975 (
            .O(N__47637),
            .I(N__47628));
    LocalMux I__9974 (
            .O(N__47634),
            .I(N__47625));
    InMux I__9973 (
            .O(N__47633),
            .I(N__47620));
    InMux I__9972 (
            .O(N__47632),
            .I(N__47617));
    InMux I__9971 (
            .O(N__47631),
            .I(N__47612));
    Span4Mux_v I__9970 (
            .O(N__47628),
            .I(N__47607));
    Span4Mux_h I__9969 (
            .O(N__47625),
            .I(N__47607));
    InMux I__9968 (
            .O(N__47624),
            .I(N__47604));
    InMux I__9967 (
            .O(N__47623),
            .I(N__47601));
    LocalMux I__9966 (
            .O(N__47620),
            .I(N__47596));
    LocalMux I__9965 (
            .O(N__47617),
            .I(N__47596));
    InMux I__9964 (
            .O(N__47616),
            .I(N__47591));
    InMux I__9963 (
            .O(N__47615),
            .I(N__47591));
    LocalMux I__9962 (
            .O(N__47612),
            .I(data_in_frame_1_5));
    Odrv4 I__9961 (
            .O(N__47607),
            .I(data_in_frame_1_5));
    LocalMux I__9960 (
            .O(N__47604),
            .I(data_in_frame_1_5));
    LocalMux I__9959 (
            .O(N__47601),
            .I(data_in_frame_1_5));
    Odrv4 I__9958 (
            .O(N__47596),
            .I(data_in_frame_1_5));
    LocalMux I__9957 (
            .O(N__47591),
            .I(data_in_frame_1_5));
    InMux I__9956 (
            .O(N__47578),
            .I(N__47575));
    LocalMux I__9955 (
            .O(N__47575),
            .I(N__47572));
    Span4Mux_h I__9954 (
            .O(N__47572),
            .I(N__47569));
    Odrv4 I__9953 (
            .O(N__47569),
            .I(\c0.n21986 ));
    CascadeMux I__9952 (
            .O(N__47566),
            .I(\c0.n13848_cascade_ ));
    InMux I__9951 (
            .O(N__47563),
            .I(N__47560));
    LocalMux I__9950 (
            .O(N__47560),
            .I(N__47557));
    Span4Mux_h I__9949 (
            .O(N__47557),
            .I(N__47554));
    Span4Mux_v I__9948 (
            .O(N__47554),
            .I(N__47551));
    Odrv4 I__9947 (
            .O(N__47551),
            .I(\c0.n13_adj_4405 ));
    InMux I__9946 (
            .O(N__47548),
            .I(N__47544));
    CascadeMux I__9945 (
            .O(N__47547),
            .I(N__47541));
    LocalMux I__9944 (
            .O(N__47544),
            .I(N__47536));
    InMux I__9943 (
            .O(N__47541),
            .I(N__47529));
    InMux I__9942 (
            .O(N__47540),
            .I(N__47529));
    InMux I__9941 (
            .O(N__47539),
            .I(N__47529));
    Odrv4 I__9940 (
            .O(N__47536),
            .I(\c0.data_in_frame_2_7 ));
    LocalMux I__9939 (
            .O(N__47529),
            .I(\c0.data_in_frame_2_7 ));
    CascadeMux I__9938 (
            .O(N__47524),
            .I(N__47519));
    CascadeMux I__9937 (
            .O(N__47523),
            .I(N__47516));
    CascadeMux I__9936 (
            .O(N__47522),
            .I(N__47513));
    InMux I__9935 (
            .O(N__47519),
            .I(N__47510));
    InMux I__9934 (
            .O(N__47516),
            .I(N__47505));
    InMux I__9933 (
            .O(N__47513),
            .I(N__47502));
    LocalMux I__9932 (
            .O(N__47510),
            .I(N__47497));
    InMux I__9931 (
            .O(N__47509),
            .I(N__47494));
    CascadeMux I__9930 (
            .O(N__47508),
            .I(N__47490));
    LocalMux I__9929 (
            .O(N__47505),
            .I(N__47487));
    LocalMux I__9928 (
            .O(N__47502),
            .I(N__47484));
    InMux I__9927 (
            .O(N__47501),
            .I(N__47479));
    InMux I__9926 (
            .O(N__47500),
            .I(N__47479));
    Span4Mux_h I__9925 (
            .O(N__47497),
            .I(N__47476));
    LocalMux I__9924 (
            .O(N__47494),
            .I(N__47473));
    InMux I__9923 (
            .O(N__47493),
            .I(N__47468));
    InMux I__9922 (
            .O(N__47490),
            .I(N__47468));
    Odrv4 I__9921 (
            .O(N__47487),
            .I(\c0.data_in_frame_0_7 ));
    Odrv4 I__9920 (
            .O(N__47484),
            .I(\c0.data_in_frame_0_7 ));
    LocalMux I__9919 (
            .O(N__47479),
            .I(\c0.data_in_frame_0_7 ));
    Odrv4 I__9918 (
            .O(N__47476),
            .I(\c0.data_in_frame_0_7 ));
    Odrv4 I__9917 (
            .O(N__47473),
            .I(\c0.data_in_frame_0_7 ));
    LocalMux I__9916 (
            .O(N__47468),
            .I(\c0.data_in_frame_0_7 ));
    InMux I__9915 (
            .O(N__47455),
            .I(N__47451));
    InMux I__9914 (
            .O(N__47454),
            .I(N__47447));
    LocalMux I__9913 (
            .O(N__47451),
            .I(N__47443));
    InMux I__9912 (
            .O(N__47450),
            .I(N__47440));
    LocalMux I__9911 (
            .O(N__47447),
            .I(N__47437));
    InMux I__9910 (
            .O(N__47446),
            .I(N__47434));
    Span4Mux_v I__9909 (
            .O(N__47443),
            .I(N__47431));
    LocalMux I__9908 (
            .O(N__47440),
            .I(\c0.data_in_frame_8_4 ));
    Odrv4 I__9907 (
            .O(N__47437),
            .I(\c0.data_in_frame_8_4 ));
    LocalMux I__9906 (
            .O(N__47434),
            .I(\c0.data_in_frame_8_4 ));
    Odrv4 I__9905 (
            .O(N__47431),
            .I(\c0.data_in_frame_8_4 ));
    CascadeMux I__9904 (
            .O(N__47422),
            .I(\c0.n21861_cascade_ ));
    InMux I__9903 (
            .O(N__47419),
            .I(N__47416));
    LocalMux I__9902 (
            .O(N__47416),
            .I(\c0.n6_adj_4258 ));
    SRMux I__9901 (
            .O(N__47413),
            .I(N__47410));
    LocalMux I__9900 (
            .O(N__47410),
            .I(N__47407));
    Span4Mux_s2_v I__9899 (
            .O(N__47407),
            .I(N__47404));
    Odrv4 I__9898 (
            .O(N__47404),
            .I(\c0.n3_adj_4474 ));
    CascadeMux I__9897 (
            .O(N__47401),
            .I(N__47398));
    InMux I__9896 (
            .O(N__47398),
            .I(N__47395));
    LocalMux I__9895 (
            .O(N__47395),
            .I(N__47392));
    Span4Mux_v I__9894 (
            .O(N__47392),
            .I(N__47388));
    CascadeMux I__9893 (
            .O(N__47391),
            .I(N__47385));
    Span4Mux_v I__9892 (
            .O(N__47388),
            .I(N__47381));
    InMux I__9891 (
            .O(N__47385),
            .I(N__47377));
    InMux I__9890 (
            .O(N__47384),
            .I(N__47374));
    Span4Mux_h I__9889 (
            .O(N__47381),
            .I(N__47371));
    InMux I__9888 (
            .O(N__47380),
            .I(N__47368));
    LocalMux I__9887 (
            .O(N__47377),
            .I(\c0.FRAME_MATCHER_i_5 ));
    LocalMux I__9886 (
            .O(N__47374),
            .I(\c0.FRAME_MATCHER_i_5 ));
    Odrv4 I__9885 (
            .O(N__47371),
            .I(\c0.FRAME_MATCHER_i_5 ));
    LocalMux I__9884 (
            .O(N__47368),
            .I(\c0.FRAME_MATCHER_i_5 ));
    CascadeMux I__9883 (
            .O(N__47359),
            .I(N__47356));
    InMux I__9882 (
            .O(N__47356),
            .I(N__47352));
    InMux I__9881 (
            .O(N__47355),
            .I(N__47349));
    LocalMux I__9880 (
            .O(N__47352),
            .I(N__47342));
    LocalMux I__9879 (
            .O(N__47349),
            .I(N__47342));
    InMux I__9878 (
            .O(N__47348),
            .I(N__47339));
    InMux I__9877 (
            .O(N__47347),
            .I(N__47336));
    Span4Mux_v I__9876 (
            .O(N__47342),
            .I(N__47333));
    LocalMux I__9875 (
            .O(N__47339),
            .I(N__47326));
    LocalMux I__9874 (
            .O(N__47336),
            .I(N__47326));
    Span4Mux_v I__9873 (
            .O(N__47333),
            .I(N__47326));
    Odrv4 I__9872 (
            .O(N__47326),
            .I(\c0.FRAME_MATCHER_i_6 ));
    InMux I__9871 (
            .O(N__47323),
            .I(N__47317));
    CascadeMux I__9870 (
            .O(N__47322),
            .I(N__47314));
    CascadeMux I__9869 (
            .O(N__47321),
            .I(N__47311));
    InMux I__9868 (
            .O(N__47320),
            .I(N__47308));
    LocalMux I__9867 (
            .O(N__47317),
            .I(N__47305));
    InMux I__9866 (
            .O(N__47314),
            .I(N__47300));
    InMux I__9865 (
            .O(N__47311),
            .I(N__47300));
    LocalMux I__9864 (
            .O(N__47308),
            .I(N__47297));
    Span4Mux_h I__9863 (
            .O(N__47305),
            .I(N__47294));
    LocalMux I__9862 (
            .O(N__47300),
            .I(N__47291));
    Span4Mux_h I__9861 (
            .O(N__47297),
            .I(N__47288));
    Span4Mux_h I__9860 (
            .O(N__47294),
            .I(N__47283));
    Span4Mux_h I__9859 (
            .O(N__47291),
            .I(N__47283));
    Span4Mux_v I__9858 (
            .O(N__47288),
            .I(N__47280));
    Span4Mux_v I__9857 (
            .O(N__47283),
            .I(N__47277));
    Span4Mux_v I__9856 (
            .O(N__47280),
            .I(N__47274));
    Span4Mux_v I__9855 (
            .O(N__47277),
            .I(N__47271));
    Odrv4 I__9854 (
            .O(N__47274),
            .I(\c0.n11_adj_4326 ));
    Odrv4 I__9853 (
            .O(N__47271),
            .I(\c0.n11_adj_4326 ));
    InMux I__9852 (
            .O(N__47266),
            .I(N__47263));
    LocalMux I__9851 (
            .O(N__47263),
            .I(N__47260));
    Span4Mux_h I__9850 (
            .O(N__47260),
            .I(N__47257));
    Odrv4 I__9849 (
            .O(N__47257),
            .I(\c0.n10_adj_4399 ));
    InMux I__9848 (
            .O(N__47254),
            .I(N__47250));
    InMux I__9847 (
            .O(N__47253),
            .I(N__47247));
    LocalMux I__9846 (
            .O(N__47250),
            .I(N__47243));
    LocalMux I__9845 (
            .O(N__47247),
            .I(N__47240));
    InMux I__9844 (
            .O(N__47246),
            .I(N__47236));
    Span4Mux_h I__9843 (
            .O(N__47243),
            .I(N__47233));
    Span4Mux_h I__9842 (
            .O(N__47240),
            .I(N__47230));
    InMux I__9841 (
            .O(N__47239),
            .I(N__47227));
    LocalMux I__9840 (
            .O(N__47236),
            .I(\c0.n13033 ));
    Odrv4 I__9839 (
            .O(N__47233),
            .I(\c0.n13033 ));
    Odrv4 I__9838 (
            .O(N__47230),
            .I(\c0.n13033 ));
    LocalMux I__9837 (
            .O(N__47227),
            .I(\c0.n13033 ));
    IoInMux I__9836 (
            .O(N__47218),
            .I(N__47203));
    CascadeMux I__9835 (
            .O(N__47217),
            .I(N__47199));
    CascadeMux I__9834 (
            .O(N__47216),
            .I(N__47195));
    CascadeMux I__9833 (
            .O(N__47215),
            .I(N__47191));
    CascadeMux I__9832 (
            .O(N__47214),
            .I(N__47186));
    CascadeMux I__9831 (
            .O(N__47213),
            .I(N__47182));
    CascadeMux I__9830 (
            .O(N__47212),
            .I(N__47178));
    CascadeMux I__9829 (
            .O(N__47211),
            .I(N__47173));
    CascadeMux I__9828 (
            .O(N__47210),
            .I(N__47169));
    CascadeMux I__9827 (
            .O(N__47209),
            .I(N__47165));
    CascadeMux I__9826 (
            .O(N__47208),
            .I(N__47160));
    CascadeMux I__9825 (
            .O(N__47207),
            .I(N__47156));
    CascadeMux I__9824 (
            .O(N__47206),
            .I(N__47152));
    LocalMux I__9823 (
            .O(N__47203),
            .I(N__47136));
    InMux I__9822 (
            .O(N__47202),
            .I(N__47121));
    InMux I__9821 (
            .O(N__47199),
            .I(N__47121));
    InMux I__9820 (
            .O(N__47198),
            .I(N__47121));
    InMux I__9819 (
            .O(N__47195),
            .I(N__47121));
    InMux I__9818 (
            .O(N__47194),
            .I(N__47121));
    InMux I__9817 (
            .O(N__47191),
            .I(N__47121));
    InMux I__9816 (
            .O(N__47190),
            .I(N__47121));
    InMux I__9815 (
            .O(N__47189),
            .I(N__47106));
    InMux I__9814 (
            .O(N__47186),
            .I(N__47106));
    InMux I__9813 (
            .O(N__47185),
            .I(N__47106));
    InMux I__9812 (
            .O(N__47182),
            .I(N__47106));
    InMux I__9811 (
            .O(N__47181),
            .I(N__47106));
    InMux I__9810 (
            .O(N__47178),
            .I(N__47106));
    InMux I__9809 (
            .O(N__47177),
            .I(N__47106));
    InMux I__9808 (
            .O(N__47176),
            .I(N__47091));
    InMux I__9807 (
            .O(N__47173),
            .I(N__47091));
    InMux I__9806 (
            .O(N__47172),
            .I(N__47091));
    InMux I__9805 (
            .O(N__47169),
            .I(N__47091));
    InMux I__9804 (
            .O(N__47168),
            .I(N__47091));
    InMux I__9803 (
            .O(N__47165),
            .I(N__47091));
    InMux I__9802 (
            .O(N__47164),
            .I(N__47091));
    InMux I__9801 (
            .O(N__47163),
            .I(N__47076));
    InMux I__9800 (
            .O(N__47160),
            .I(N__47076));
    InMux I__9799 (
            .O(N__47159),
            .I(N__47076));
    InMux I__9798 (
            .O(N__47156),
            .I(N__47076));
    InMux I__9797 (
            .O(N__47155),
            .I(N__47076));
    InMux I__9796 (
            .O(N__47152),
            .I(N__47076));
    InMux I__9795 (
            .O(N__47151),
            .I(N__47076));
    CascadeMux I__9794 (
            .O(N__47150),
            .I(N__47072));
    CascadeMux I__9793 (
            .O(N__47149),
            .I(N__47068));
    CascadeMux I__9792 (
            .O(N__47148),
            .I(N__47064));
    CascadeMux I__9791 (
            .O(N__47147),
            .I(N__47059));
    CascadeMux I__9790 (
            .O(N__47146),
            .I(N__47055));
    CascadeMux I__9789 (
            .O(N__47145),
            .I(N__47051));
    CascadeMux I__9788 (
            .O(N__47144),
            .I(N__47046));
    CascadeMux I__9787 (
            .O(N__47143),
            .I(N__47042));
    CascadeMux I__9786 (
            .O(N__47142),
            .I(N__47038));
    CascadeMux I__9785 (
            .O(N__47141),
            .I(N__47033));
    CascadeMux I__9784 (
            .O(N__47140),
            .I(N__47029));
    CascadeMux I__9783 (
            .O(N__47139),
            .I(N__47025));
    IoSpan4Mux I__9782 (
            .O(N__47136),
            .I(N__47003));
    LocalMux I__9781 (
            .O(N__47121),
            .I(N__47003));
    LocalMux I__9780 (
            .O(N__47106),
            .I(N__47003));
    LocalMux I__9779 (
            .O(N__47091),
            .I(N__47003));
    LocalMux I__9778 (
            .O(N__47076),
            .I(N__47000));
    InMux I__9777 (
            .O(N__47075),
            .I(N__46985));
    InMux I__9776 (
            .O(N__47072),
            .I(N__46985));
    InMux I__9775 (
            .O(N__47071),
            .I(N__46985));
    InMux I__9774 (
            .O(N__47068),
            .I(N__46985));
    InMux I__9773 (
            .O(N__47067),
            .I(N__46985));
    InMux I__9772 (
            .O(N__47064),
            .I(N__46985));
    InMux I__9771 (
            .O(N__47063),
            .I(N__46985));
    InMux I__9770 (
            .O(N__47062),
            .I(N__46970));
    InMux I__9769 (
            .O(N__47059),
            .I(N__46970));
    InMux I__9768 (
            .O(N__47058),
            .I(N__46970));
    InMux I__9767 (
            .O(N__47055),
            .I(N__46970));
    InMux I__9766 (
            .O(N__47054),
            .I(N__46970));
    InMux I__9765 (
            .O(N__47051),
            .I(N__46970));
    InMux I__9764 (
            .O(N__47050),
            .I(N__46970));
    InMux I__9763 (
            .O(N__47049),
            .I(N__46955));
    InMux I__9762 (
            .O(N__47046),
            .I(N__46955));
    InMux I__9761 (
            .O(N__47045),
            .I(N__46955));
    InMux I__9760 (
            .O(N__47042),
            .I(N__46955));
    InMux I__9759 (
            .O(N__47041),
            .I(N__46955));
    InMux I__9758 (
            .O(N__47038),
            .I(N__46955));
    InMux I__9757 (
            .O(N__47037),
            .I(N__46955));
    InMux I__9756 (
            .O(N__47036),
            .I(N__46940));
    InMux I__9755 (
            .O(N__47033),
            .I(N__46940));
    InMux I__9754 (
            .O(N__47032),
            .I(N__46940));
    InMux I__9753 (
            .O(N__47029),
            .I(N__46940));
    InMux I__9752 (
            .O(N__47028),
            .I(N__46940));
    InMux I__9751 (
            .O(N__47025),
            .I(N__46940));
    InMux I__9750 (
            .O(N__47024),
            .I(N__46940));
    CascadeMux I__9749 (
            .O(N__47023),
            .I(N__46936));
    CascadeMux I__9748 (
            .O(N__47022),
            .I(N__46932));
    CascadeMux I__9747 (
            .O(N__47021),
            .I(N__46928));
    CascadeMux I__9746 (
            .O(N__47020),
            .I(N__46923));
    CascadeMux I__9745 (
            .O(N__47019),
            .I(N__46919));
    CascadeMux I__9744 (
            .O(N__47018),
            .I(N__46915));
    CascadeMux I__9743 (
            .O(N__47017),
            .I(N__46910));
    CascadeMux I__9742 (
            .O(N__47016),
            .I(N__46906));
    CascadeMux I__9741 (
            .O(N__47015),
            .I(N__46902));
    CascadeMux I__9740 (
            .O(N__47014),
            .I(N__46897));
    CascadeMux I__9739 (
            .O(N__47013),
            .I(N__46893));
    CascadeMux I__9738 (
            .O(N__47012),
            .I(N__46889));
    Span4Mux_s3_v I__9737 (
            .O(N__47003),
            .I(N__46865));
    Span4Mux_h I__9736 (
            .O(N__47000),
            .I(N__46865));
    LocalMux I__9735 (
            .O(N__46985),
            .I(N__46865));
    LocalMux I__9734 (
            .O(N__46970),
            .I(N__46865));
    LocalMux I__9733 (
            .O(N__46955),
            .I(N__46865));
    LocalMux I__9732 (
            .O(N__46940),
            .I(N__46862));
    InMux I__9731 (
            .O(N__46939),
            .I(N__46847));
    InMux I__9730 (
            .O(N__46936),
            .I(N__46847));
    InMux I__9729 (
            .O(N__46935),
            .I(N__46847));
    InMux I__9728 (
            .O(N__46932),
            .I(N__46847));
    InMux I__9727 (
            .O(N__46931),
            .I(N__46847));
    InMux I__9726 (
            .O(N__46928),
            .I(N__46847));
    InMux I__9725 (
            .O(N__46927),
            .I(N__46847));
    InMux I__9724 (
            .O(N__46926),
            .I(N__46832));
    InMux I__9723 (
            .O(N__46923),
            .I(N__46832));
    InMux I__9722 (
            .O(N__46922),
            .I(N__46832));
    InMux I__9721 (
            .O(N__46919),
            .I(N__46832));
    InMux I__9720 (
            .O(N__46918),
            .I(N__46832));
    InMux I__9719 (
            .O(N__46915),
            .I(N__46832));
    InMux I__9718 (
            .O(N__46914),
            .I(N__46832));
    InMux I__9717 (
            .O(N__46913),
            .I(N__46817));
    InMux I__9716 (
            .O(N__46910),
            .I(N__46817));
    InMux I__9715 (
            .O(N__46909),
            .I(N__46817));
    InMux I__9714 (
            .O(N__46906),
            .I(N__46817));
    InMux I__9713 (
            .O(N__46905),
            .I(N__46817));
    InMux I__9712 (
            .O(N__46902),
            .I(N__46817));
    InMux I__9711 (
            .O(N__46901),
            .I(N__46817));
    InMux I__9710 (
            .O(N__46900),
            .I(N__46802));
    InMux I__9709 (
            .O(N__46897),
            .I(N__46802));
    InMux I__9708 (
            .O(N__46896),
            .I(N__46802));
    InMux I__9707 (
            .O(N__46893),
            .I(N__46802));
    InMux I__9706 (
            .O(N__46892),
            .I(N__46802));
    InMux I__9705 (
            .O(N__46889),
            .I(N__46802));
    InMux I__9704 (
            .O(N__46888),
            .I(N__46802));
    CascadeMux I__9703 (
            .O(N__46887),
            .I(N__46798));
    CascadeMux I__9702 (
            .O(N__46886),
            .I(N__46794));
    CascadeMux I__9701 (
            .O(N__46885),
            .I(N__46790));
    CascadeMux I__9700 (
            .O(N__46884),
            .I(N__46785));
    CascadeMux I__9699 (
            .O(N__46883),
            .I(N__46781));
    CascadeMux I__9698 (
            .O(N__46882),
            .I(N__46777));
    CascadeMux I__9697 (
            .O(N__46881),
            .I(N__46772));
    CascadeMux I__9696 (
            .O(N__46880),
            .I(N__46768));
    CascadeMux I__9695 (
            .O(N__46879),
            .I(N__46764));
    CascadeMux I__9694 (
            .O(N__46878),
            .I(N__46759));
    CascadeMux I__9693 (
            .O(N__46877),
            .I(N__46755));
    CascadeMux I__9692 (
            .O(N__46876),
            .I(N__46751));
    Span4Mux_v I__9691 (
            .O(N__46865),
            .I(N__46730));
    Span4Mux_h I__9690 (
            .O(N__46862),
            .I(N__46730));
    LocalMux I__9689 (
            .O(N__46847),
            .I(N__46730));
    LocalMux I__9688 (
            .O(N__46832),
            .I(N__46730));
    LocalMux I__9687 (
            .O(N__46817),
            .I(N__46730));
    LocalMux I__9686 (
            .O(N__46802),
            .I(N__46727));
    InMux I__9685 (
            .O(N__46801),
            .I(N__46712));
    InMux I__9684 (
            .O(N__46798),
            .I(N__46712));
    InMux I__9683 (
            .O(N__46797),
            .I(N__46712));
    InMux I__9682 (
            .O(N__46794),
            .I(N__46712));
    InMux I__9681 (
            .O(N__46793),
            .I(N__46712));
    InMux I__9680 (
            .O(N__46790),
            .I(N__46712));
    InMux I__9679 (
            .O(N__46789),
            .I(N__46712));
    InMux I__9678 (
            .O(N__46788),
            .I(N__46697));
    InMux I__9677 (
            .O(N__46785),
            .I(N__46697));
    InMux I__9676 (
            .O(N__46784),
            .I(N__46697));
    InMux I__9675 (
            .O(N__46781),
            .I(N__46697));
    InMux I__9674 (
            .O(N__46780),
            .I(N__46697));
    InMux I__9673 (
            .O(N__46777),
            .I(N__46697));
    InMux I__9672 (
            .O(N__46776),
            .I(N__46697));
    InMux I__9671 (
            .O(N__46775),
            .I(N__46682));
    InMux I__9670 (
            .O(N__46772),
            .I(N__46682));
    InMux I__9669 (
            .O(N__46771),
            .I(N__46682));
    InMux I__9668 (
            .O(N__46768),
            .I(N__46682));
    InMux I__9667 (
            .O(N__46767),
            .I(N__46682));
    InMux I__9666 (
            .O(N__46764),
            .I(N__46682));
    InMux I__9665 (
            .O(N__46763),
            .I(N__46682));
    InMux I__9664 (
            .O(N__46762),
            .I(N__46667));
    InMux I__9663 (
            .O(N__46759),
            .I(N__46667));
    InMux I__9662 (
            .O(N__46758),
            .I(N__46667));
    InMux I__9661 (
            .O(N__46755),
            .I(N__46667));
    InMux I__9660 (
            .O(N__46754),
            .I(N__46667));
    InMux I__9659 (
            .O(N__46751),
            .I(N__46667));
    InMux I__9658 (
            .O(N__46750),
            .I(N__46667));
    CascadeMux I__9657 (
            .O(N__46749),
            .I(N__46663));
    CascadeMux I__9656 (
            .O(N__46748),
            .I(N__46659));
    CascadeMux I__9655 (
            .O(N__46747),
            .I(N__46655));
    CascadeMux I__9654 (
            .O(N__46746),
            .I(N__46650));
    CascadeMux I__9653 (
            .O(N__46745),
            .I(N__46646));
    CascadeMux I__9652 (
            .O(N__46744),
            .I(N__46642));
    CascadeMux I__9651 (
            .O(N__46743),
            .I(N__46637));
    CascadeMux I__9650 (
            .O(N__46742),
            .I(N__46633));
    CascadeMux I__9649 (
            .O(N__46741),
            .I(N__46629));
    Span4Mux_v I__9648 (
            .O(N__46730),
            .I(N__46603));
    Span4Mux_h I__9647 (
            .O(N__46727),
            .I(N__46603));
    LocalMux I__9646 (
            .O(N__46712),
            .I(N__46603));
    LocalMux I__9645 (
            .O(N__46697),
            .I(N__46603));
    LocalMux I__9644 (
            .O(N__46682),
            .I(N__46603));
    LocalMux I__9643 (
            .O(N__46667),
            .I(N__46603));
    InMux I__9642 (
            .O(N__46666),
            .I(N__46588));
    InMux I__9641 (
            .O(N__46663),
            .I(N__46588));
    InMux I__9640 (
            .O(N__46662),
            .I(N__46588));
    InMux I__9639 (
            .O(N__46659),
            .I(N__46588));
    InMux I__9638 (
            .O(N__46658),
            .I(N__46588));
    InMux I__9637 (
            .O(N__46655),
            .I(N__46588));
    InMux I__9636 (
            .O(N__46654),
            .I(N__46588));
    InMux I__9635 (
            .O(N__46653),
            .I(N__46573));
    InMux I__9634 (
            .O(N__46650),
            .I(N__46573));
    InMux I__9633 (
            .O(N__46649),
            .I(N__46573));
    InMux I__9632 (
            .O(N__46646),
            .I(N__46573));
    InMux I__9631 (
            .O(N__46645),
            .I(N__46573));
    InMux I__9630 (
            .O(N__46642),
            .I(N__46573));
    InMux I__9629 (
            .O(N__46641),
            .I(N__46573));
    InMux I__9628 (
            .O(N__46640),
            .I(N__46558));
    InMux I__9627 (
            .O(N__46637),
            .I(N__46558));
    InMux I__9626 (
            .O(N__46636),
            .I(N__46558));
    InMux I__9625 (
            .O(N__46633),
            .I(N__46558));
    InMux I__9624 (
            .O(N__46632),
            .I(N__46558));
    InMux I__9623 (
            .O(N__46629),
            .I(N__46558));
    InMux I__9622 (
            .O(N__46628),
            .I(N__46558));
    CascadeMux I__9621 (
            .O(N__46627),
            .I(N__46554));
    CascadeMux I__9620 (
            .O(N__46626),
            .I(N__46550));
    CascadeMux I__9619 (
            .O(N__46625),
            .I(N__46546));
    CascadeMux I__9618 (
            .O(N__46624),
            .I(N__46541));
    CascadeMux I__9617 (
            .O(N__46623),
            .I(N__46537));
    CascadeMux I__9616 (
            .O(N__46622),
            .I(N__46533));
    CascadeMux I__9615 (
            .O(N__46621),
            .I(N__46504));
    CascadeMux I__9614 (
            .O(N__46620),
            .I(N__46500));
    CascadeMux I__9613 (
            .O(N__46619),
            .I(N__46496));
    CascadeMux I__9612 (
            .O(N__46618),
            .I(N__46488));
    CascadeMux I__9611 (
            .O(N__46617),
            .I(N__46484));
    CascadeMux I__9610 (
            .O(N__46616),
            .I(N__46480));
    Span4Mux_v I__9609 (
            .O(N__46603),
            .I(N__46470));
    LocalMux I__9608 (
            .O(N__46588),
            .I(N__46470));
    LocalMux I__9607 (
            .O(N__46573),
            .I(N__46470));
    LocalMux I__9606 (
            .O(N__46558),
            .I(N__46470));
    InMux I__9605 (
            .O(N__46557),
            .I(N__46455));
    InMux I__9604 (
            .O(N__46554),
            .I(N__46455));
    InMux I__9603 (
            .O(N__46553),
            .I(N__46455));
    InMux I__9602 (
            .O(N__46550),
            .I(N__46455));
    InMux I__9601 (
            .O(N__46549),
            .I(N__46455));
    InMux I__9600 (
            .O(N__46546),
            .I(N__46455));
    InMux I__9599 (
            .O(N__46545),
            .I(N__46455));
    InMux I__9598 (
            .O(N__46544),
            .I(N__46440));
    InMux I__9597 (
            .O(N__46541),
            .I(N__46440));
    InMux I__9596 (
            .O(N__46540),
            .I(N__46440));
    InMux I__9595 (
            .O(N__46537),
            .I(N__46440));
    InMux I__9594 (
            .O(N__46536),
            .I(N__46440));
    InMux I__9593 (
            .O(N__46533),
            .I(N__46440));
    InMux I__9592 (
            .O(N__46532),
            .I(N__46440));
    InMux I__9591 (
            .O(N__46531),
            .I(N__46433));
    InMux I__9590 (
            .O(N__46530),
            .I(N__46433));
    InMux I__9589 (
            .O(N__46529),
            .I(N__46433));
    InMux I__9588 (
            .O(N__46528),
            .I(N__46424));
    InMux I__9587 (
            .O(N__46527),
            .I(N__46424));
    InMux I__9586 (
            .O(N__46526),
            .I(N__46424));
    InMux I__9585 (
            .O(N__46525),
            .I(N__46424));
    InMux I__9584 (
            .O(N__46524),
            .I(N__46417));
    InMux I__9583 (
            .O(N__46523),
            .I(N__46417));
    InMux I__9582 (
            .O(N__46522),
            .I(N__46417));
    InMux I__9581 (
            .O(N__46521),
            .I(N__46408));
    InMux I__9580 (
            .O(N__46520),
            .I(N__46408));
    InMux I__9579 (
            .O(N__46519),
            .I(N__46408));
    InMux I__9578 (
            .O(N__46518),
            .I(N__46408));
    InMux I__9577 (
            .O(N__46517),
            .I(N__46401));
    InMux I__9576 (
            .O(N__46516),
            .I(N__46401));
    InMux I__9575 (
            .O(N__46515),
            .I(N__46401));
    InMux I__9574 (
            .O(N__46514),
            .I(N__46392));
    InMux I__9573 (
            .O(N__46513),
            .I(N__46392));
    InMux I__9572 (
            .O(N__46512),
            .I(N__46392));
    InMux I__9571 (
            .O(N__46511),
            .I(N__46392));
    CascadeMux I__9570 (
            .O(N__46510),
            .I(N__46388));
    CascadeMux I__9569 (
            .O(N__46509),
            .I(N__46384));
    CascadeMux I__9568 (
            .O(N__46508),
            .I(N__46380));
    InMux I__9567 (
            .O(N__46507),
            .I(N__46364));
    InMux I__9566 (
            .O(N__46504),
            .I(N__46364));
    InMux I__9565 (
            .O(N__46503),
            .I(N__46364));
    InMux I__9564 (
            .O(N__46500),
            .I(N__46364));
    InMux I__9563 (
            .O(N__46499),
            .I(N__46364));
    InMux I__9562 (
            .O(N__46496),
            .I(N__46364));
    InMux I__9561 (
            .O(N__46495),
            .I(N__46364));
    CascadeMux I__9560 (
            .O(N__46494),
            .I(N__46360));
    CascadeMux I__9559 (
            .O(N__46493),
            .I(N__46356));
    CascadeMux I__9558 (
            .O(N__46492),
            .I(N__46352));
    InMux I__9557 (
            .O(N__46491),
            .I(N__46336));
    InMux I__9556 (
            .O(N__46488),
            .I(N__46336));
    InMux I__9555 (
            .O(N__46487),
            .I(N__46336));
    InMux I__9554 (
            .O(N__46484),
            .I(N__46336));
    InMux I__9553 (
            .O(N__46483),
            .I(N__46336));
    InMux I__9552 (
            .O(N__46480),
            .I(N__46336));
    InMux I__9551 (
            .O(N__46479),
            .I(N__46336));
    Span4Mux_v I__9550 (
            .O(N__46470),
            .I(N__46329));
    LocalMux I__9549 (
            .O(N__46455),
            .I(N__46329));
    LocalMux I__9548 (
            .O(N__46440),
            .I(N__46329));
    LocalMux I__9547 (
            .O(N__46433),
            .I(N__46316));
    LocalMux I__9546 (
            .O(N__46424),
            .I(N__46316));
    LocalMux I__9545 (
            .O(N__46417),
            .I(N__46316));
    LocalMux I__9544 (
            .O(N__46408),
            .I(N__46316));
    LocalMux I__9543 (
            .O(N__46401),
            .I(N__46316));
    LocalMux I__9542 (
            .O(N__46392),
            .I(N__46316));
    InMux I__9541 (
            .O(N__46391),
            .I(N__46301));
    InMux I__9540 (
            .O(N__46388),
            .I(N__46301));
    InMux I__9539 (
            .O(N__46387),
            .I(N__46301));
    InMux I__9538 (
            .O(N__46384),
            .I(N__46301));
    InMux I__9537 (
            .O(N__46383),
            .I(N__46301));
    InMux I__9536 (
            .O(N__46380),
            .I(N__46301));
    InMux I__9535 (
            .O(N__46379),
            .I(N__46301));
    LocalMux I__9534 (
            .O(N__46364),
            .I(N__46298));
    InMux I__9533 (
            .O(N__46363),
            .I(N__46283));
    InMux I__9532 (
            .O(N__46360),
            .I(N__46283));
    InMux I__9531 (
            .O(N__46359),
            .I(N__46283));
    InMux I__9530 (
            .O(N__46356),
            .I(N__46283));
    InMux I__9529 (
            .O(N__46355),
            .I(N__46283));
    InMux I__9528 (
            .O(N__46352),
            .I(N__46283));
    InMux I__9527 (
            .O(N__46351),
            .I(N__46283));
    LocalMux I__9526 (
            .O(N__46336),
            .I(N__46259));
    Span4Mux_v I__9525 (
            .O(N__46329),
            .I(N__46252));
    Span4Mux_v I__9524 (
            .O(N__46316),
            .I(N__46252));
    LocalMux I__9523 (
            .O(N__46301),
            .I(N__46252));
    Span4Mux_v I__9522 (
            .O(N__46298),
            .I(N__46247));
    LocalMux I__9521 (
            .O(N__46283),
            .I(N__46247));
    InMux I__9520 (
            .O(N__46282),
            .I(N__46240));
    InMux I__9519 (
            .O(N__46281),
            .I(N__46240));
    InMux I__9518 (
            .O(N__46280),
            .I(N__46240));
    InMux I__9517 (
            .O(N__46279),
            .I(N__46231));
    InMux I__9516 (
            .O(N__46278),
            .I(N__46231));
    InMux I__9515 (
            .O(N__46277),
            .I(N__46231));
    InMux I__9514 (
            .O(N__46276),
            .I(N__46231));
    InMux I__9513 (
            .O(N__46275),
            .I(N__46224));
    InMux I__9512 (
            .O(N__46274),
            .I(N__46224));
    InMux I__9511 (
            .O(N__46273),
            .I(N__46224));
    InMux I__9510 (
            .O(N__46272),
            .I(N__46215));
    InMux I__9509 (
            .O(N__46271),
            .I(N__46215));
    InMux I__9508 (
            .O(N__46270),
            .I(N__46215));
    InMux I__9507 (
            .O(N__46269),
            .I(N__46215));
    InMux I__9506 (
            .O(N__46268),
            .I(N__46208));
    InMux I__9505 (
            .O(N__46267),
            .I(N__46208));
    InMux I__9504 (
            .O(N__46266),
            .I(N__46208));
    InMux I__9503 (
            .O(N__46265),
            .I(N__46199));
    InMux I__9502 (
            .O(N__46264),
            .I(N__46199));
    InMux I__9501 (
            .O(N__46263),
            .I(N__46199));
    InMux I__9500 (
            .O(N__46262),
            .I(N__46199));
    Odrv4 I__9499 (
            .O(N__46259),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__9498 (
            .O(N__46252),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__9497 (
            .O(N__46247),
            .I(CONSTANT_ONE_NET));
    LocalMux I__9496 (
            .O(N__46240),
            .I(CONSTANT_ONE_NET));
    LocalMux I__9495 (
            .O(N__46231),
            .I(CONSTANT_ONE_NET));
    LocalMux I__9494 (
            .O(N__46224),
            .I(CONSTANT_ONE_NET));
    LocalMux I__9493 (
            .O(N__46215),
            .I(CONSTANT_ONE_NET));
    LocalMux I__9492 (
            .O(N__46208),
            .I(CONSTANT_ONE_NET));
    LocalMux I__9491 (
            .O(N__46199),
            .I(CONSTANT_ONE_NET));
    InMux I__9490 (
            .O(N__46180),
            .I(bfn_19_32_0_));
    CascadeMux I__9489 (
            .O(N__46177),
            .I(N__46171));
    InMux I__9488 (
            .O(N__46176),
            .I(N__46168));
    CascadeMux I__9487 (
            .O(N__46175),
            .I(N__46165));
    CascadeMux I__9486 (
            .O(N__46174),
            .I(N__46162));
    InMux I__9485 (
            .O(N__46171),
            .I(N__46159));
    LocalMux I__9484 (
            .O(N__46168),
            .I(N__46155));
    InMux I__9483 (
            .O(N__46165),
            .I(N__46152));
    InMux I__9482 (
            .O(N__46162),
            .I(N__46149));
    LocalMux I__9481 (
            .O(N__46159),
            .I(N__46144));
    InMux I__9480 (
            .O(N__46158),
            .I(N__46141));
    Span4Mux_v I__9479 (
            .O(N__46155),
            .I(N__46138));
    LocalMux I__9478 (
            .O(N__46152),
            .I(N__46135));
    LocalMux I__9477 (
            .O(N__46149),
            .I(N__46132));
    InMux I__9476 (
            .O(N__46148),
            .I(N__46129));
    InMux I__9475 (
            .O(N__46147),
            .I(N__46126));
    Span4Mux_h I__9474 (
            .O(N__46144),
            .I(N__46121));
    LocalMux I__9473 (
            .O(N__46141),
            .I(N__46121));
    Span4Mux_h I__9472 (
            .O(N__46138),
            .I(N__46116));
    Span4Mux_v I__9471 (
            .O(N__46135),
            .I(N__46116));
    Span4Mux_h I__9470 (
            .O(N__46132),
            .I(N__46113));
    LocalMux I__9469 (
            .O(N__46129),
            .I(N__46110));
    LocalMux I__9468 (
            .O(N__46126),
            .I(N__46104));
    Span4Mux_h I__9467 (
            .O(N__46121),
            .I(N__46104));
    Span4Mux_h I__9466 (
            .O(N__46116),
            .I(N__46099));
    Span4Mux_v I__9465 (
            .O(N__46113),
            .I(N__46099));
    Span12Mux_h I__9464 (
            .O(N__46110),
            .I(N__46096));
    InMux I__9463 (
            .O(N__46109),
            .I(N__46093));
    Sp12to4 I__9462 (
            .O(N__46104),
            .I(N__46090));
    Span4Mux_v I__9461 (
            .O(N__46099),
            .I(N__46087));
    Span12Mux_v I__9460 (
            .O(N__46096),
            .I(N__46084));
    LocalMux I__9459 (
            .O(N__46093),
            .I(\c0.FRAME_MATCHER_i_31 ));
    Odrv12 I__9458 (
            .O(N__46090),
            .I(\c0.FRAME_MATCHER_i_31 ));
    Odrv4 I__9457 (
            .O(N__46087),
            .I(\c0.FRAME_MATCHER_i_31 ));
    Odrv12 I__9456 (
            .O(N__46084),
            .I(\c0.FRAME_MATCHER_i_31 ));
    SRMux I__9455 (
            .O(N__46075),
            .I(N__46072));
    LocalMux I__9454 (
            .O(N__46072),
            .I(N__46069));
    Span4Mux_s1_v I__9453 (
            .O(N__46069),
            .I(N__46066));
    Span4Mux_v I__9452 (
            .O(N__46066),
            .I(N__46063));
    Odrv4 I__9451 (
            .O(N__46063),
            .I(\c0.n3_adj_4421 ));
    SRMux I__9450 (
            .O(N__46060),
            .I(N__46057));
    LocalMux I__9449 (
            .O(N__46057),
            .I(\c0.n3_adj_4475 ));
    InMux I__9448 (
            .O(N__46054),
            .I(N__46051));
    LocalMux I__9447 (
            .O(N__46051),
            .I(N__46045));
    InMux I__9446 (
            .O(N__46050),
            .I(N__46040));
    InMux I__9445 (
            .O(N__46049),
            .I(N__46040));
    InMux I__9444 (
            .O(N__46048),
            .I(N__46036));
    Span4Mux_h I__9443 (
            .O(N__46045),
            .I(N__46031));
    LocalMux I__9442 (
            .O(N__46040),
            .I(N__46031));
    InMux I__9441 (
            .O(N__46039),
            .I(N__46027));
    LocalMux I__9440 (
            .O(N__46036),
            .I(N__46024));
    Span4Mux_v I__9439 (
            .O(N__46031),
            .I(N__46021));
    InMux I__9438 (
            .O(N__46030),
            .I(N__46018));
    LocalMux I__9437 (
            .O(N__46027),
            .I(N__46015));
    Span4Mux_v I__9436 (
            .O(N__46024),
            .I(N__46011));
    Span4Mux_v I__9435 (
            .O(N__46021),
            .I(N__46006));
    LocalMux I__9434 (
            .O(N__46018),
            .I(N__46006));
    Span4Mux_h I__9433 (
            .O(N__46015),
            .I(N__46003));
    CascadeMux I__9432 (
            .O(N__46014),
            .I(N__46000));
    Span4Mux_v I__9431 (
            .O(N__46011),
            .I(N__45996));
    Span4Mux_h I__9430 (
            .O(N__46006),
            .I(N__45993));
    Sp12to4 I__9429 (
            .O(N__46003),
            .I(N__45990));
    InMux I__9428 (
            .O(N__46000),
            .I(N__45987));
    InMux I__9427 (
            .O(N__45999),
            .I(N__45984));
    Span4Mux_v I__9426 (
            .O(N__45996),
            .I(N__45981));
    Span4Mux_v I__9425 (
            .O(N__45993),
            .I(N__45978));
    Span12Mux_v I__9424 (
            .O(N__45990),
            .I(N__45975));
    LocalMux I__9423 (
            .O(N__45987),
            .I(\c0.FRAME_MATCHER_i_3 ));
    LocalMux I__9422 (
            .O(N__45984),
            .I(\c0.FRAME_MATCHER_i_3 ));
    Odrv4 I__9421 (
            .O(N__45981),
            .I(\c0.FRAME_MATCHER_i_3 ));
    Odrv4 I__9420 (
            .O(N__45978),
            .I(\c0.FRAME_MATCHER_i_3 ));
    Odrv12 I__9419 (
            .O(N__45975),
            .I(\c0.FRAME_MATCHER_i_3 ));
    SRMux I__9418 (
            .O(N__45964),
            .I(N__45961));
    LocalMux I__9417 (
            .O(N__45961),
            .I(N__45958));
    Odrv4 I__9416 (
            .O(N__45958),
            .I(\c0.n3_adj_4472 ));
    SRMux I__9415 (
            .O(N__45955),
            .I(N__45952));
    LocalMux I__9414 (
            .O(N__45952),
            .I(N__45949));
    Span4Mux_s3_v I__9413 (
            .O(N__45949),
            .I(N__45946));
    Odrv4 I__9412 (
            .O(N__45946),
            .I(\c0.n3_adj_4428 ));
    InMux I__9411 (
            .O(N__45943),
            .I(N__45937));
    InMux I__9410 (
            .O(N__45942),
            .I(N__45937));
    LocalMux I__9409 (
            .O(N__45937),
            .I(N__45933));
    InMux I__9408 (
            .O(N__45936),
            .I(N__45930));
    Span4Mux_v I__9407 (
            .O(N__45933),
            .I(N__45927));
    LocalMux I__9406 (
            .O(N__45930),
            .I(\c0.FRAME_MATCHER_i_30 ));
    Odrv4 I__9405 (
            .O(N__45927),
            .I(\c0.FRAME_MATCHER_i_30 ));
    InMux I__9404 (
            .O(N__45922),
            .I(bfn_19_31_0_));
    SRMux I__9403 (
            .O(N__45919),
            .I(N__45916));
    LocalMux I__9402 (
            .O(N__45916),
            .I(N__45913));
    Span4Mux_v I__9401 (
            .O(N__45913),
            .I(N__45910));
    Odrv4 I__9400 (
            .O(N__45910),
            .I(\c0.n3_adj_4426 ));
    InMux I__9399 (
            .O(N__45907),
            .I(bfn_19_29_0_));
    InMux I__9398 (
            .O(N__45904),
            .I(N__45900));
    InMux I__9397 (
            .O(N__45903),
            .I(N__45897));
    LocalMux I__9396 (
            .O(N__45900),
            .I(N__45891));
    LocalMux I__9395 (
            .O(N__45897),
            .I(N__45891));
    InMux I__9394 (
            .O(N__45896),
            .I(N__45888));
    Span4Mux_v I__9393 (
            .O(N__45891),
            .I(N__45885));
    LocalMux I__9392 (
            .O(N__45888),
            .I(\c0.FRAME_MATCHER_i_29 ));
    Odrv4 I__9391 (
            .O(N__45885),
            .I(\c0.FRAME_MATCHER_i_29 ));
    InMux I__9390 (
            .O(N__45880),
            .I(bfn_19_30_0_));
    InMux I__9389 (
            .O(N__45877),
            .I(N__45873));
    CascadeMux I__9388 (
            .O(N__45876),
            .I(N__45870));
    LocalMux I__9387 (
            .O(N__45873),
            .I(N__45866));
    InMux I__9386 (
            .O(N__45870),
            .I(N__45863));
    InMux I__9385 (
            .O(N__45869),
            .I(N__45860));
    Sp12to4 I__9384 (
            .O(N__45866),
            .I(N__45857));
    LocalMux I__9383 (
            .O(N__45863),
            .I(\c0.FRAME_MATCHER_i_27 ));
    LocalMux I__9382 (
            .O(N__45860),
            .I(\c0.FRAME_MATCHER_i_27 ));
    Odrv12 I__9381 (
            .O(N__45857),
            .I(\c0.FRAME_MATCHER_i_27 ));
    InMux I__9380 (
            .O(N__45850),
            .I(bfn_19_28_0_));
    SRMux I__9379 (
            .O(N__45847),
            .I(N__45844));
    LocalMux I__9378 (
            .O(N__45844),
            .I(N__45841));
    Odrv4 I__9377 (
            .O(N__45841),
            .I(\c0.n3_adj_4432 ));
    InMux I__9376 (
            .O(N__45838),
            .I(N__45834));
    CascadeMux I__9375 (
            .O(N__45837),
            .I(N__45831));
    LocalMux I__9374 (
            .O(N__45834),
            .I(N__45827));
    InMux I__9373 (
            .O(N__45831),
            .I(N__45824));
    InMux I__9372 (
            .O(N__45830),
            .I(N__45821));
    Span4Mux_v I__9371 (
            .O(N__45827),
            .I(N__45818));
    LocalMux I__9370 (
            .O(N__45824),
            .I(\c0.FRAME_MATCHER_i_26 ));
    LocalMux I__9369 (
            .O(N__45821),
            .I(\c0.FRAME_MATCHER_i_26 ));
    Odrv4 I__9368 (
            .O(N__45818),
            .I(\c0.FRAME_MATCHER_i_26 ));
    InMux I__9367 (
            .O(N__45811),
            .I(bfn_19_27_0_));
    SRMux I__9366 (
            .O(N__45808),
            .I(N__45805));
    LocalMux I__9365 (
            .O(N__45805),
            .I(\c0.n3_adj_4433 ));
    CascadeMux I__9364 (
            .O(N__45802),
            .I(N__45799));
    InMux I__9363 (
            .O(N__45799),
            .I(N__45795));
    CascadeMux I__9362 (
            .O(N__45798),
            .I(N__45792));
    LocalMux I__9361 (
            .O(N__45795),
            .I(N__45788));
    InMux I__9360 (
            .O(N__45792),
            .I(N__45785));
    InMux I__9359 (
            .O(N__45791),
            .I(N__45782));
    Span4Mux_v I__9358 (
            .O(N__45788),
            .I(N__45779));
    LocalMux I__9357 (
            .O(N__45785),
            .I(\c0.FRAME_MATCHER_i_25 ));
    LocalMux I__9356 (
            .O(N__45782),
            .I(\c0.FRAME_MATCHER_i_25 ));
    Odrv4 I__9355 (
            .O(N__45779),
            .I(\c0.FRAME_MATCHER_i_25 ));
    InMux I__9354 (
            .O(N__45772),
            .I(bfn_19_26_0_));
    SRMux I__9353 (
            .O(N__45769),
            .I(N__45766));
    LocalMux I__9352 (
            .O(N__45766),
            .I(N__45763));
    Odrv4 I__9351 (
            .O(N__45763),
            .I(\c0.n3_adj_4434 ));
    CascadeMux I__9350 (
            .O(N__45760),
            .I(N__45756));
    CascadeMux I__9349 (
            .O(N__45759),
            .I(N__45753));
    InMux I__9348 (
            .O(N__45756),
            .I(N__45750));
    InMux I__9347 (
            .O(N__45753),
            .I(N__45746));
    LocalMux I__9346 (
            .O(N__45750),
            .I(N__45743));
    InMux I__9345 (
            .O(N__45749),
            .I(N__45740));
    LocalMux I__9344 (
            .O(N__45746),
            .I(N__45737));
    Odrv4 I__9343 (
            .O(N__45743),
            .I(\c0.FRAME_MATCHER_i_24 ));
    LocalMux I__9342 (
            .O(N__45740),
            .I(\c0.FRAME_MATCHER_i_24 ));
    Odrv4 I__9341 (
            .O(N__45737),
            .I(\c0.FRAME_MATCHER_i_24 ));
    InMux I__9340 (
            .O(N__45730),
            .I(bfn_19_25_0_));
    SRMux I__9339 (
            .O(N__45727),
            .I(N__45724));
    LocalMux I__9338 (
            .O(N__45724),
            .I(N__45721));
    Span4Mux_h I__9337 (
            .O(N__45721),
            .I(N__45718));
    Odrv4 I__9336 (
            .O(N__45718),
            .I(\c0.n3_adj_4435 ));
    InMux I__9335 (
            .O(N__45715),
            .I(N__45711));
    CascadeMux I__9334 (
            .O(N__45714),
            .I(N__45708));
    LocalMux I__9333 (
            .O(N__45711),
            .I(N__45704));
    InMux I__9332 (
            .O(N__45708),
            .I(N__45701));
    InMux I__9331 (
            .O(N__45707),
            .I(N__45698));
    Span4Mux_h I__9330 (
            .O(N__45704),
            .I(N__45695));
    LocalMux I__9329 (
            .O(N__45701),
            .I(\c0.FRAME_MATCHER_i_23 ));
    LocalMux I__9328 (
            .O(N__45698),
            .I(\c0.FRAME_MATCHER_i_23 ));
    Odrv4 I__9327 (
            .O(N__45695),
            .I(\c0.FRAME_MATCHER_i_23 ));
    InMux I__9326 (
            .O(N__45688),
            .I(bfn_19_24_0_));
    SRMux I__9325 (
            .O(N__45685),
            .I(N__45682));
    LocalMux I__9324 (
            .O(N__45682),
            .I(N__45679));
    Odrv12 I__9323 (
            .O(N__45679),
            .I(\c0.n3_adj_4436 ));
    InMux I__9322 (
            .O(N__45676),
            .I(N__45671));
    InMux I__9321 (
            .O(N__45675),
            .I(N__45668));
    InMux I__9320 (
            .O(N__45674),
            .I(N__45665));
    LocalMux I__9319 (
            .O(N__45671),
            .I(N__45662));
    LocalMux I__9318 (
            .O(N__45668),
            .I(\c0.FRAME_MATCHER_i_22 ));
    LocalMux I__9317 (
            .O(N__45665),
            .I(\c0.FRAME_MATCHER_i_22 ));
    Odrv4 I__9316 (
            .O(N__45662),
            .I(\c0.FRAME_MATCHER_i_22 ));
    InMux I__9315 (
            .O(N__45655),
            .I(bfn_19_23_0_));
    SRMux I__9314 (
            .O(N__45652),
            .I(N__45649));
    LocalMux I__9313 (
            .O(N__45649),
            .I(N__45646));
    Span4Mux_h I__9312 (
            .O(N__45646),
            .I(N__45643));
    Odrv4 I__9311 (
            .O(N__45643),
            .I(\c0.n3_adj_4438 ));
    CascadeMux I__9310 (
            .O(N__45640),
            .I(N__45637));
    InMux I__9309 (
            .O(N__45637),
            .I(N__45634));
    LocalMux I__9308 (
            .O(N__45634),
            .I(N__45631));
    Span4Mux_h I__9307 (
            .O(N__45631),
            .I(N__45626));
    InMux I__9306 (
            .O(N__45630),
            .I(N__45623));
    InMux I__9305 (
            .O(N__45629),
            .I(N__45620));
    Odrv4 I__9304 (
            .O(N__45626),
            .I(\c0.FRAME_MATCHER_i_21 ));
    LocalMux I__9303 (
            .O(N__45623),
            .I(\c0.FRAME_MATCHER_i_21 ));
    LocalMux I__9302 (
            .O(N__45620),
            .I(\c0.FRAME_MATCHER_i_21 ));
    InMux I__9301 (
            .O(N__45613),
            .I(bfn_19_22_0_));
    SRMux I__9300 (
            .O(N__45610),
            .I(N__45607));
    LocalMux I__9299 (
            .O(N__45607),
            .I(N__45604));
    Odrv4 I__9298 (
            .O(N__45604),
            .I(\c0.n3_adj_4440 ));
    SRMux I__9297 (
            .O(N__45601),
            .I(N__45598));
    LocalMux I__9296 (
            .O(N__45598),
            .I(N__45595));
    Span4Mux_h I__9295 (
            .O(N__45595),
            .I(N__45592));
    Span4Mux_h I__9294 (
            .O(N__45592),
            .I(N__45589));
    Odrv4 I__9293 (
            .O(N__45589),
            .I(\c0.n3_adj_4444 ));
    InMux I__9292 (
            .O(N__45586),
            .I(bfn_19_21_0_));
    CascadeMux I__9291 (
            .O(N__45583),
            .I(N__45580));
    InMux I__9290 (
            .O(N__45580),
            .I(N__45576));
    InMux I__9289 (
            .O(N__45579),
            .I(N__45573));
    LocalMux I__9288 (
            .O(N__45576),
            .I(N__45570));
    LocalMux I__9287 (
            .O(N__45573),
            .I(N__45566));
    Span4Mux_h I__9286 (
            .O(N__45570),
            .I(N__45563));
    InMux I__9285 (
            .O(N__45569),
            .I(N__45560));
    Span4Mux_h I__9284 (
            .O(N__45566),
            .I(N__45557));
    Odrv4 I__9283 (
            .O(N__45563),
            .I(\c0.FRAME_MATCHER_i_18 ));
    LocalMux I__9282 (
            .O(N__45560),
            .I(\c0.FRAME_MATCHER_i_18 ));
    Odrv4 I__9281 (
            .O(N__45557),
            .I(\c0.FRAME_MATCHER_i_18 ));
    InMux I__9280 (
            .O(N__45550),
            .I(bfn_19_19_0_));
    SRMux I__9279 (
            .O(N__45547),
            .I(N__45544));
    LocalMux I__9278 (
            .O(N__45544),
            .I(N__45541));
    Span4Mux_v I__9277 (
            .O(N__45541),
            .I(N__45538));
    Odrv4 I__9276 (
            .O(N__45538),
            .I(\c0.n3_adj_4446 ));
    CascadeMux I__9275 (
            .O(N__45535),
            .I(N__45531));
    InMux I__9274 (
            .O(N__45534),
            .I(N__45528));
    InMux I__9273 (
            .O(N__45531),
            .I(N__45525));
    LocalMux I__9272 (
            .O(N__45528),
            .I(N__45521));
    LocalMux I__9271 (
            .O(N__45525),
            .I(N__45518));
    InMux I__9270 (
            .O(N__45524),
            .I(N__45515));
    Span4Mux_v I__9269 (
            .O(N__45521),
            .I(N__45512));
    Odrv4 I__9268 (
            .O(N__45518),
            .I(\c0.FRAME_MATCHER_i_19 ));
    LocalMux I__9267 (
            .O(N__45515),
            .I(\c0.FRAME_MATCHER_i_19 ));
    Odrv4 I__9266 (
            .O(N__45512),
            .I(\c0.FRAME_MATCHER_i_19 ));
    InMux I__9265 (
            .O(N__45505),
            .I(bfn_19_20_0_));
    CascadeMux I__9264 (
            .O(N__45502),
            .I(N__45499));
    InMux I__9263 (
            .O(N__45499),
            .I(N__45495));
    InMux I__9262 (
            .O(N__45498),
            .I(N__45492));
    LocalMux I__9261 (
            .O(N__45495),
            .I(N__45488));
    LocalMux I__9260 (
            .O(N__45492),
            .I(N__45485));
    InMux I__9259 (
            .O(N__45491),
            .I(N__45482));
    Span4Mux_v I__9258 (
            .O(N__45488),
            .I(N__45477));
    Span4Mux_v I__9257 (
            .O(N__45485),
            .I(N__45477));
    LocalMux I__9256 (
            .O(N__45482),
            .I(\c0.FRAME_MATCHER_i_17 ));
    Odrv4 I__9255 (
            .O(N__45477),
            .I(\c0.FRAME_MATCHER_i_17 ));
    InMux I__9254 (
            .O(N__45472),
            .I(bfn_19_18_0_));
    SRMux I__9253 (
            .O(N__45469),
            .I(N__45466));
    LocalMux I__9252 (
            .O(N__45466),
            .I(N__45463));
    Span4Mux_h I__9251 (
            .O(N__45463),
            .I(N__45460));
    Span4Mux_v I__9250 (
            .O(N__45460),
            .I(N__45457));
    Odrv4 I__9249 (
            .O(N__45457),
            .I(\c0.n3_adj_4448 ));
    InMux I__9248 (
            .O(N__45454),
            .I(bfn_19_17_0_));
    SRMux I__9247 (
            .O(N__45451),
            .I(N__45448));
    LocalMux I__9246 (
            .O(N__45448),
            .I(N__45445));
    Odrv12 I__9245 (
            .O(N__45445),
            .I(\c0.n3_adj_4450 ));
    InMux I__9244 (
            .O(N__45442),
            .I(bfn_19_16_0_));
    CascadeMux I__9243 (
            .O(N__45439),
            .I(N__45436));
    InMux I__9242 (
            .O(N__45436),
            .I(N__45432));
    InMux I__9241 (
            .O(N__45435),
            .I(N__45429));
    LocalMux I__9240 (
            .O(N__45432),
            .I(N__45426));
    LocalMux I__9239 (
            .O(N__45429),
            .I(N__45422));
    Span4Mux_h I__9238 (
            .O(N__45426),
            .I(N__45419));
    InMux I__9237 (
            .O(N__45425),
            .I(N__45416));
    Span4Mux_v I__9236 (
            .O(N__45422),
            .I(N__45413));
    Odrv4 I__9235 (
            .O(N__45419),
            .I(\c0.FRAME_MATCHER_i_14 ));
    LocalMux I__9234 (
            .O(N__45416),
            .I(\c0.FRAME_MATCHER_i_14 ));
    Odrv4 I__9233 (
            .O(N__45413),
            .I(\c0.FRAME_MATCHER_i_14 ));
    InMux I__9232 (
            .O(N__45406),
            .I(bfn_19_15_0_));
    SRMux I__9231 (
            .O(N__45403),
            .I(N__45400));
    LocalMux I__9230 (
            .O(N__45400),
            .I(N__45397));
    Span4Mux_v I__9229 (
            .O(N__45397),
            .I(N__45394));
    Sp12to4 I__9228 (
            .O(N__45394),
            .I(N__45391));
    Odrv12 I__9227 (
            .O(N__45391),
            .I(\c0.n3_adj_4453 ));
    InMux I__9226 (
            .O(N__45388),
            .I(bfn_19_14_0_));
    CascadeMux I__9225 (
            .O(N__45385),
            .I(N__45381));
    CascadeMux I__9224 (
            .O(N__45384),
            .I(N__45378));
    InMux I__9223 (
            .O(N__45381),
            .I(N__45375));
    InMux I__9222 (
            .O(N__45378),
            .I(N__45372));
    LocalMux I__9221 (
            .O(N__45375),
            .I(N__45369));
    LocalMux I__9220 (
            .O(N__45372),
            .I(N__45366));
    Span4Mux_h I__9219 (
            .O(N__45369),
            .I(N__45363));
    Span4Mux_h I__9218 (
            .O(N__45366),
            .I(N__45359));
    Span4Mux_v I__9217 (
            .O(N__45363),
            .I(N__45356));
    InMux I__9216 (
            .O(N__45362),
            .I(N__45353));
    Odrv4 I__9215 (
            .O(N__45359),
            .I(\c0.FRAME_MATCHER_i_12 ));
    Odrv4 I__9214 (
            .O(N__45356),
            .I(\c0.FRAME_MATCHER_i_12 ));
    LocalMux I__9213 (
            .O(N__45353),
            .I(\c0.FRAME_MATCHER_i_12 ));
    InMux I__9212 (
            .O(N__45346),
            .I(bfn_19_13_0_));
    SRMux I__9211 (
            .O(N__45343),
            .I(N__45340));
    LocalMux I__9210 (
            .O(N__45340),
            .I(N__45337));
    Span4Mux_v I__9209 (
            .O(N__45337),
            .I(N__45334));
    Odrv4 I__9208 (
            .O(N__45334),
            .I(\c0.n3_adj_4456 ));
    InMux I__9207 (
            .O(N__45331),
            .I(N__45328));
    LocalMux I__9206 (
            .O(N__45328),
            .I(N__45324));
    InMux I__9205 (
            .O(N__45327),
            .I(N__45321));
    Sp12to4 I__9204 (
            .O(N__45324),
            .I(N__45318));
    LocalMux I__9203 (
            .O(N__45321),
            .I(N__45315));
    Span12Mux_h I__9202 (
            .O(N__45318),
            .I(N__45309));
    Sp12to4 I__9201 (
            .O(N__45315),
            .I(N__45309));
    InMux I__9200 (
            .O(N__45314),
            .I(N__45306));
    Odrv12 I__9199 (
            .O(N__45309),
            .I(\c0.FRAME_MATCHER_i_11 ));
    LocalMux I__9198 (
            .O(N__45306),
            .I(\c0.FRAME_MATCHER_i_11 ));
    InMux I__9197 (
            .O(N__45301),
            .I(bfn_19_12_0_));
    SRMux I__9196 (
            .O(N__45298),
            .I(N__45295));
    LocalMux I__9195 (
            .O(N__45295),
            .I(N__45292));
    Span4Mux_h I__9194 (
            .O(N__45292),
            .I(N__45289));
    Span4Mux_v I__9193 (
            .O(N__45289),
            .I(N__45286));
    Span4Mux_v I__9192 (
            .O(N__45286),
            .I(N__45283));
    Odrv4 I__9191 (
            .O(N__45283),
            .I(\c0.n3_adj_4458 ));
    CascadeMux I__9190 (
            .O(N__45280),
            .I(N__45276));
    InMux I__9189 (
            .O(N__45279),
            .I(N__45273));
    InMux I__9188 (
            .O(N__45276),
            .I(N__45270));
    LocalMux I__9187 (
            .O(N__45273),
            .I(N__45267));
    LocalMux I__9186 (
            .O(N__45270),
            .I(N__45261));
    Span4Mux_v I__9185 (
            .O(N__45267),
            .I(N__45261));
    InMux I__9184 (
            .O(N__45266),
            .I(N__45258));
    Sp12to4 I__9183 (
            .O(N__45261),
            .I(N__45255));
    LocalMux I__9182 (
            .O(N__45258),
            .I(\c0.FRAME_MATCHER_i_9 ));
    Odrv12 I__9181 (
            .O(N__45255),
            .I(\c0.FRAME_MATCHER_i_9 ));
    InMux I__9180 (
            .O(N__45250),
            .I(bfn_19_10_0_));
    SRMux I__9179 (
            .O(N__45247),
            .I(N__45244));
    LocalMux I__9178 (
            .O(N__45244),
            .I(N__45241));
    Span4Mux_v I__9177 (
            .O(N__45241),
            .I(N__45238));
    Span4Mux_h I__9176 (
            .O(N__45238),
            .I(N__45235));
    Odrv4 I__9175 (
            .O(N__45235),
            .I(\c0.n3_adj_4462 ));
    InMux I__9174 (
            .O(N__45232),
            .I(bfn_19_11_0_));
    InMux I__9173 (
            .O(N__45229),
            .I(N__45226));
    LocalMux I__9172 (
            .O(N__45226),
            .I(N__45222));
    InMux I__9171 (
            .O(N__45225),
            .I(N__45219));
    Span4Mux_v I__9170 (
            .O(N__45222),
            .I(N__45216));
    LocalMux I__9169 (
            .O(N__45219),
            .I(N__45212));
    Span4Mux_v I__9168 (
            .O(N__45216),
            .I(N__45209));
    InMux I__9167 (
            .O(N__45215),
            .I(N__45206));
    Sp12to4 I__9166 (
            .O(N__45212),
            .I(N__45203));
    Odrv4 I__9165 (
            .O(N__45209),
            .I(\c0.FRAME_MATCHER_i_8 ));
    LocalMux I__9164 (
            .O(N__45206),
            .I(\c0.FRAME_MATCHER_i_8 ));
    Odrv12 I__9163 (
            .O(N__45203),
            .I(\c0.FRAME_MATCHER_i_8 ));
    InMux I__9162 (
            .O(N__45196),
            .I(bfn_19_9_0_));
    SRMux I__9161 (
            .O(N__45193),
            .I(N__45190));
    LocalMux I__9160 (
            .O(N__45190),
            .I(N__45187));
    Span4Mux_h I__9159 (
            .O(N__45187),
            .I(N__45184));
    Span4Mux_v I__9158 (
            .O(N__45184),
            .I(N__45181));
    Odrv4 I__9157 (
            .O(N__45181),
            .I(\c0.n3_adj_4463 ));
    InMux I__9156 (
            .O(N__45178),
            .I(N__45175));
    LocalMux I__9155 (
            .O(N__45175),
            .I(N__45171));
    InMux I__9154 (
            .O(N__45174),
            .I(N__45168));
    Sp12to4 I__9153 (
            .O(N__45171),
            .I(N__45165));
    LocalMux I__9152 (
            .O(N__45168),
            .I(N__45162));
    Span12Mux_h I__9151 (
            .O(N__45165),
            .I(N__45159));
    Span4Mux_v I__9150 (
            .O(N__45162),
            .I(N__45156));
    Span12Mux_v I__9149 (
            .O(N__45159),
            .I(N__45152));
    Span4Mux_v I__9148 (
            .O(N__45156),
            .I(N__45149));
    InMux I__9147 (
            .O(N__45155),
            .I(N__45146));
    Odrv12 I__9146 (
            .O(N__45152),
            .I(\c0.FRAME_MATCHER_i_7 ));
    Odrv4 I__9145 (
            .O(N__45149),
            .I(\c0.FRAME_MATCHER_i_7 ));
    LocalMux I__9144 (
            .O(N__45146),
            .I(\c0.FRAME_MATCHER_i_7 ));
    InMux I__9143 (
            .O(N__45139),
            .I(bfn_19_8_0_));
    SRMux I__9142 (
            .O(N__45136),
            .I(N__45133));
    LocalMux I__9141 (
            .O(N__45133),
            .I(N__45130));
    Sp12to4 I__9140 (
            .O(N__45130),
            .I(N__45127));
    Span12Mux_h I__9139 (
            .O(N__45127),
            .I(N__45124));
    Span12Mux_v I__9138 (
            .O(N__45124),
            .I(N__45121));
    Odrv12 I__9137 (
            .O(N__45121),
            .I(\c0.n3_adj_4465 ));
    InMux I__9136 (
            .O(N__45118),
            .I(bfn_19_7_0_));
    SRMux I__9135 (
            .O(N__45115),
            .I(N__45112));
    LocalMux I__9134 (
            .O(N__45112),
            .I(N__45109));
    Span4Mux_v I__9133 (
            .O(N__45109),
            .I(N__45106));
    Span4Mux_v I__9132 (
            .O(N__45106),
            .I(N__45103));
    Odrv4 I__9131 (
            .O(N__45103),
            .I(\c0.n3_adj_4467 ));
    InMux I__9130 (
            .O(N__45100),
            .I(bfn_19_6_0_));
    SRMux I__9129 (
            .O(N__45097),
            .I(N__45094));
    LocalMux I__9128 (
            .O(N__45094),
            .I(N__45091));
    Span4Mux_v I__9127 (
            .O(N__45091),
            .I(N__45088));
    Odrv4 I__9126 (
            .O(N__45088),
            .I(\c0.n3_adj_4468 ));
    CascadeMux I__9125 (
            .O(N__45085),
            .I(N__45082));
    InMux I__9124 (
            .O(N__45082),
            .I(N__45078));
    InMux I__9123 (
            .O(N__45081),
            .I(N__45074));
    LocalMux I__9122 (
            .O(N__45078),
            .I(N__45070));
    CascadeMux I__9121 (
            .O(N__45077),
            .I(N__45066));
    LocalMux I__9120 (
            .O(N__45074),
            .I(N__45061));
    InMux I__9119 (
            .O(N__45073),
            .I(N__45058));
    Span4Mux_v I__9118 (
            .O(N__45070),
            .I(N__45055));
    InMux I__9117 (
            .O(N__45069),
            .I(N__45052));
    InMux I__9116 (
            .O(N__45066),
            .I(N__45049));
    InMux I__9115 (
            .O(N__45065),
            .I(N__45044));
    InMux I__9114 (
            .O(N__45064),
            .I(N__45044));
    Span4Mux_h I__9113 (
            .O(N__45061),
            .I(N__45039));
    LocalMux I__9112 (
            .O(N__45058),
            .I(N__45039));
    Span4Mux_h I__9111 (
            .O(N__45055),
            .I(N__45034));
    LocalMux I__9110 (
            .O(N__45052),
            .I(N__45034));
    LocalMux I__9109 (
            .O(N__45049),
            .I(N__45027));
    LocalMux I__9108 (
            .O(N__45044),
            .I(N__45027));
    Span4Mux_v I__9107 (
            .O(N__45039),
            .I(N__45027));
    Span4Mux_v I__9106 (
            .O(N__45034),
            .I(N__45022));
    Span4Mux_v I__9105 (
            .O(N__45027),
            .I(N__45022));
    Span4Mux_v I__9104 (
            .O(N__45022),
            .I(N__45019));
    Span4Mux_v I__9103 (
            .O(N__45019),
            .I(N__45015));
    InMux I__9102 (
            .O(N__45018),
            .I(N__45012));
    Odrv4 I__9101 (
            .O(N__45015),
            .I(\c0.FRAME_MATCHER_i_4 ));
    LocalMux I__9100 (
            .O(N__45012),
            .I(\c0.FRAME_MATCHER_i_4 ));
    InMux I__9099 (
            .O(N__45007),
            .I(bfn_19_5_0_));
    SRMux I__9098 (
            .O(N__45004),
            .I(N__45001));
    LocalMux I__9097 (
            .O(N__45001),
            .I(N__44998));
    Span4Mux_v I__9096 (
            .O(N__44998),
            .I(N__44995));
    Span4Mux_v I__9095 (
            .O(N__44995),
            .I(N__44992));
    Span4Mux_v I__9094 (
            .O(N__44992),
            .I(N__44989));
    Odrv4 I__9093 (
            .O(N__44989),
            .I(\c0.n3_adj_4470 ));
    InMux I__9092 (
            .O(N__44986),
            .I(bfn_19_4_0_));
    InMux I__9091 (
            .O(N__44983),
            .I(bfn_19_3_0_));
    SRMux I__9090 (
            .O(N__44980),
            .I(N__44977));
    LocalMux I__9089 (
            .O(N__44977),
            .I(N__44974));
    Span4Mux_s2_v I__9088 (
            .O(N__44974),
            .I(N__44971));
    Odrv4 I__9087 (
            .O(N__44971),
            .I(\c0.n3 ));
    InMux I__9086 (
            .O(N__44968),
            .I(bfn_19_2_0_));
    InMux I__9085 (
            .O(N__44965),
            .I(N__44962));
    LocalMux I__9084 (
            .O(N__44962),
            .I(N__44959));
    Span4Mux_h I__9083 (
            .O(N__44959),
            .I(N__44956));
    Odrv4 I__9082 (
            .O(N__44956),
            .I(\c0.n29_adj_4382 ));
    CascadeMux I__9081 (
            .O(N__44953),
            .I(N__44950));
    InMux I__9080 (
            .O(N__44950),
            .I(N__44947));
    LocalMux I__9079 (
            .O(N__44947),
            .I(N__44944));
    Span4Mux_s1_v I__9078 (
            .O(N__44944),
            .I(N__44941));
    Span4Mux_v I__9077 (
            .O(N__44941),
            .I(N__44938));
    Span4Mux_h I__9076 (
            .O(N__44938),
            .I(N__44935));
    Span4Mux_h I__9075 (
            .O(N__44935),
            .I(N__44932));
    Odrv4 I__9074 (
            .O(N__44932),
            .I(\c0.n161 ));
    InMux I__9073 (
            .O(N__44929),
            .I(N__44926));
    LocalMux I__9072 (
            .O(N__44926),
            .I(N__44922));
    InMux I__9071 (
            .O(N__44925),
            .I(N__44918));
    Span4Mux_h I__9070 (
            .O(N__44922),
            .I(N__44915));
    InMux I__9069 (
            .O(N__44921),
            .I(N__44912));
    LocalMux I__9068 (
            .O(N__44918),
            .I(data_in_frame_22_1));
    Odrv4 I__9067 (
            .O(N__44915),
            .I(data_in_frame_22_1));
    LocalMux I__9066 (
            .O(N__44912),
            .I(data_in_frame_22_1));
    CascadeMux I__9065 (
            .O(N__44905),
            .I(\c0.rx.n22611_cascade_ ));
    CascadeMux I__9064 (
            .O(N__44902),
            .I(\c0.rx.n8_cascade_ ));
    CascadeMux I__9063 (
            .O(N__44899),
            .I(N__44895));
    CascadeMux I__9062 (
            .O(N__44898),
            .I(N__44892));
    InMux I__9061 (
            .O(N__44895),
            .I(N__44889));
    InMux I__9060 (
            .O(N__44892),
            .I(N__44886));
    LocalMux I__9059 (
            .O(N__44889),
            .I(\c0.data_in_frame_29_2 ));
    LocalMux I__9058 (
            .O(N__44886),
            .I(\c0.data_in_frame_29_2 ));
    InMux I__9057 (
            .O(N__44881),
            .I(N__44877));
    InMux I__9056 (
            .O(N__44880),
            .I(N__44874));
    LocalMux I__9055 (
            .O(N__44877),
            .I(N__44871));
    LocalMux I__9054 (
            .O(N__44874),
            .I(\c0.data_in_frame_29_1 ));
    Odrv12 I__9053 (
            .O(N__44871),
            .I(\c0.data_in_frame_29_1 ));
    CascadeMux I__9052 (
            .O(N__44866),
            .I(\c0.n23388_cascade_ ));
    InMux I__9051 (
            .O(N__44863),
            .I(N__44860));
    LocalMux I__9050 (
            .O(N__44860),
            .I(\c0.n30_adj_4299 ));
    CascadeMux I__9049 (
            .O(N__44857),
            .I(\c0.n15_adj_4376_cascade_ ));
    InMux I__9048 (
            .O(N__44854),
            .I(N__44851));
    LocalMux I__9047 (
            .O(N__44851),
            .I(N__44848));
    Odrv12 I__9046 (
            .O(N__44848),
            .I(\c0.n17_adj_4378 ));
    CascadeMux I__9045 (
            .O(N__44845),
            .I(\c0.n18_adj_4379_cascade_ ));
    InMux I__9044 (
            .O(N__44842),
            .I(N__44839));
    LocalMux I__9043 (
            .O(N__44839),
            .I(\c0.n27_adj_4383 ));
    CascadeMux I__9042 (
            .O(N__44836),
            .I(\c0.n30_adj_4380_cascade_ ));
    InMux I__9041 (
            .O(N__44833),
            .I(N__44830));
    LocalMux I__9040 (
            .O(N__44830),
            .I(N__44827));
    Span4Mux_v I__9039 (
            .O(N__44827),
            .I(N__44824));
    Odrv4 I__9038 (
            .O(N__44824),
            .I(\c0.n28_adj_4381 ));
    InMux I__9037 (
            .O(N__44821),
            .I(N__44818));
    LocalMux I__9036 (
            .O(N__44818),
            .I(N__44814));
    InMux I__9035 (
            .O(N__44817),
            .I(N__44811));
    Odrv4 I__9034 (
            .O(N__44814),
            .I(\c0.n13000 ));
    LocalMux I__9033 (
            .O(N__44811),
            .I(\c0.n13000 ));
    CascadeMux I__9032 (
            .O(N__44806),
            .I(\c0.n10_adj_4286_cascade_ ));
    CascadeMux I__9031 (
            .O(N__44803),
            .I(N__44799));
    InMux I__9030 (
            .O(N__44802),
            .I(N__44794));
    InMux I__9029 (
            .O(N__44799),
            .I(N__44794));
    LocalMux I__9028 (
            .O(N__44794),
            .I(\c0.data_in_frame_28_2 ));
    CascadeMux I__9027 (
            .O(N__44791),
            .I(N__44787));
    InMux I__9026 (
            .O(N__44790),
            .I(N__44784));
    InMux I__9025 (
            .O(N__44787),
            .I(N__44781));
    LocalMux I__9024 (
            .O(N__44784),
            .I(N__44778));
    LocalMux I__9023 (
            .O(N__44781),
            .I(\c0.data_in_frame_29_0 ));
    Odrv4 I__9022 (
            .O(N__44778),
            .I(\c0.data_in_frame_29_0 ));
    InMux I__9021 (
            .O(N__44773),
            .I(N__44770));
    LocalMux I__9020 (
            .O(N__44770),
            .I(N__44767));
    Span4Mux_h I__9019 (
            .O(N__44767),
            .I(N__44764));
    Span4Mux_v I__9018 (
            .O(N__44764),
            .I(N__44761));
    Span4Mux_v I__9017 (
            .O(N__44761),
            .I(N__44758));
    Odrv4 I__9016 (
            .O(N__44758),
            .I(\c0.n17600 ));
    CascadeMux I__9015 (
            .O(N__44755),
            .I(\c0.n19_cascade_ ));
    InMux I__9014 (
            .O(N__44752),
            .I(N__44749));
    LocalMux I__9013 (
            .O(N__44749),
            .I(\c0.n23389 ));
    CascadeMux I__9012 (
            .O(N__44746),
            .I(\c0.n32_adj_4295_cascade_ ));
    InMux I__9011 (
            .O(N__44743),
            .I(N__44740));
    LocalMux I__9010 (
            .O(N__44740),
            .I(N__44737));
    Odrv4 I__9009 (
            .O(N__44737),
            .I(\c0.n23523 ));
    InMux I__9008 (
            .O(N__44734),
            .I(N__44731));
    LocalMux I__9007 (
            .O(N__44731),
            .I(\c0.n34 ));
    InMux I__9006 (
            .O(N__44728),
            .I(N__44725));
    LocalMux I__9005 (
            .O(N__44725),
            .I(N__44720));
    InMux I__9004 (
            .O(N__44724),
            .I(N__44715));
    InMux I__9003 (
            .O(N__44723),
            .I(N__44715));
    Odrv4 I__9002 (
            .O(N__44720),
            .I(\c0.n17790 ));
    LocalMux I__9001 (
            .O(N__44715),
            .I(\c0.n17790 ));
    InMux I__9000 (
            .O(N__44710),
            .I(N__44707));
    LocalMux I__8999 (
            .O(N__44707),
            .I(N__44704));
    Span4Mux_v I__8998 (
            .O(N__44704),
            .I(N__44699));
    CascadeMux I__8997 (
            .O(N__44703),
            .I(N__44692));
    InMux I__8996 (
            .O(N__44702),
            .I(N__44689));
    Span4Mux_v I__8995 (
            .O(N__44699),
            .I(N__44686));
    InMux I__8994 (
            .O(N__44698),
            .I(N__44683));
    InMux I__8993 (
            .O(N__44697),
            .I(N__44678));
    InMux I__8992 (
            .O(N__44696),
            .I(N__44678));
    InMux I__8991 (
            .O(N__44695),
            .I(N__44673));
    InMux I__8990 (
            .O(N__44692),
            .I(N__44673));
    LocalMux I__8989 (
            .O(N__44689),
            .I(data_in_frame_1_0));
    Odrv4 I__8988 (
            .O(N__44686),
            .I(data_in_frame_1_0));
    LocalMux I__8987 (
            .O(N__44683),
            .I(data_in_frame_1_0));
    LocalMux I__8986 (
            .O(N__44678),
            .I(data_in_frame_1_0));
    LocalMux I__8985 (
            .O(N__44673),
            .I(data_in_frame_1_0));
    CascadeMux I__8984 (
            .O(N__44662),
            .I(N__44656));
    InMux I__8983 (
            .O(N__44661),
            .I(N__44650));
    InMux I__8982 (
            .O(N__44660),
            .I(N__44647));
    InMux I__8981 (
            .O(N__44659),
            .I(N__44644));
    InMux I__8980 (
            .O(N__44656),
            .I(N__44637));
    InMux I__8979 (
            .O(N__44655),
            .I(N__44637));
    InMux I__8978 (
            .O(N__44654),
            .I(N__44637));
    InMux I__8977 (
            .O(N__44653),
            .I(N__44634));
    LocalMux I__8976 (
            .O(N__44650),
            .I(n23726));
    LocalMux I__8975 (
            .O(N__44647),
            .I(n23726));
    LocalMux I__8974 (
            .O(N__44644),
            .I(n23726));
    LocalMux I__8973 (
            .O(N__44637),
            .I(n23726));
    LocalMux I__8972 (
            .O(N__44634),
            .I(n23726));
    CascadeMux I__8971 (
            .O(N__44623),
            .I(N__44620));
    InMux I__8970 (
            .O(N__44620),
            .I(N__44615));
    InMux I__8969 (
            .O(N__44619),
            .I(N__44612));
    CascadeMux I__8968 (
            .O(N__44618),
            .I(N__44609));
    LocalMux I__8967 (
            .O(N__44615),
            .I(N__44603));
    LocalMux I__8966 (
            .O(N__44612),
            .I(N__44600));
    InMux I__8965 (
            .O(N__44609),
            .I(N__44597));
    InMux I__8964 (
            .O(N__44608),
            .I(N__44592));
    InMux I__8963 (
            .O(N__44607),
            .I(N__44592));
    InMux I__8962 (
            .O(N__44606),
            .I(N__44588));
    Span4Mux_v I__8961 (
            .O(N__44603),
            .I(N__44583));
    Span4Mux_v I__8960 (
            .O(N__44600),
            .I(N__44583));
    LocalMux I__8959 (
            .O(N__44597),
            .I(N__44578));
    LocalMux I__8958 (
            .O(N__44592),
            .I(N__44578));
    InMux I__8957 (
            .O(N__44591),
            .I(N__44575));
    LocalMux I__8956 (
            .O(N__44588),
            .I(N__44572));
    Span4Mux_h I__8955 (
            .O(N__44583),
            .I(N__44567));
    Span4Mux_v I__8954 (
            .O(N__44578),
            .I(N__44567));
    LocalMux I__8953 (
            .O(N__44575),
            .I(control_mode_0));
    Odrv4 I__8952 (
            .O(N__44572),
            .I(control_mode_0));
    Odrv4 I__8951 (
            .O(N__44567),
            .I(control_mode_0));
    CascadeMux I__8950 (
            .O(N__44560),
            .I(N__44556));
    InMux I__8949 (
            .O(N__44559),
            .I(N__44553));
    InMux I__8948 (
            .O(N__44556),
            .I(N__44550));
    LocalMux I__8947 (
            .O(N__44553),
            .I(\c0.data_in_frame_29_4 ));
    LocalMux I__8946 (
            .O(N__44550),
            .I(\c0.data_in_frame_29_4 ));
    CascadeMux I__8945 (
            .O(N__44545),
            .I(n4_cascade_));
    CascadeMux I__8944 (
            .O(N__44542),
            .I(N__44538));
    CascadeMux I__8943 (
            .O(N__44541),
            .I(N__44535));
    InMux I__8942 (
            .O(N__44538),
            .I(N__44529));
    InMux I__8941 (
            .O(N__44535),
            .I(N__44529));
    InMux I__8940 (
            .O(N__44534),
            .I(N__44526));
    LocalMux I__8939 (
            .O(N__44529),
            .I(N__44523));
    LocalMux I__8938 (
            .O(N__44526),
            .I(\c0.data_in_frame_4_6 ));
    Odrv12 I__8937 (
            .O(N__44523),
            .I(\c0.data_in_frame_4_6 ));
    InMux I__8936 (
            .O(N__44518),
            .I(N__44515));
    LocalMux I__8935 (
            .O(N__44515),
            .I(N__44512));
    Odrv4 I__8934 (
            .O(N__44512),
            .I(n4));
    CascadeMux I__8933 (
            .O(N__44509),
            .I(\c0.n21758_cascade_ ));
    CascadeMux I__8932 (
            .O(N__44506),
            .I(N__44502));
    CascadeMux I__8931 (
            .O(N__44505),
            .I(N__44499));
    InMux I__8930 (
            .O(N__44502),
            .I(N__44496));
    InMux I__8929 (
            .O(N__44499),
            .I(N__44493));
    LocalMux I__8928 (
            .O(N__44496),
            .I(N__44488));
    LocalMux I__8927 (
            .O(N__44493),
            .I(N__44485));
    InMux I__8926 (
            .O(N__44492),
            .I(N__44480));
    InMux I__8925 (
            .O(N__44491),
            .I(N__44480));
    Odrv4 I__8924 (
            .O(N__44488),
            .I(\c0.data_in_frame_2_4 ));
    Odrv12 I__8923 (
            .O(N__44485),
            .I(\c0.data_in_frame_2_4 ));
    LocalMux I__8922 (
            .O(N__44480),
            .I(\c0.data_in_frame_2_4 ));
    CascadeMux I__8921 (
            .O(N__44473),
            .I(N__44470));
    InMux I__8920 (
            .O(N__44470),
            .I(N__44465));
    InMux I__8919 (
            .O(N__44469),
            .I(N__44462));
    InMux I__8918 (
            .O(N__44468),
            .I(N__44459));
    LocalMux I__8917 (
            .O(N__44465),
            .I(N__44454));
    LocalMux I__8916 (
            .O(N__44462),
            .I(N__44454));
    LocalMux I__8915 (
            .O(N__44459),
            .I(\c0.data_in_frame_5_0 ));
    Odrv4 I__8914 (
            .O(N__44454),
            .I(\c0.data_in_frame_5_0 ));
    InMux I__8913 (
            .O(N__44449),
            .I(N__44445));
    CascadeMux I__8912 (
            .O(N__44448),
            .I(N__44440));
    LocalMux I__8911 (
            .O(N__44445),
            .I(N__44437));
    InMux I__8910 (
            .O(N__44444),
            .I(N__44432));
    InMux I__8909 (
            .O(N__44443),
            .I(N__44432));
    InMux I__8908 (
            .O(N__44440),
            .I(N__44429));
    Sp12to4 I__8907 (
            .O(N__44437),
            .I(N__44424));
    LocalMux I__8906 (
            .O(N__44432),
            .I(N__44424));
    LocalMux I__8905 (
            .O(N__44429),
            .I(\c0.data_in_frame_2_0 ));
    Odrv12 I__8904 (
            .O(N__44424),
            .I(\c0.data_in_frame_2_0 ));
    InMux I__8903 (
            .O(N__44419),
            .I(N__44416));
    LocalMux I__8902 (
            .O(N__44416),
            .I(N__44412));
    InMux I__8901 (
            .O(N__44415),
            .I(N__44409));
    Span4Mux_v I__8900 (
            .O(N__44412),
            .I(N__44406));
    LocalMux I__8899 (
            .O(N__44409),
            .I(data_in_frame_6_1));
    Odrv4 I__8898 (
            .O(N__44406),
            .I(data_in_frame_6_1));
    InMux I__8897 (
            .O(N__44401),
            .I(N__44395));
    InMux I__8896 (
            .O(N__44400),
            .I(N__44388));
    InMux I__8895 (
            .O(N__44399),
            .I(N__44388));
    InMux I__8894 (
            .O(N__44398),
            .I(N__44388));
    LocalMux I__8893 (
            .O(N__44395),
            .I(\c0.data_in_frame_4_7 ));
    LocalMux I__8892 (
            .O(N__44388),
            .I(\c0.data_in_frame_4_7 ));
    CascadeMux I__8891 (
            .O(N__44383),
            .I(N__44380));
    InMux I__8890 (
            .O(N__44380),
            .I(N__44375));
    InMux I__8889 (
            .O(N__44379),
            .I(N__44372));
    InMux I__8888 (
            .O(N__44378),
            .I(N__44369));
    LocalMux I__8887 (
            .O(N__44375),
            .I(\c0.data_in_frame_5_1 ));
    LocalMux I__8886 (
            .O(N__44372),
            .I(\c0.data_in_frame_5_1 ));
    LocalMux I__8885 (
            .O(N__44369),
            .I(\c0.data_in_frame_5_1 ));
    InMux I__8884 (
            .O(N__44362),
            .I(N__44356));
    InMux I__8883 (
            .O(N__44361),
            .I(N__44356));
    LocalMux I__8882 (
            .O(N__44356),
            .I(N__44352));
    InMux I__8881 (
            .O(N__44355),
            .I(N__44349));
    Odrv12 I__8880 (
            .O(N__44352),
            .I(\c0.n21992 ));
    LocalMux I__8879 (
            .O(N__44349),
            .I(\c0.n21992 ));
    CascadeMux I__8878 (
            .O(N__44344),
            .I(N__44340));
    CascadeMux I__8877 (
            .O(N__44343),
            .I(N__44337));
    InMux I__8876 (
            .O(N__44340),
            .I(N__44333));
    InMux I__8875 (
            .O(N__44337),
            .I(N__44330));
    InMux I__8874 (
            .O(N__44336),
            .I(N__44327));
    LocalMux I__8873 (
            .O(N__44333),
            .I(\c0.data_in_frame_2_2 ));
    LocalMux I__8872 (
            .O(N__44330),
            .I(\c0.data_in_frame_2_2 ));
    LocalMux I__8871 (
            .O(N__44327),
            .I(\c0.data_in_frame_2_2 ));
    CascadeMux I__8870 (
            .O(N__44320),
            .I(N__44317));
    InMux I__8869 (
            .O(N__44317),
            .I(N__44314));
    LocalMux I__8868 (
            .O(N__44314),
            .I(N__44311));
    Span4Mux_v I__8867 (
            .O(N__44311),
            .I(N__44305));
    InMux I__8866 (
            .O(N__44310),
            .I(N__44302));
    CascadeMux I__8865 (
            .O(N__44309),
            .I(N__44299));
    CascadeMux I__8864 (
            .O(N__44308),
            .I(N__44294));
    Span4Mux_v I__8863 (
            .O(N__44305),
            .I(N__44287));
    LocalMux I__8862 (
            .O(N__44302),
            .I(N__44287));
    InMux I__8861 (
            .O(N__44299),
            .I(N__44282));
    InMux I__8860 (
            .O(N__44298),
            .I(N__44282));
    InMux I__8859 (
            .O(N__44297),
            .I(N__44279));
    InMux I__8858 (
            .O(N__44294),
            .I(N__44272));
    InMux I__8857 (
            .O(N__44293),
            .I(N__44272));
    InMux I__8856 (
            .O(N__44292),
            .I(N__44272));
    Odrv4 I__8855 (
            .O(N__44287),
            .I(data_in_frame_1_7));
    LocalMux I__8854 (
            .O(N__44282),
            .I(data_in_frame_1_7));
    LocalMux I__8853 (
            .O(N__44279),
            .I(data_in_frame_1_7));
    LocalMux I__8852 (
            .O(N__44272),
            .I(data_in_frame_1_7));
    InMux I__8851 (
            .O(N__44263),
            .I(N__44260));
    LocalMux I__8850 (
            .O(N__44260),
            .I(\c0.n39_adj_4406 ));
    CascadeMux I__8849 (
            .O(N__44257),
            .I(N__44252));
    InMux I__8848 (
            .O(N__44256),
            .I(N__44248));
    InMux I__8847 (
            .O(N__44255),
            .I(N__44245));
    InMux I__8846 (
            .O(N__44252),
            .I(N__44242));
    InMux I__8845 (
            .O(N__44251),
            .I(N__44239));
    LocalMux I__8844 (
            .O(N__44248),
            .I(N__44236));
    LocalMux I__8843 (
            .O(N__44245),
            .I(data_in_frame_6_7));
    LocalMux I__8842 (
            .O(N__44242),
            .I(data_in_frame_6_7));
    LocalMux I__8841 (
            .O(N__44239),
            .I(data_in_frame_6_7));
    Odrv4 I__8840 (
            .O(N__44236),
            .I(data_in_frame_6_7));
    InMux I__8839 (
            .O(N__44227),
            .I(N__44224));
    LocalMux I__8838 (
            .O(N__44224),
            .I(\c0.n21882 ));
    InMux I__8837 (
            .O(N__44221),
            .I(N__44217));
    InMux I__8836 (
            .O(N__44220),
            .I(N__44214));
    LocalMux I__8835 (
            .O(N__44217),
            .I(N__44211));
    LocalMux I__8834 (
            .O(N__44214),
            .I(\c0.n21928 ));
    Odrv4 I__8833 (
            .O(N__44211),
            .I(\c0.n21928 ));
    CascadeMux I__8832 (
            .O(N__44206),
            .I(\c0.n14037_cascade_ ));
    InMux I__8831 (
            .O(N__44203),
            .I(N__44200));
    LocalMux I__8830 (
            .O(N__44200),
            .I(\c0.n6_adj_4369 ));
    InMux I__8829 (
            .O(N__44197),
            .I(N__44194));
    LocalMux I__8828 (
            .O(N__44194),
            .I(\c0.n5_adj_4368 ));
    InMux I__8827 (
            .O(N__44191),
            .I(N__44188));
    LocalMux I__8826 (
            .O(N__44188),
            .I(\c0.data_out_frame_29__7__N_1474 ));
    CascadeMux I__8825 (
            .O(N__44185),
            .I(N__44182));
    InMux I__8824 (
            .O(N__44182),
            .I(N__44178));
    InMux I__8823 (
            .O(N__44181),
            .I(N__44175));
    LocalMux I__8822 (
            .O(N__44178),
            .I(N__44172));
    LocalMux I__8821 (
            .O(N__44175),
            .I(data_in_frame_6_6));
    Odrv4 I__8820 (
            .O(N__44172),
            .I(data_in_frame_6_6));
    InMux I__8819 (
            .O(N__44167),
            .I(N__44162));
    InMux I__8818 (
            .O(N__44166),
            .I(N__44159));
    InMux I__8817 (
            .O(N__44165),
            .I(N__44156));
    LocalMux I__8816 (
            .O(N__44162),
            .I(N__44153));
    LocalMux I__8815 (
            .O(N__44159),
            .I(N__44150));
    LocalMux I__8814 (
            .O(N__44156),
            .I(N__44147));
    Span4Mux_h I__8813 (
            .O(N__44153),
            .I(N__44142));
    Span4Mux_v I__8812 (
            .O(N__44150),
            .I(N__44137));
    Span4Mux_h I__8811 (
            .O(N__44147),
            .I(N__44137));
    CascadeMux I__8810 (
            .O(N__44146),
            .I(N__44132));
    InMux I__8809 (
            .O(N__44145),
            .I(N__44129));
    Span4Mux_v I__8808 (
            .O(N__44142),
            .I(N__44126));
    Span4Mux_v I__8807 (
            .O(N__44137),
            .I(N__44123));
    InMux I__8806 (
            .O(N__44136),
            .I(N__44120));
    InMux I__8805 (
            .O(N__44135),
            .I(N__44115));
    InMux I__8804 (
            .O(N__44132),
            .I(N__44115));
    LocalMux I__8803 (
            .O(N__44129),
            .I(\c0.data_in_frame_0_2 ));
    Odrv4 I__8802 (
            .O(N__44126),
            .I(\c0.data_in_frame_0_2 ));
    Odrv4 I__8801 (
            .O(N__44123),
            .I(\c0.data_in_frame_0_2 ));
    LocalMux I__8800 (
            .O(N__44120),
            .I(\c0.data_in_frame_0_2 ));
    LocalMux I__8799 (
            .O(N__44115),
            .I(\c0.data_in_frame_0_2 ));
    CascadeMux I__8798 (
            .O(N__44104),
            .I(N__44100));
    InMux I__8797 (
            .O(N__44103),
            .I(N__44096));
    InMux I__8796 (
            .O(N__44100),
            .I(N__44093));
    InMux I__8795 (
            .O(N__44099),
            .I(N__44090));
    LocalMux I__8794 (
            .O(N__44096),
            .I(N__44087));
    LocalMux I__8793 (
            .O(N__44093),
            .I(\c0.data_in_frame_3_6 ));
    LocalMux I__8792 (
            .O(N__44090),
            .I(\c0.data_in_frame_3_6 ));
    Odrv4 I__8791 (
            .O(N__44087),
            .I(\c0.data_in_frame_3_6 ));
    InMux I__8790 (
            .O(N__44080),
            .I(N__44073));
    InMux I__8789 (
            .O(N__44079),
            .I(N__44073));
    InMux I__8788 (
            .O(N__44078),
            .I(N__44070));
    LocalMux I__8787 (
            .O(N__44073),
            .I(\c0.data_in_frame_4_1 ));
    LocalMux I__8786 (
            .O(N__44070),
            .I(\c0.data_in_frame_4_1 ));
    InMux I__8785 (
            .O(N__44065),
            .I(N__44061));
    InMux I__8784 (
            .O(N__44064),
            .I(N__44058));
    LocalMux I__8783 (
            .O(N__44061),
            .I(\c0.n22218 ));
    LocalMux I__8782 (
            .O(N__44058),
            .I(\c0.n22218 ));
    CascadeMux I__8781 (
            .O(N__44053),
            .I(\c0.n21928_cascade_ ));
    InMux I__8780 (
            .O(N__44050),
            .I(N__44045));
    CascadeMux I__8779 (
            .O(N__44049),
            .I(N__44042));
    CascadeMux I__8778 (
            .O(N__44048),
            .I(N__44039));
    LocalMux I__8777 (
            .O(N__44045),
            .I(N__44035));
    InMux I__8776 (
            .O(N__44042),
            .I(N__44032));
    InMux I__8775 (
            .O(N__44039),
            .I(N__44029));
    InMux I__8774 (
            .O(N__44038),
            .I(N__44026));
    Span4Mux_h I__8773 (
            .O(N__44035),
            .I(N__44021));
    LocalMux I__8772 (
            .O(N__44032),
            .I(N__44021));
    LocalMux I__8771 (
            .O(N__44029),
            .I(\c0.data_in_frame_2_3 ));
    LocalMux I__8770 (
            .O(N__44026),
            .I(\c0.data_in_frame_2_3 ));
    Odrv4 I__8769 (
            .O(N__44021),
            .I(\c0.data_in_frame_2_3 ));
    InMux I__8768 (
            .O(N__44014),
            .I(N__44009));
    InMux I__8767 (
            .O(N__44013),
            .I(N__44006));
    InMux I__8766 (
            .O(N__44012),
            .I(N__44003));
    LocalMux I__8765 (
            .O(N__44009),
            .I(N__44000));
    LocalMux I__8764 (
            .O(N__44006),
            .I(\c0.n21791 ));
    LocalMux I__8763 (
            .O(N__44003),
            .I(\c0.n21791 ));
    Odrv4 I__8762 (
            .O(N__44000),
            .I(\c0.n21791 ));
    CascadeMux I__8761 (
            .O(N__43993),
            .I(\c0.n21882_cascade_ ));
    InMux I__8760 (
            .O(N__43990),
            .I(N__43987));
    LocalMux I__8759 (
            .O(N__43987),
            .I(N__43984));
    Span4Mux_v I__8758 (
            .O(N__43984),
            .I(N__43981));
    Odrv4 I__8757 (
            .O(N__43981),
            .I(\c0.data_out_frame_0__7__N_2744 ));
    CascadeMux I__8756 (
            .O(N__43978),
            .I(\c0.data_out_frame_0__7__N_2744_cascade_ ));
    CascadeMux I__8755 (
            .O(N__43975),
            .I(\c0.n6_adj_4272_cascade_ ));
    CascadeMux I__8754 (
            .O(N__43972),
            .I(N__43967));
    InMux I__8753 (
            .O(N__43971),
            .I(N__43962));
    InMux I__8752 (
            .O(N__43970),
            .I(N__43962));
    InMux I__8751 (
            .O(N__43967),
            .I(N__43959));
    LocalMux I__8750 (
            .O(N__43962),
            .I(N__43956));
    LocalMux I__8749 (
            .O(N__43959),
            .I(\c0.data_in_frame_3_7 ));
    Odrv4 I__8748 (
            .O(N__43956),
            .I(\c0.data_in_frame_3_7 ));
    InMux I__8747 (
            .O(N__43951),
            .I(N__43948));
    LocalMux I__8746 (
            .O(N__43948),
            .I(\c0.n21803 ));
    InMux I__8745 (
            .O(N__43945),
            .I(N__43942));
    LocalMux I__8744 (
            .O(N__43942),
            .I(N__43939));
    Odrv12 I__8743 (
            .O(N__43939),
            .I(\c0.n18_adj_4370 ));
    InMux I__8742 (
            .O(N__43936),
            .I(N__43933));
    LocalMux I__8741 (
            .O(N__43933),
            .I(\c0.n22194 ));
    CascadeMux I__8740 (
            .O(N__43930),
            .I(\c0.n21803_cascade_ ));
    InMux I__8739 (
            .O(N__43927),
            .I(N__43924));
    LocalMux I__8738 (
            .O(N__43924),
            .I(\c0.n30_adj_4371 ));
    InMux I__8737 (
            .O(N__43921),
            .I(N__43915));
    InMux I__8736 (
            .O(N__43920),
            .I(N__43910));
    InMux I__8735 (
            .O(N__43919),
            .I(N__43910));
    InMux I__8734 (
            .O(N__43918),
            .I(N__43907));
    LocalMux I__8733 (
            .O(N__43915),
            .I(N__43904));
    LocalMux I__8732 (
            .O(N__43910),
            .I(N__43901));
    LocalMux I__8731 (
            .O(N__43907),
            .I(N__43892));
    Span4Mux_v I__8730 (
            .O(N__43904),
            .I(N__43892));
    Span4Mux_h I__8729 (
            .O(N__43901),
            .I(N__43892));
    InMux I__8728 (
            .O(N__43900),
            .I(N__43889));
    InMux I__8727 (
            .O(N__43899),
            .I(N__43886));
    Odrv4 I__8726 (
            .O(N__43892),
            .I(\c0.data_in_frame_0_1 ));
    LocalMux I__8725 (
            .O(N__43889),
            .I(\c0.data_in_frame_0_1 ));
    LocalMux I__8724 (
            .O(N__43886),
            .I(\c0.data_in_frame_0_1 ));
    CascadeMux I__8723 (
            .O(N__43879),
            .I(N__43875));
    InMux I__8722 (
            .O(N__43878),
            .I(N__43872));
    InMux I__8721 (
            .O(N__43875),
            .I(N__43865));
    LocalMux I__8720 (
            .O(N__43872),
            .I(N__43862));
    InMux I__8719 (
            .O(N__43871),
            .I(N__43859));
    InMux I__8718 (
            .O(N__43870),
            .I(N__43856));
    InMux I__8717 (
            .O(N__43869),
            .I(N__43851));
    InMux I__8716 (
            .O(N__43868),
            .I(N__43851));
    LocalMux I__8715 (
            .O(N__43865),
            .I(N__43848));
    Odrv12 I__8714 (
            .O(N__43862),
            .I(\c0.data_in_frame_0_0 ));
    LocalMux I__8713 (
            .O(N__43859),
            .I(\c0.data_in_frame_0_0 ));
    LocalMux I__8712 (
            .O(N__43856),
            .I(\c0.data_in_frame_0_0 ));
    LocalMux I__8711 (
            .O(N__43851),
            .I(\c0.data_in_frame_0_0 ));
    Odrv4 I__8710 (
            .O(N__43848),
            .I(\c0.data_in_frame_0_0 ));
    CascadeMux I__8709 (
            .O(N__43837),
            .I(\c0.n13376_cascade_ ));
    InMux I__8708 (
            .O(N__43834),
            .I(N__43830));
    InMux I__8707 (
            .O(N__43833),
            .I(N__43827));
    LocalMux I__8706 (
            .O(N__43830),
            .I(\c0.n13376 ));
    LocalMux I__8705 (
            .O(N__43827),
            .I(\c0.n13376 ));
    InMux I__8704 (
            .O(N__43822),
            .I(N__43819));
    LocalMux I__8703 (
            .O(N__43819),
            .I(N__43814));
    InMux I__8702 (
            .O(N__43818),
            .I(N__43811));
    InMux I__8701 (
            .O(N__43817),
            .I(N__43803));
    Span4Mux_v I__8700 (
            .O(N__43814),
            .I(N__43800));
    LocalMux I__8699 (
            .O(N__43811),
            .I(N__43797));
    InMux I__8698 (
            .O(N__43810),
            .I(N__43794));
    InMux I__8697 (
            .O(N__43809),
            .I(N__43791));
    InMux I__8696 (
            .O(N__43808),
            .I(N__43784));
    InMux I__8695 (
            .O(N__43807),
            .I(N__43784));
    InMux I__8694 (
            .O(N__43806),
            .I(N__43784));
    LocalMux I__8693 (
            .O(N__43803),
            .I(data_in_frame_1_6));
    Odrv4 I__8692 (
            .O(N__43800),
            .I(data_in_frame_1_6));
    Odrv12 I__8691 (
            .O(N__43797),
            .I(data_in_frame_1_6));
    LocalMux I__8690 (
            .O(N__43794),
            .I(data_in_frame_1_6));
    LocalMux I__8689 (
            .O(N__43791),
            .I(data_in_frame_1_6));
    LocalMux I__8688 (
            .O(N__43784),
            .I(data_in_frame_1_6));
    InMux I__8687 (
            .O(N__43771),
            .I(N__43767));
    InMux I__8686 (
            .O(N__43770),
            .I(N__43764));
    LocalMux I__8685 (
            .O(N__43767),
            .I(data_in_frame_6_2));
    LocalMux I__8684 (
            .O(N__43764),
            .I(data_in_frame_6_2));
    CascadeMux I__8683 (
            .O(N__43759),
            .I(\c0.n13386_cascade_ ));
    CascadeMux I__8682 (
            .O(N__43756),
            .I(N__43753));
    InMux I__8681 (
            .O(N__43753),
            .I(N__43748));
    InMux I__8680 (
            .O(N__43752),
            .I(N__43745));
    InMux I__8679 (
            .O(N__43751),
            .I(N__43742));
    LocalMux I__8678 (
            .O(N__43748),
            .I(\c0.data_in_frame_4_4 ));
    LocalMux I__8677 (
            .O(N__43745),
            .I(\c0.data_in_frame_4_4 ));
    LocalMux I__8676 (
            .O(N__43742),
            .I(\c0.data_in_frame_4_4 ));
    InMux I__8675 (
            .O(N__43735),
            .I(N__43732));
    LocalMux I__8674 (
            .O(N__43732),
            .I(\c0.n22261 ));
    CascadeMux I__8673 (
            .O(N__43729),
            .I(N__43725));
    InMux I__8672 (
            .O(N__43728),
            .I(N__43720));
    InMux I__8671 (
            .O(N__43725),
            .I(N__43715));
    InMux I__8670 (
            .O(N__43724),
            .I(N__43715));
    InMux I__8669 (
            .O(N__43723),
            .I(N__43712));
    LocalMux I__8668 (
            .O(N__43720),
            .I(\c0.data_in_frame_2_1 ));
    LocalMux I__8667 (
            .O(N__43715),
            .I(\c0.data_in_frame_2_1 ));
    LocalMux I__8666 (
            .O(N__43712),
            .I(\c0.data_in_frame_2_1 ));
    CascadeMux I__8665 (
            .O(N__43705),
            .I(\c0.n22261_cascade_ ));
    InMux I__8664 (
            .O(N__43702),
            .I(N__43699));
    LocalMux I__8663 (
            .O(N__43699),
            .I(\c0.n22320 ));
    InMux I__8662 (
            .O(N__43696),
            .I(N__43693));
    LocalMux I__8661 (
            .O(N__43693),
            .I(\c0.n28_adj_4372 ));
    InMux I__8660 (
            .O(N__43690),
            .I(N__43687));
    LocalMux I__8659 (
            .O(N__43687),
            .I(\c0.n22290 ));
    CascadeMux I__8658 (
            .O(N__43684),
            .I(N__43681));
    InMux I__8657 (
            .O(N__43681),
            .I(N__43678));
    LocalMux I__8656 (
            .O(N__43678),
            .I(\c0.n22258 ));
    CascadeMux I__8655 (
            .O(N__43675),
            .I(\c0.n22258_cascade_ ));
    InMux I__8654 (
            .O(N__43672),
            .I(N__43669));
    LocalMux I__8653 (
            .O(N__43669),
            .I(\c0.n29_adj_4374 ));
    CascadeMux I__8652 (
            .O(N__43666),
            .I(\c0.n27_adj_4377_cascade_ ));
    CascadeMux I__8651 (
            .O(N__43663),
            .I(\c0.n14072_cascade_ ));
    InMux I__8650 (
            .O(N__43660),
            .I(N__43657));
    LocalMux I__8649 (
            .O(N__43657),
            .I(\c0.n14072 ));
    CascadeMux I__8648 (
            .O(N__43654),
            .I(\c0.n6_adj_4385_cascade_ ));
    CascadeMux I__8647 (
            .O(N__43651),
            .I(\c0.n21902_cascade_ ));
    CascadeMux I__8646 (
            .O(N__43648),
            .I(N__43645));
    InMux I__8645 (
            .O(N__43645),
            .I(N__43639));
    InMux I__8644 (
            .O(N__43644),
            .I(N__43639));
    LocalMux I__8643 (
            .O(N__43639),
            .I(\c0.data_in_frame_3_0 ));
    InMux I__8642 (
            .O(N__43636),
            .I(N__43633));
    LocalMux I__8641 (
            .O(N__43633),
            .I(\c0.n21902 ));
    CascadeMux I__8640 (
            .O(N__43630),
            .I(N__43626));
    CascadeMux I__8639 (
            .O(N__43629),
            .I(N__43623));
    InMux I__8638 (
            .O(N__43626),
            .I(N__43620));
    InMux I__8637 (
            .O(N__43623),
            .I(N__43617));
    LocalMux I__8636 (
            .O(N__43620),
            .I(\c0.data_in_frame_5_2 ));
    LocalMux I__8635 (
            .O(N__43617),
            .I(\c0.data_in_frame_5_2 ));
    CascadeMux I__8634 (
            .O(N__43612),
            .I(\c0.n21879_cascade_ ));
    CascadeMux I__8633 (
            .O(N__43609),
            .I(N__43606));
    InMux I__8632 (
            .O(N__43606),
            .I(N__43599));
    InMux I__8631 (
            .O(N__43605),
            .I(N__43599));
    InMux I__8630 (
            .O(N__43604),
            .I(N__43596));
    LocalMux I__8629 (
            .O(N__43599),
            .I(\c0.data_in_frame_3_4 ));
    LocalMux I__8628 (
            .O(N__43596),
            .I(\c0.data_in_frame_3_4 ));
    InMux I__8627 (
            .O(N__43591),
            .I(N__43588));
    LocalMux I__8626 (
            .O(N__43588),
            .I(N__43585));
    Odrv4 I__8625 (
            .O(N__43585),
            .I(\c0.n21957 ));
    CascadeMux I__8624 (
            .O(N__43582),
            .I(\c0.n21957_cascade_ ));
    InMux I__8623 (
            .O(N__43579),
            .I(N__43576));
    LocalMux I__8622 (
            .O(N__43576),
            .I(\c0.n22287 ));
    InMux I__8621 (
            .O(N__43573),
            .I(N__43564));
    InMux I__8620 (
            .O(N__43572),
            .I(N__43564));
    InMux I__8619 (
            .O(N__43571),
            .I(N__43564));
    LocalMux I__8618 (
            .O(N__43564),
            .I(\c0.data_in_frame_3_3 ));
    CascadeMux I__8617 (
            .O(N__43561),
            .I(N__43558));
    InMux I__8616 (
            .O(N__43558),
            .I(N__43552));
    InMux I__8615 (
            .O(N__43557),
            .I(N__43552));
    LocalMux I__8614 (
            .O(N__43552),
            .I(\c0.data_in_frame_5_4 ));
    InMux I__8613 (
            .O(N__43549),
            .I(N__43546));
    LocalMux I__8612 (
            .O(N__43546),
            .I(N__43543));
    Odrv4 I__8611 (
            .O(N__43543),
            .I(\c0.n23838 ));
    InMux I__8610 (
            .O(N__43540),
            .I(N__43536));
    InMux I__8609 (
            .O(N__43539),
            .I(N__43533));
    LocalMux I__8608 (
            .O(N__43536),
            .I(N__43526));
    LocalMux I__8607 (
            .O(N__43533),
            .I(N__43526));
    InMux I__8606 (
            .O(N__43532),
            .I(N__43523));
    InMux I__8605 (
            .O(N__43531),
            .I(N__43520));
    Span4Mux_h I__8604 (
            .O(N__43526),
            .I(N__43517));
    LocalMux I__8603 (
            .O(N__43523),
            .I(\c0.FRAME_MATCHER_state_28 ));
    LocalMux I__8602 (
            .O(N__43520),
            .I(\c0.FRAME_MATCHER_state_28 ));
    Odrv4 I__8601 (
            .O(N__43517),
            .I(\c0.FRAME_MATCHER_state_28 ));
    SRMux I__8600 (
            .O(N__43510),
            .I(N__43507));
    LocalMux I__8599 (
            .O(N__43507),
            .I(\c0.n21378 ));
    InMux I__8598 (
            .O(N__43504),
            .I(N__43499));
    InMux I__8597 (
            .O(N__43503),
            .I(N__43496));
    CascadeMux I__8596 (
            .O(N__43502),
            .I(N__43493));
    LocalMux I__8595 (
            .O(N__43499),
            .I(N__43488));
    LocalMux I__8594 (
            .O(N__43496),
            .I(N__43488));
    InMux I__8593 (
            .O(N__43493),
            .I(N__43484));
    Span4Mux_v I__8592 (
            .O(N__43488),
            .I(N__43481));
    InMux I__8591 (
            .O(N__43487),
            .I(N__43478));
    LocalMux I__8590 (
            .O(N__43484),
            .I(N__43475));
    Span4Mux_h I__8589 (
            .O(N__43481),
            .I(N__43472));
    LocalMux I__8588 (
            .O(N__43478),
            .I(\c0.FRAME_MATCHER_state_31 ));
    Odrv4 I__8587 (
            .O(N__43475),
            .I(\c0.FRAME_MATCHER_state_31 ));
    Odrv4 I__8586 (
            .O(N__43472),
            .I(\c0.FRAME_MATCHER_state_31 ));
    SRMux I__8585 (
            .O(N__43465),
            .I(N__43462));
    LocalMux I__8584 (
            .O(N__43462),
            .I(N__43459));
    Odrv4 I__8583 (
            .O(N__43459),
            .I(\c0.n21332 ));
    CascadeMux I__8582 (
            .O(N__43456),
            .I(N__43452));
    InMux I__8581 (
            .O(N__43455),
            .I(N__43448));
    InMux I__8580 (
            .O(N__43452),
            .I(N__43445));
    InMux I__8579 (
            .O(N__43451),
            .I(N__43441));
    LocalMux I__8578 (
            .O(N__43448),
            .I(N__43436));
    LocalMux I__8577 (
            .O(N__43445),
            .I(N__43436));
    InMux I__8576 (
            .O(N__43444),
            .I(N__43433));
    LocalMux I__8575 (
            .O(N__43441),
            .I(N__43430));
    Span4Mux_h I__8574 (
            .O(N__43436),
            .I(N__43427));
    LocalMux I__8573 (
            .O(N__43433),
            .I(\c0.FRAME_MATCHER_state_13 ));
    Odrv12 I__8572 (
            .O(N__43430),
            .I(\c0.FRAME_MATCHER_state_13 ));
    Odrv4 I__8571 (
            .O(N__43427),
            .I(\c0.FRAME_MATCHER_state_13 ));
    SRMux I__8570 (
            .O(N__43420),
            .I(N__43417));
    LocalMux I__8569 (
            .O(N__43417),
            .I(N__43414));
    Odrv4 I__8568 (
            .O(N__43414),
            .I(\c0.n21354 ));
    InMux I__8567 (
            .O(N__43411),
            .I(N__43407));
    CascadeMux I__8566 (
            .O(N__43410),
            .I(N__43404));
    LocalMux I__8565 (
            .O(N__43407),
            .I(N__43401));
    InMux I__8564 (
            .O(N__43404),
            .I(N__43398));
    Span4Mux_h I__8563 (
            .O(N__43401),
            .I(N__43395));
    LocalMux I__8562 (
            .O(N__43398),
            .I(N__43388));
    Span4Mux_v I__8561 (
            .O(N__43395),
            .I(N__43388));
    InMux I__8560 (
            .O(N__43394),
            .I(N__43385));
    InMux I__8559 (
            .O(N__43393),
            .I(N__43382));
    Span4Mux_h I__8558 (
            .O(N__43388),
            .I(N__43379));
    LocalMux I__8557 (
            .O(N__43385),
            .I(\c0.FRAME_MATCHER_state_15 ));
    LocalMux I__8556 (
            .O(N__43382),
            .I(\c0.FRAME_MATCHER_state_15 ));
    Odrv4 I__8555 (
            .O(N__43379),
            .I(\c0.FRAME_MATCHER_state_15 ));
    SRMux I__8554 (
            .O(N__43372),
            .I(N__43369));
    LocalMux I__8553 (
            .O(N__43369),
            .I(N__43366));
    Odrv4 I__8552 (
            .O(N__43366),
            .I(\c0.n21358 ));
    InMux I__8551 (
            .O(N__43363),
            .I(N__43358));
    InMux I__8550 (
            .O(N__43362),
            .I(N__43353));
    InMux I__8549 (
            .O(N__43361),
            .I(N__43353));
    LocalMux I__8548 (
            .O(N__43358),
            .I(N__43350));
    LocalMux I__8547 (
            .O(N__43353),
            .I(\c0.n21734 ));
    Odrv4 I__8546 (
            .O(N__43350),
            .I(\c0.n21734 ));
    InMux I__8545 (
            .O(N__43345),
            .I(N__43333));
    InMux I__8544 (
            .O(N__43344),
            .I(N__43333));
    InMux I__8543 (
            .O(N__43343),
            .I(N__43333));
    InMux I__8542 (
            .O(N__43342),
            .I(N__43330));
    InMux I__8541 (
            .O(N__43341),
            .I(N__43325));
    InMux I__8540 (
            .O(N__43340),
            .I(N__43325));
    LocalMux I__8539 (
            .O(N__43333),
            .I(N__43322));
    LocalMux I__8538 (
            .O(N__43330),
            .I(N__43319));
    LocalMux I__8537 (
            .O(N__43325),
            .I(N__43314));
    Span4Mux_h I__8536 (
            .O(N__43322),
            .I(N__43314));
    Span4Mux_h I__8535 (
            .O(N__43319),
            .I(N__43311));
    Odrv4 I__8534 (
            .O(N__43314),
            .I(\c0.n13021 ));
    Odrv4 I__8533 (
            .O(N__43311),
            .I(\c0.n13021 ));
    CascadeMux I__8532 (
            .O(N__43306),
            .I(N__43303));
    InMux I__8531 (
            .O(N__43303),
            .I(N__43300));
    LocalMux I__8530 (
            .O(N__43300),
            .I(N__43297));
    Span4Mux_h I__8529 (
            .O(N__43297),
            .I(N__43294));
    Odrv4 I__8528 (
            .O(N__43294),
            .I(\c0.n23965 ));
    InMux I__8527 (
            .O(N__43291),
            .I(N__43287));
    InMux I__8526 (
            .O(N__43290),
            .I(N__43284));
    LocalMux I__8525 (
            .O(N__43287),
            .I(\c0.n22575 ));
    LocalMux I__8524 (
            .O(N__43284),
            .I(\c0.n22575 ));
    InMux I__8523 (
            .O(N__43279),
            .I(N__43276));
    LocalMux I__8522 (
            .O(N__43276),
            .I(\c0.n45_adj_4389 ));
    CascadeMux I__8521 (
            .O(N__43273),
            .I(N__43270));
    InMux I__8520 (
            .O(N__43270),
            .I(N__43251));
    InMux I__8519 (
            .O(N__43269),
            .I(N__43251));
    InMux I__8518 (
            .O(N__43268),
            .I(N__43251));
    InMux I__8517 (
            .O(N__43267),
            .I(N__43246));
    InMux I__8516 (
            .O(N__43266),
            .I(N__43246));
    CascadeMux I__8515 (
            .O(N__43265),
            .I(N__43240));
    InMux I__8514 (
            .O(N__43264),
            .I(N__43236));
    InMux I__8513 (
            .O(N__43263),
            .I(N__43233));
    InMux I__8512 (
            .O(N__43262),
            .I(N__43230));
    InMux I__8511 (
            .O(N__43261),
            .I(N__43227));
    InMux I__8510 (
            .O(N__43260),
            .I(N__43220));
    InMux I__8509 (
            .O(N__43259),
            .I(N__43220));
    InMux I__8508 (
            .O(N__43258),
            .I(N__43220));
    LocalMux I__8507 (
            .O(N__43251),
            .I(N__43210));
    LocalMux I__8506 (
            .O(N__43246),
            .I(N__43210));
    InMux I__8505 (
            .O(N__43245),
            .I(N__43199));
    InMux I__8504 (
            .O(N__43244),
            .I(N__43199));
    InMux I__8503 (
            .O(N__43243),
            .I(N__43199));
    InMux I__8502 (
            .O(N__43240),
            .I(N__43199));
    InMux I__8501 (
            .O(N__43239),
            .I(N__43199));
    LocalMux I__8500 (
            .O(N__43236),
            .I(N__43194));
    LocalMux I__8499 (
            .O(N__43233),
            .I(N__43194));
    LocalMux I__8498 (
            .O(N__43230),
            .I(N__43185));
    LocalMux I__8497 (
            .O(N__43227),
            .I(N__43185));
    LocalMux I__8496 (
            .O(N__43220),
            .I(N__43185));
    InMux I__8495 (
            .O(N__43219),
            .I(N__43182));
    InMux I__8494 (
            .O(N__43218),
            .I(N__43179));
    InMux I__8493 (
            .O(N__43217),
            .I(N__43176));
    InMux I__8492 (
            .O(N__43216),
            .I(N__43172));
    InMux I__8491 (
            .O(N__43215),
            .I(N__43166));
    Span4Mux_v I__8490 (
            .O(N__43210),
            .I(N__43161));
    LocalMux I__8489 (
            .O(N__43199),
            .I(N__43161));
    Span4Mux_v I__8488 (
            .O(N__43194),
            .I(N__43158));
    InMux I__8487 (
            .O(N__43193),
            .I(N__43151));
    InMux I__8486 (
            .O(N__43192),
            .I(N__43148));
    Span4Mux_v I__8485 (
            .O(N__43185),
            .I(N__43139));
    LocalMux I__8484 (
            .O(N__43182),
            .I(N__43139));
    LocalMux I__8483 (
            .O(N__43179),
            .I(N__43139));
    LocalMux I__8482 (
            .O(N__43176),
            .I(N__43139));
    InMux I__8481 (
            .O(N__43175),
            .I(N__43136));
    LocalMux I__8480 (
            .O(N__43172),
            .I(N__43133));
    InMux I__8479 (
            .O(N__43171),
            .I(N__43130));
    InMux I__8478 (
            .O(N__43170),
            .I(N__43125));
    InMux I__8477 (
            .O(N__43169),
            .I(N__43125));
    LocalMux I__8476 (
            .O(N__43166),
            .I(N__43120));
    Span4Mux_h I__8475 (
            .O(N__43161),
            .I(N__43120));
    Sp12to4 I__8474 (
            .O(N__43158),
            .I(N__43117));
    InMux I__8473 (
            .O(N__43157),
            .I(N__43112));
    InMux I__8472 (
            .O(N__43156),
            .I(N__43112));
    InMux I__8471 (
            .O(N__43155),
            .I(N__43106));
    InMux I__8470 (
            .O(N__43154),
            .I(N__43103));
    LocalMux I__8469 (
            .O(N__43151),
            .I(N__43096));
    LocalMux I__8468 (
            .O(N__43148),
            .I(N__43096));
    Span4Mux_h I__8467 (
            .O(N__43139),
            .I(N__43096));
    LocalMux I__8466 (
            .O(N__43136),
            .I(N__43091));
    Span4Mux_v I__8465 (
            .O(N__43133),
            .I(N__43091));
    LocalMux I__8464 (
            .O(N__43130),
            .I(N__43080));
    LocalMux I__8463 (
            .O(N__43125),
            .I(N__43080));
    Sp12to4 I__8462 (
            .O(N__43120),
            .I(N__43080));
    Span12Mux_h I__8461 (
            .O(N__43117),
            .I(N__43080));
    LocalMux I__8460 (
            .O(N__43112),
            .I(N__43080));
    InMux I__8459 (
            .O(N__43111),
            .I(N__43072));
    InMux I__8458 (
            .O(N__43110),
            .I(N__43072));
    InMux I__8457 (
            .O(N__43109),
            .I(N__43072));
    LocalMux I__8456 (
            .O(N__43106),
            .I(N__43067));
    LocalMux I__8455 (
            .O(N__43103),
            .I(N__43067));
    Span4Mux_v I__8454 (
            .O(N__43096),
            .I(N__43064));
    Sp12to4 I__8453 (
            .O(N__43091),
            .I(N__43059));
    Span12Mux_v I__8452 (
            .O(N__43080),
            .I(N__43059));
    InMux I__8451 (
            .O(N__43079),
            .I(N__43056));
    LocalMux I__8450 (
            .O(N__43072),
            .I(rx_data_ready));
    Odrv12 I__8449 (
            .O(N__43067),
            .I(rx_data_ready));
    Odrv4 I__8448 (
            .O(N__43064),
            .I(rx_data_ready));
    Odrv12 I__8447 (
            .O(N__43059),
            .I(rx_data_ready));
    LocalMux I__8446 (
            .O(N__43056),
            .I(rx_data_ready));
    InMux I__8445 (
            .O(N__43045),
            .I(N__43038));
    InMux I__8444 (
            .O(N__43044),
            .I(N__43038));
    InMux I__8443 (
            .O(N__43043),
            .I(N__43035));
    LocalMux I__8442 (
            .O(N__43038),
            .I(N__43032));
    LocalMux I__8441 (
            .O(N__43035),
            .I(N__43028));
    Span4Mux_h I__8440 (
            .O(N__43032),
            .I(N__43025));
    InMux I__8439 (
            .O(N__43031),
            .I(N__43022));
    Span4Mux_v I__8438 (
            .O(N__43028),
            .I(N__43019));
    Span4Mux_h I__8437 (
            .O(N__43025),
            .I(N__43016));
    LocalMux I__8436 (
            .O(N__43022),
            .I(data_in_3_1));
    Odrv4 I__8435 (
            .O(N__43019),
            .I(data_in_3_1));
    Odrv4 I__8434 (
            .O(N__43016),
            .I(data_in_3_1));
    InMux I__8433 (
            .O(N__43009),
            .I(N__43004));
    InMux I__8432 (
            .O(N__43008),
            .I(N__43001));
    InMux I__8431 (
            .O(N__43007),
            .I(N__42998));
    LocalMux I__8430 (
            .O(N__43004),
            .I(N__42995));
    LocalMux I__8429 (
            .O(N__43001),
            .I(N__42990));
    LocalMux I__8428 (
            .O(N__42998),
            .I(N__42990));
    Odrv4 I__8427 (
            .O(N__42995),
            .I(\c0.n1 ));
    Odrv12 I__8426 (
            .O(N__42990),
            .I(\c0.n1 ));
    InMux I__8425 (
            .O(N__42985),
            .I(N__42982));
    LocalMux I__8424 (
            .O(N__42982),
            .I(N__42979));
    Span4Mux_v I__8423 (
            .O(N__42979),
            .I(N__42975));
    InMux I__8422 (
            .O(N__42978),
            .I(N__42972));
    Span4Mux_h I__8421 (
            .O(N__42975),
            .I(N__42966));
    LocalMux I__8420 (
            .O(N__42972),
            .I(N__42966));
    InMux I__8419 (
            .O(N__42971),
            .I(N__42963));
    Sp12to4 I__8418 (
            .O(N__42966),
            .I(N__42958));
    LocalMux I__8417 (
            .O(N__42963),
            .I(N__42958));
    Odrv12 I__8416 (
            .O(N__42958),
            .I(\c0.n19783 ));
    InMux I__8415 (
            .O(N__42955),
            .I(N__42951));
    InMux I__8414 (
            .O(N__42954),
            .I(N__42948));
    LocalMux I__8413 (
            .O(N__42951),
            .I(N__42943));
    LocalMux I__8412 (
            .O(N__42948),
            .I(N__42943));
    Span4Mux_h I__8411 (
            .O(N__42943),
            .I(N__42940));
    Odrv4 I__8410 (
            .O(N__42940),
            .I(\c0.n937 ));
    InMux I__8409 (
            .O(N__42937),
            .I(N__42932));
    CascadeMux I__8408 (
            .O(N__42936),
            .I(N__42929));
    InMux I__8407 (
            .O(N__42935),
            .I(N__42925));
    LocalMux I__8406 (
            .O(N__42932),
            .I(N__42922));
    InMux I__8405 (
            .O(N__42929),
            .I(N__42919));
    InMux I__8404 (
            .O(N__42928),
            .I(N__42916));
    LocalMux I__8403 (
            .O(N__42925),
            .I(N__42913));
    Span4Mux_h I__8402 (
            .O(N__42922),
            .I(N__42910));
    LocalMux I__8401 (
            .O(N__42919),
            .I(N__42907));
    LocalMux I__8400 (
            .O(N__42916),
            .I(\c0.FRAME_MATCHER_state_12 ));
    Odrv4 I__8399 (
            .O(N__42913),
            .I(\c0.FRAME_MATCHER_state_12 ));
    Odrv4 I__8398 (
            .O(N__42910),
            .I(\c0.FRAME_MATCHER_state_12 ));
    Odrv12 I__8397 (
            .O(N__42907),
            .I(\c0.FRAME_MATCHER_state_12 ));
    SRMux I__8396 (
            .O(N__42898),
            .I(N__42895));
    LocalMux I__8395 (
            .O(N__42895),
            .I(N__42892));
    Span4Mux_h I__8394 (
            .O(N__42892),
            .I(N__42889));
    Odrv4 I__8393 (
            .O(N__42889),
            .I(\c0.n21352 ));
    CascadeMux I__8392 (
            .O(N__42886),
            .I(N__42881));
    InMux I__8391 (
            .O(N__42885),
            .I(N__42877));
    InMux I__8390 (
            .O(N__42884),
            .I(N__42874));
    InMux I__8389 (
            .O(N__42881),
            .I(N__42871));
    InMux I__8388 (
            .O(N__42880),
            .I(N__42867));
    LocalMux I__8387 (
            .O(N__42877),
            .I(N__42864));
    LocalMux I__8386 (
            .O(N__42874),
            .I(N__42859));
    LocalMux I__8385 (
            .O(N__42871),
            .I(N__42859));
    InMux I__8384 (
            .O(N__42870),
            .I(N__42856));
    LocalMux I__8383 (
            .O(N__42867),
            .I(N__42853));
    Span4Mux_v I__8382 (
            .O(N__42864),
            .I(N__42850));
    Span4Mux_v I__8381 (
            .O(N__42859),
            .I(N__42847));
    LocalMux I__8380 (
            .O(N__42856),
            .I(N__42844));
    Odrv12 I__8379 (
            .O(N__42853),
            .I(\c0.n20_adj_4327 ));
    Odrv4 I__8378 (
            .O(N__42850),
            .I(\c0.n20_adj_4327 ));
    Odrv4 I__8377 (
            .O(N__42847),
            .I(\c0.n20_adj_4327 ));
    Odrv12 I__8376 (
            .O(N__42844),
            .I(\c0.n20_adj_4327 ));
    InMux I__8375 (
            .O(N__42835),
            .I(N__42830));
    InMux I__8374 (
            .O(N__42834),
            .I(N__42827));
    InMux I__8373 (
            .O(N__42833),
            .I(N__42822));
    LocalMux I__8372 (
            .O(N__42830),
            .I(N__42819));
    LocalMux I__8371 (
            .O(N__42827),
            .I(N__42816));
    InMux I__8370 (
            .O(N__42826),
            .I(N__42813));
    InMux I__8369 (
            .O(N__42825),
            .I(N__42810));
    LocalMux I__8368 (
            .O(N__42822),
            .I(\c0.n12992 ));
    Odrv4 I__8367 (
            .O(N__42819),
            .I(\c0.n12992 ));
    Odrv12 I__8366 (
            .O(N__42816),
            .I(\c0.n12992 ));
    LocalMux I__8365 (
            .O(N__42813),
            .I(\c0.n12992 ));
    LocalMux I__8364 (
            .O(N__42810),
            .I(\c0.n12992 ));
    InMux I__8363 (
            .O(N__42799),
            .I(N__42782));
    InMux I__8362 (
            .O(N__42798),
            .I(N__42779));
    InMux I__8361 (
            .O(N__42797),
            .I(N__42770));
    InMux I__8360 (
            .O(N__42796),
            .I(N__42770));
    InMux I__8359 (
            .O(N__42795),
            .I(N__42770));
    InMux I__8358 (
            .O(N__42794),
            .I(N__42770));
    InMux I__8357 (
            .O(N__42793),
            .I(N__42755));
    InMux I__8356 (
            .O(N__42792),
            .I(N__42755));
    InMux I__8355 (
            .O(N__42791),
            .I(N__42755));
    InMux I__8354 (
            .O(N__42790),
            .I(N__42755));
    InMux I__8353 (
            .O(N__42789),
            .I(N__42755));
    InMux I__8352 (
            .O(N__42788),
            .I(N__42752));
    InMux I__8351 (
            .O(N__42787),
            .I(N__42745));
    InMux I__8350 (
            .O(N__42786),
            .I(N__42745));
    InMux I__8349 (
            .O(N__42785),
            .I(N__42745));
    LocalMux I__8348 (
            .O(N__42782),
            .I(N__42740));
    LocalMux I__8347 (
            .O(N__42779),
            .I(N__42737));
    LocalMux I__8346 (
            .O(N__42770),
            .I(N__42734));
    InMux I__8345 (
            .O(N__42769),
            .I(N__42729));
    InMux I__8344 (
            .O(N__42768),
            .I(N__42729));
    InMux I__8343 (
            .O(N__42767),
            .I(N__42724));
    InMux I__8342 (
            .O(N__42766),
            .I(N__42724));
    LocalMux I__8341 (
            .O(N__42755),
            .I(N__42721));
    LocalMux I__8340 (
            .O(N__42752),
            .I(N__42716));
    LocalMux I__8339 (
            .O(N__42745),
            .I(N__42716));
    InMux I__8338 (
            .O(N__42744),
            .I(N__42711));
    InMux I__8337 (
            .O(N__42743),
            .I(N__42711));
    Span4Mux_v I__8336 (
            .O(N__42740),
            .I(N__42700));
    Span4Mux_h I__8335 (
            .O(N__42737),
            .I(N__42693));
    Span4Mux_h I__8334 (
            .O(N__42734),
            .I(N__42693));
    LocalMux I__8333 (
            .O(N__42729),
            .I(N__42693));
    LocalMux I__8332 (
            .O(N__42724),
            .I(N__42690));
    Span4Mux_h I__8331 (
            .O(N__42721),
            .I(N__42687));
    Span4Mux_v I__8330 (
            .O(N__42716),
            .I(N__42682));
    LocalMux I__8329 (
            .O(N__42711),
            .I(N__42682));
    InMux I__8328 (
            .O(N__42710),
            .I(N__42675));
    InMux I__8327 (
            .O(N__42709),
            .I(N__42675));
    InMux I__8326 (
            .O(N__42708),
            .I(N__42675));
    InMux I__8325 (
            .O(N__42707),
            .I(N__42664));
    InMux I__8324 (
            .O(N__42706),
            .I(N__42664));
    InMux I__8323 (
            .O(N__42705),
            .I(N__42664));
    InMux I__8322 (
            .O(N__42704),
            .I(N__42664));
    InMux I__8321 (
            .O(N__42703),
            .I(N__42664));
    Odrv4 I__8320 (
            .O(N__42700),
            .I(\c0.n9668 ));
    Odrv4 I__8319 (
            .O(N__42693),
            .I(\c0.n9668 ));
    Odrv4 I__8318 (
            .O(N__42690),
            .I(\c0.n9668 ));
    Odrv4 I__8317 (
            .O(N__42687),
            .I(\c0.n9668 ));
    Odrv4 I__8316 (
            .O(N__42682),
            .I(\c0.n9668 ));
    LocalMux I__8315 (
            .O(N__42675),
            .I(\c0.n9668 ));
    LocalMux I__8314 (
            .O(N__42664),
            .I(\c0.n9668 ));
    InMux I__8313 (
            .O(N__42649),
            .I(N__42646));
    LocalMux I__8312 (
            .O(N__42646),
            .I(\c0.n7_adj_4356 ));
    InMux I__8311 (
            .O(N__42643),
            .I(N__42640));
    LocalMux I__8310 (
            .O(N__42640),
            .I(N__42635));
    InMux I__8309 (
            .O(N__42639),
            .I(N__42632));
    InMux I__8308 (
            .O(N__42638),
            .I(N__42629));
    Span4Mux_v I__8307 (
            .O(N__42635),
            .I(N__42624));
    LocalMux I__8306 (
            .O(N__42632),
            .I(N__42624));
    LocalMux I__8305 (
            .O(N__42629),
            .I(N__42621));
    Odrv4 I__8304 (
            .O(N__42624),
            .I(\c0.n12876 ));
    Odrv4 I__8303 (
            .O(N__42621),
            .I(\c0.n12876 ));
    CascadeMux I__8302 (
            .O(N__42616),
            .I(N__42612));
    InMux I__8301 (
            .O(N__42615),
            .I(N__42605));
    InMux I__8300 (
            .O(N__42612),
            .I(N__42605));
    InMux I__8299 (
            .O(N__42611),
            .I(N__42602));
    InMux I__8298 (
            .O(N__42610),
            .I(N__42599));
    LocalMux I__8297 (
            .O(N__42605),
            .I(N__42594));
    LocalMux I__8296 (
            .O(N__42602),
            .I(N__42594));
    LocalMux I__8295 (
            .O(N__42599),
            .I(\c0.n21022 ));
    Odrv4 I__8294 (
            .O(N__42594),
            .I(\c0.n21022 ));
    InMux I__8293 (
            .O(N__42589),
            .I(N__42586));
    LocalMux I__8292 (
            .O(N__42586),
            .I(N__42581));
    InMux I__8291 (
            .O(N__42585),
            .I(N__42578));
    InMux I__8290 (
            .O(N__42584),
            .I(N__42575));
    Odrv4 I__8289 (
            .O(N__42581),
            .I(\c0.n12991 ));
    LocalMux I__8288 (
            .O(N__42578),
            .I(\c0.n12991 ));
    LocalMux I__8287 (
            .O(N__42575),
            .I(\c0.n12991 ));
    InMux I__8286 (
            .O(N__42568),
            .I(N__42564));
    CascadeMux I__8285 (
            .O(N__42567),
            .I(N__42561));
    LocalMux I__8284 (
            .O(N__42564),
            .I(N__42558));
    InMux I__8283 (
            .O(N__42561),
            .I(N__42555));
    Odrv4 I__8282 (
            .O(N__42558),
            .I(\c0.n5024 ));
    LocalMux I__8281 (
            .O(N__42555),
            .I(\c0.n5024 ));
    CascadeMux I__8280 (
            .O(N__42550),
            .I(\c0.n5_adj_4342_cascade_ ));
    InMux I__8279 (
            .O(N__42547),
            .I(N__42542));
    InMux I__8278 (
            .O(N__42546),
            .I(N__42539));
    CascadeMux I__8277 (
            .O(N__42545),
            .I(N__42535));
    LocalMux I__8276 (
            .O(N__42542),
            .I(N__42532));
    LocalMux I__8275 (
            .O(N__42539),
            .I(N__42529));
    InMux I__8274 (
            .O(N__42538),
            .I(N__42524));
    InMux I__8273 (
            .O(N__42535),
            .I(N__42524));
    Span4Mux_v I__8272 (
            .O(N__42532),
            .I(N__42521));
    Span4Mux_v I__8271 (
            .O(N__42529),
            .I(N__42518));
    LocalMux I__8270 (
            .O(N__42524),
            .I(N__42515));
    Odrv4 I__8269 (
            .O(N__42521),
            .I(\c0.n21686 ));
    Odrv4 I__8268 (
            .O(N__42518),
            .I(\c0.n21686 ));
    Odrv4 I__8267 (
            .O(N__42515),
            .I(\c0.n21686 ));
    CascadeMux I__8266 (
            .O(N__42508),
            .I(N__42503));
    CascadeMux I__8265 (
            .O(N__42507),
            .I(N__42499));
    InMux I__8264 (
            .O(N__42506),
            .I(N__42495));
    InMux I__8263 (
            .O(N__42503),
            .I(N__42490));
    InMux I__8262 (
            .O(N__42502),
            .I(N__42487));
    InMux I__8261 (
            .O(N__42499),
            .I(N__42484));
    InMux I__8260 (
            .O(N__42498),
            .I(N__42481));
    LocalMux I__8259 (
            .O(N__42495),
            .I(N__42478));
    InMux I__8258 (
            .O(N__42494),
            .I(N__42473));
    InMux I__8257 (
            .O(N__42493),
            .I(N__42473));
    LocalMux I__8256 (
            .O(N__42490),
            .I(N__42470));
    LocalMux I__8255 (
            .O(N__42487),
            .I(N__42463));
    LocalMux I__8254 (
            .O(N__42484),
            .I(N__42463));
    LocalMux I__8253 (
            .O(N__42481),
            .I(N__42463));
    Span4Mux_h I__8252 (
            .O(N__42478),
            .I(N__42460));
    LocalMux I__8251 (
            .O(N__42473),
            .I(N__42453));
    Span4Mux_v I__8250 (
            .O(N__42470),
            .I(N__42453));
    Span4Mux_v I__8249 (
            .O(N__42463),
            .I(N__42453));
    Odrv4 I__8248 (
            .O(N__42460),
            .I(\c0.FRAME_MATCHER_state_3 ));
    Odrv4 I__8247 (
            .O(N__42453),
            .I(\c0.FRAME_MATCHER_state_3 ));
    CascadeMux I__8246 (
            .O(N__42448),
            .I(\c0.n21686_cascade_ ));
    SRMux I__8245 (
            .O(N__42445),
            .I(N__42442));
    LocalMux I__8244 (
            .O(N__42442),
            .I(N__42439));
    Span4Mux_h I__8243 (
            .O(N__42439),
            .I(N__42436));
    Odrv4 I__8242 (
            .O(N__42436),
            .I(\c0.n21334 ));
    CascadeMux I__8241 (
            .O(N__42433),
            .I(N__42430));
    InMux I__8240 (
            .O(N__42430),
            .I(N__42426));
    InMux I__8239 (
            .O(N__42429),
            .I(N__42423));
    LocalMux I__8238 (
            .O(N__42426),
            .I(N__42420));
    LocalMux I__8237 (
            .O(N__42423),
            .I(N__42417));
    Span4Mux_h I__8236 (
            .O(N__42420),
            .I(N__42412));
    Span4Mux_h I__8235 (
            .O(N__42417),
            .I(N__42412));
    Odrv4 I__8234 (
            .O(N__42412),
            .I(\c0.n44_adj_4336 ));
    InMux I__8233 (
            .O(N__42409),
            .I(N__42406));
    LocalMux I__8232 (
            .O(N__42406),
            .I(\c0.n1_adj_4349 ));
    CascadeMux I__8231 (
            .O(N__42403),
            .I(N__42400));
    InMux I__8230 (
            .O(N__42400),
            .I(N__42397));
    LocalMux I__8229 (
            .O(N__42397),
            .I(N__42392));
    InMux I__8228 (
            .O(N__42396),
            .I(N__42389));
    InMux I__8227 (
            .O(N__42395),
            .I(N__42386));
    Span4Mux_v I__8226 (
            .O(N__42392),
            .I(N__42382));
    LocalMux I__8225 (
            .O(N__42389),
            .I(N__42379));
    LocalMux I__8224 (
            .O(N__42386),
            .I(N__42376));
    InMux I__8223 (
            .O(N__42385),
            .I(N__42372));
    Sp12to4 I__8222 (
            .O(N__42382),
            .I(N__42367));
    Span12Mux_v I__8221 (
            .O(N__42379),
            .I(N__42367));
    Span4Mux_v I__8220 (
            .O(N__42376),
            .I(N__42364));
    InMux I__8219 (
            .O(N__42375),
            .I(N__42361));
    LocalMux I__8218 (
            .O(N__42372),
            .I(control_mode_4));
    Odrv12 I__8217 (
            .O(N__42367),
            .I(control_mode_4));
    Odrv4 I__8216 (
            .O(N__42364),
            .I(control_mode_4));
    LocalMux I__8215 (
            .O(N__42361),
            .I(control_mode_4));
    CascadeMux I__8214 (
            .O(N__42352),
            .I(N__42348));
    InMux I__8213 (
            .O(N__42351),
            .I(N__42345));
    InMux I__8212 (
            .O(N__42348),
            .I(N__42342));
    LocalMux I__8211 (
            .O(N__42345),
            .I(N__42339));
    LocalMux I__8210 (
            .O(N__42342),
            .I(N__42333));
    Span4Mux_h I__8209 (
            .O(N__42339),
            .I(N__42330));
    InMux I__8208 (
            .O(N__42338),
            .I(N__42325));
    InMux I__8207 (
            .O(N__42337),
            .I(N__42325));
    InMux I__8206 (
            .O(N__42336),
            .I(N__42322));
    Span4Mux_h I__8205 (
            .O(N__42333),
            .I(N__42315));
    Span4Mux_v I__8204 (
            .O(N__42330),
            .I(N__42315));
    LocalMux I__8203 (
            .O(N__42325),
            .I(N__42315));
    LocalMux I__8202 (
            .O(N__42322),
            .I(control_mode_7));
    Odrv4 I__8201 (
            .O(N__42315),
            .I(control_mode_7));
    CascadeMux I__8200 (
            .O(N__42310),
            .I(n23726_cascade_));
    InMux I__8199 (
            .O(N__42307),
            .I(N__42303));
    CascadeMux I__8198 (
            .O(N__42306),
            .I(N__42300));
    LocalMux I__8197 (
            .O(N__42303),
            .I(N__42297));
    InMux I__8196 (
            .O(N__42300),
            .I(N__42294));
    Span4Mux_v I__8195 (
            .O(N__42297),
            .I(N__42290));
    LocalMux I__8194 (
            .O(N__42294),
            .I(N__42287));
    InMux I__8193 (
            .O(N__42293),
            .I(N__42283));
    Sp12to4 I__8192 (
            .O(N__42290),
            .I(N__42280));
    Span4Mux_h I__8191 (
            .O(N__42287),
            .I(N__42277));
    InMux I__8190 (
            .O(N__42286),
            .I(N__42274));
    LocalMux I__8189 (
            .O(N__42283),
            .I(control_mode_6));
    Odrv12 I__8188 (
            .O(N__42280),
            .I(control_mode_6));
    Odrv4 I__8187 (
            .O(N__42277),
            .I(control_mode_6));
    LocalMux I__8186 (
            .O(N__42274),
            .I(control_mode_6));
    InMux I__8185 (
            .O(N__42265),
            .I(N__42262));
    LocalMux I__8184 (
            .O(N__42262),
            .I(N__42259));
    Span4Mux_h I__8183 (
            .O(N__42259),
            .I(N__42256));
    Odrv4 I__8182 (
            .O(N__42256),
            .I(n2249));
    CascadeMux I__8181 (
            .O(N__42253),
            .I(N__42245));
    CascadeMux I__8180 (
            .O(N__42252),
            .I(N__42242));
    InMux I__8179 (
            .O(N__42251),
            .I(N__42224));
    InMux I__8178 (
            .O(N__42250),
            .I(N__42224));
    InMux I__8177 (
            .O(N__42249),
            .I(N__42224));
    InMux I__8176 (
            .O(N__42248),
            .I(N__42210));
    InMux I__8175 (
            .O(N__42245),
            .I(N__42210));
    InMux I__8174 (
            .O(N__42242),
            .I(N__42210));
    InMux I__8173 (
            .O(N__42241),
            .I(N__42210));
    InMux I__8172 (
            .O(N__42240),
            .I(N__42210));
    CascadeMux I__8171 (
            .O(N__42239),
            .I(N__42205));
    InMux I__8170 (
            .O(N__42238),
            .I(N__42199));
    InMux I__8169 (
            .O(N__42237),
            .I(N__42190));
    InMux I__8168 (
            .O(N__42236),
            .I(N__42190));
    InMux I__8167 (
            .O(N__42235),
            .I(N__42190));
    InMux I__8166 (
            .O(N__42234),
            .I(N__42190));
    InMux I__8165 (
            .O(N__42233),
            .I(N__42187));
    InMux I__8164 (
            .O(N__42232),
            .I(N__42184));
    CascadeMux I__8163 (
            .O(N__42231),
            .I(N__42181));
    LocalMux I__8162 (
            .O(N__42224),
            .I(N__42177));
    InMux I__8161 (
            .O(N__42223),
            .I(N__42172));
    InMux I__8160 (
            .O(N__42222),
            .I(N__42172));
    CascadeMux I__8159 (
            .O(N__42221),
            .I(N__42169));
    LocalMux I__8158 (
            .O(N__42210),
            .I(N__42164));
    InMux I__8157 (
            .O(N__42209),
            .I(N__42155));
    InMux I__8156 (
            .O(N__42208),
            .I(N__42155));
    InMux I__8155 (
            .O(N__42205),
            .I(N__42155));
    InMux I__8154 (
            .O(N__42204),
            .I(N__42155));
    CascadeMux I__8153 (
            .O(N__42203),
            .I(N__42152));
    InMux I__8152 (
            .O(N__42202),
            .I(N__42147));
    LocalMux I__8151 (
            .O(N__42199),
            .I(N__42138));
    LocalMux I__8150 (
            .O(N__42190),
            .I(N__42138));
    LocalMux I__8149 (
            .O(N__42187),
            .I(N__42138));
    LocalMux I__8148 (
            .O(N__42184),
            .I(N__42138));
    InMux I__8147 (
            .O(N__42181),
            .I(N__42133));
    InMux I__8146 (
            .O(N__42180),
            .I(N__42133));
    Span4Mux_h I__8145 (
            .O(N__42177),
            .I(N__42128));
    LocalMux I__8144 (
            .O(N__42172),
            .I(N__42128));
    InMux I__8143 (
            .O(N__42169),
            .I(N__42123));
    InMux I__8142 (
            .O(N__42168),
            .I(N__42123));
    InMux I__8141 (
            .O(N__42167),
            .I(N__42120));
    Span4Mux_v I__8140 (
            .O(N__42164),
            .I(N__42115));
    LocalMux I__8139 (
            .O(N__42155),
            .I(N__42115));
    InMux I__8138 (
            .O(N__42152),
            .I(N__42108));
    InMux I__8137 (
            .O(N__42151),
            .I(N__42108));
    InMux I__8136 (
            .O(N__42150),
            .I(N__42108));
    LocalMux I__8135 (
            .O(N__42147),
            .I(N__42103));
    Span4Mux_v I__8134 (
            .O(N__42138),
            .I(N__42100));
    LocalMux I__8133 (
            .O(N__42133),
            .I(N__42097));
    Span4Mux_h I__8132 (
            .O(N__42128),
            .I(N__42090));
    LocalMux I__8131 (
            .O(N__42123),
            .I(N__42090));
    LocalMux I__8130 (
            .O(N__42120),
            .I(N__42090));
    Span4Mux_v I__8129 (
            .O(N__42115),
            .I(N__42085));
    LocalMux I__8128 (
            .O(N__42108),
            .I(N__42085));
    InMux I__8127 (
            .O(N__42107),
            .I(N__42082));
    InMux I__8126 (
            .O(N__42106),
            .I(N__42079));
    Span4Mux_v I__8125 (
            .O(N__42103),
            .I(N__42076));
    Span4Mux_h I__8124 (
            .O(N__42100),
            .I(N__42071));
    Span4Mux_v I__8123 (
            .O(N__42097),
            .I(N__42071));
    Span4Mux_v I__8122 (
            .O(N__42090),
            .I(N__42062));
    Span4Mux_h I__8121 (
            .O(N__42085),
            .I(N__42062));
    LocalMux I__8120 (
            .O(N__42082),
            .I(N__42062));
    LocalMux I__8119 (
            .O(N__42079),
            .I(N__42062));
    Span4Mux_v I__8118 (
            .O(N__42076),
            .I(N__42059));
    Span4Mux_v I__8117 (
            .O(N__42071),
            .I(N__42056));
    Span4Mux_h I__8116 (
            .O(N__42062),
            .I(N__42053));
    Odrv4 I__8115 (
            .O(N__42059),
            .I(count_enable));
    Odrv4 I__8114 (
            .O(N__42056),
            .I(count_enable));
    Odrv4 I__8113 (
            .O(N__42053),
            .I(count_enable));
    InMux I__8112 (
            .O(N__42046),
            .I(N__42042));
    InMux I__8111 (
            .O(N__42045),
            .I(N__42038));
    LocalMux I__8110 (
            .O(N__42042),
            .I(N__42035));
    CascadeMux I__8109 (
            .O(N__42041),
            .I(N__42031));
    LocalMux I__8108 (
            .O(N__42038),
            .I(N__42027));
    Span4Mux_h I__8107 (
            .O(N__42035),
            .I(N__42024));
    InMux I__8106 (
            .O(N__42034),
            .I(N__42021));
    InMux I__8105 (
            .O(N__42031),
            .I(N__42018));
    InMux I__8104 (
            .O(N__42030),
            .I(N__42015));
    Span4Mux_h I__8103 (
            .O(N__42027),
            .I(N__42010));
    Span4Mux_v I__8102 (
            .O(N__42024),
            .I(N__42010));
    LocalMux I__8101 (
            .O(N__42021),
            .I(N__42007));
    LocalMux I__8100 (
            .O(N__42018),
            .I(encoder0_position_22));
    LocalMux I__8099 (
            .O(N__42015),
            .I(encoder0_position_22));
    Odrv4 I__8098 (
            .O(N__42010),
            .I(encoder0_position_22));
    Odrv4 I__8097 (
            .O(N__42007),
            .I(encoder0_position_22));
    InMux I__8096 (
            .O(N__41998),
            .I(N__41995));
    LocalMux I__8095 (
            .O(N__41995),
            .I(N__41989));
    InMux I__8094 (
            .O(N__41994),
            .I(N__41986));
    InMux I__8093 (
            .O(N__41993),
            .I(N__41981));
    InMux I__8092 (
            .O(N__41992),
            .I(N__41981));
    Span4Mux_v I__8091 (
            .O(N__41989),
            .I(N__41976));
    LocalMux I__8090 (
            .O(N__41986),
            .I(N__41976));
    LocalMux I__8089 (
            .O(N__41981),
            .I(N__41971));
    Span4Mux_h I__8088 (
            .O(N__41976),
            .I(N__41971));
    Odrv4 I__8087 (
            .O(N__41971),
            .I(data_in_2_4));
    InMux I__8086 (
            .O(N__41968),
            .I(N__41964));
    InMux I__8085 (
            .O(N__41967),
            .I(N__41961));
    LocalMux I__8084 (
            .O(N__41964),
            .I(N__41957));
    LocalMux I__8083 (
            .O(N__41961),
            .I(N__41954));
    CascadeMux I__8082 (
            .O(N__41960),
            .I(N__41951));
    Span4Mux_v I__8081 (
            .O(N__41957),
            .I(N__41947));
    Span4Mux_v I__8080 (
            .O(N__41954),
            .I(N__41944));
    InMux I__8079 (
            .O(N__41951),
            .I(N__41941));
    InMux I__8078 (
            .O(N__41950),
            .I(N__41938));
    Span4Mux_h I__8077 (
            .O(N__41947),
            .I(N__41935));
    Sp12to4 I__8076 (
            .O(N__41944),
            .I(N__41930));
    LocalMux I__8075 (
            .O(N__41941),
            .I(N__41930));
    LocalMux I__8074 (
            .O(N__41938),
            .I(data_in_1_4));
    Odrv4 I__8073 (
            .O(N__41935),
            .I(data_in_1_4));
    Odrv12 I__8072 (
            .O(N__41930),
            .I(data_in_1_4));
    InMux I__8071 (
            .O(N__41923),
            .I(N__41920));
    LocalMux I__8070 (
            .O(N__41920),
            .I(N__41917));
    Span4Mux_h I__8069 (
            .O(N__41917),
            .I(N__41914));
    Span4Mux_h I__8068 (
            .O(N__41914),
            .I(N__41910));
    InMux I__8067 (
            .O(N__41913),
            .I(N__41907));
    Span4Mux_v I__8066 (
            .O(N__41910),
            .I(N__41904));
    LocalMux I__8065 (
            .O(N__41907),
            .I(\c0.FRAME_MATCHER_rx_data_ready_prev ));
    Odrv4 I__8064 (
            .O(N__41904),
            .I(\c0.FRAME_MATCHER_rx_data_ready_prev ));
    CascadeMux I__8063 (
            .O(N__41899),
            .I(\c0.n17790_cascade_ ));
    CascadeMux I__8062 (
            .O(N__41896),
            .I(\c0.n21775_cascade_ ));
    InMux I__8061 (
            .O(N__41893),
            .I(N__41890));
    LocalMux I__8060 (
            .O(N__41890),
            .I(N__41885));
    InMux I__8059 (
            .O(N__41889),
            .I(N__41880));
    InMux I__8058 (
            .O(N__41888),
            .I(N__41880));
    Span4Mux_h I__8057 (
            .O(N__41885),
            .I(N__41877));
    LocalMux I__8056 (
            .O(N__41880),
            .I(data_in_3_4));
    Odrv4 I__8055 (
            .O(N__41877),
            .I(data_in_3_4));
    InMux I__8054 (
            .O(N__41872),
            .I(N__41866));
    InMux I__8053 (
            .O(N__41871),
            .I(N__41863));
    InMux I__8052 (
            .O(N__41870),
            .I(N__41859));
    InMux I__8051 (
            .O(N__41869),
            .I(N__41856));
    LocalMux I__8050 (
            .O(N__41866),
            .I(N__41853));
    LocalMux I__8049 (
            .O(N__41863),
            .I(N__41850));
    InMux I__8048 (
            .O(N__41862),
            .I(N__41847));
    LocalMux I__8047 (
            .O(N__41859),
            .I(N__41844));
    LocalMux I__8046 (
            .O(N__41856),
            .I(N__41840));
    Span4Mux_v I__8045 (
            .O(N__41853),
            .I(N__41833));
    Span4Mux_v I__8044 (
            .O(N__41850),
            .I(N__41833));
    LocalMux I__8043 (
            .O(N__41847),
            .I(N__41833));
    Span4Mux_h I__8042 (
            .O(N__41844),
            .I(N__41830));
    InMux I__8041 (
            .O(N__41843),
            .I(N__41827));
    Span4Mux_v I__8040 (
            .O(N__41840),
            .I(N__41822));
    Span4Mux_h I__8039 (
            .O(N__41833),
            .I(N__41822));
    Odrv4 I__8038 (
            .O(N__41830),
            .I(control_mode_1));
    LocalMux I__8037 (
            .O(N__41827),
            .I(control_mode_1));
    Odrv4 I__8036 (
            .O(N__41822),
            .I(control_mode_1));
    CascadeMux I__8035 (
            .O(N__41815),
            .I(N__41812));
    InMux I__8034 (
            .O(N__41812),
            .I(N__41807));
    InMux I__8033 (
            .O(N__41811),
            .I(N__41804));
    InMux I__8032 (
            .O(N__41810),
            .I(N__41801));
    LocalMux I__8031 (
            .O(N__41807),
            .I(N__41796));
    LocalMux I__8030 (
            .O(N__41804),
            .I(N__41791));
    LocalMux I__8029 (
            .O(N__41801),
            .I(N__41791));
    InMux I__8028 (
            .O(N__41800),
            .I(N__41788));
    InMux I__8027 (
            .O(N__41799),
            .I(N__41785));
    Span4Mux_v I__8026 (
            .O(N__41796),
            .I(N__41781));
    Span4Mux_v I__8025 (
            .O(N__41791),
            .I(N__41774));
    LocalMux I__8024 (
            .O(N__41788),
            .I(N__41774));
    LocalMux I__8023 (
            .O(N__41785),
            .I(N__41774));
    InMux I__8022 (
            .O(N__41784),
            .I(N__41771));
    Span4Mux_h I__8021 (
            .O(N__41781),
            .I(N__41768));
    Span4Mux_h I__8020 (
            .O(N__41774),
            .I(N__41765));
    LocalMux I__8019 (
            .O(N__41771),
            .I(control_mode_3));
    Odrv4 I__8018 (
            .O(N__41768),
            .I(control_mode_3));
    Odrv4 I__8017 (
            .O(N__41765),
            .I(control_mode_3));
    CascadeMux I__8016 (
            .O(N__41758),
            .I(N__41755));
    InMux I__8015 (
            .O(N__41755),
            .I(N__41751));
    InMux I__8014 (
            .O(N__41754),
            .I(N__41747));
    LocalMux I__8013 (
            .O(N__41751),
            .I(N__41741));
    InMux I__8012 (
            .O(N__41750),
            .I(N__41738));
    LocalMux I__8011 (
            .O(N__41747),
            .I(N__41735));
    InMux I__8010 (
            .O(N__41746),
            .I(N__41728));
    InMux I__8009 (
            .O(N__41745),
            .I(N__41728));
    InMux I__8008 (
            .O(N__41744),
            .I(N__41728));
    Span4Mux_h I__8007 (
            .O(N__41741),
            .I(N__41723));
    LocalMux I__8006 (
            .O(N__41738),
            .I(N__41723));
    Span4Mux_h I__8005 (
            .O(N__41735),
            .I(N__41719));
    LocalMux I__8004 (
            .O(N__41728),
            .I(N__41714));
    Span4Mux_h I__8003 (
            .O(N__41723),
            .I(N__41714));
    InMux I__8002 (
            .O(N__41722),
            .I(N__41711));
    Odrv4 I__8001 (
            .O(N__41719),
            .I(encoder0_position_18));
    Odrv4 I__8000 (
            .O(N__41714),
            .I(encoder0_position_18));
    LocalMux I__7999 (
            .O(N__41711),
            .I(encoder0_position_18));
    CascadeMux I__7998 (
            .O(N__41704),
            .I(N__41701));
    InMux I__7997 (
            .O(N__41701),
            .I(N__41697));
    InMux I__7996 (
            .O(N__41700),
            .I(N__41693));
    LocalMux I__7995 (
            .O(N__41697),
            .I(N__41690));
    InMux I__7994 (
            .O(N__41696),
            .I(N__41687));
    LocalMux I__7993 (
            .O(N__41693),
            .I(N__41684));
    Span4Mux_v I__7992 (
            .O(N__41690),
            .I(N__41679));
    LocalMux I__7991 (
            .O(N__41687),
            .I(N__41674));
    Span4Mux_v I__7990 (
            .O(N__41684),
            .I(N__41674));
    CascadeMux I__7989 (
            .O(N__41683),
            .I(N__41670));
    InMux I__7988 (
            .O(N__41682),
            .I(N__41667));
    Span4Mux_h I__7987 (
            .O(N__41679),
            .I(N__41662));
    Span4Mux_h I__7986 (
            .O(N__41674),
            .I(N__41662));
    InMux I__7985 (
            .O(N__41673),
            .I(N__41657));
    InMux I__7984 (
            .O(N__41670),
            .I(N__41657));
    LocalMux I__7983 (
            .O(N__41667),
            .I(encoder0_position_3));
    Odrv4 I__7982 (
            .O(N__41662),
            .I(encoder0_position_3));
    LocalMux I__7981 (
            .O(N__41657),
            .I(encoder0_position_3));
    InMux I__7980 (
            .O(N__41650),
            .I(N__41642));
    InMux I__7979 (
            .O(N__41649),
            .I(N__41635));
    InMux I__7978 (
            .O(N__41648),
            .I(N__41635));
    InMux I__7977 (
            .O(N__41647),
            .I(N__41635));
    InMux I__7976 (
            .O(N__41646),
            .I(N__41632));
    CascadeMux I__7975 (
            .O(N__41645),
            .I(N__41629));
    LocalMux I__7974 (
            .O(N__41642),
            .I(N__41623));
    LocalMux I__7973 (
            .O(N__41635),
            .I(N__41623));
    LocalMux I__7972 (
            .O(N__41632),
            .I(N__41620));
    InMux I__7971 (
            .O(N__41629),
            .I(N__41615));
    InMux I__7970 (
            .O(N__41628),
            .I(N__41615));
    Span4Mux_h I__7969 (
            .O(N__41623),
            .I(N__41612));
    Odrv12 I__7968 (
            .O(N__41620),
            .I(encoder0_position_31));
    LocalMux I__7967 (
            .O(N__41615),
            .I(encoder0_position_31));
    Odrv4 I__7966 (
            .O(N__41612),
            .I(encoder0_position_31));
    CascadeMux I__7965 (
            .O(N__41605),
            .I(N__41602));
    InMux I__7964 (
            .O(N__41602),
            .I(N__41598));
    InMux I__7963 (
            .O(N__41601),
            .I(N__41595));
    LocalMux I__7962 (
            .O(N__41598),
            .I(N__41592));
    LocalMux I__7961 (
            .O(N__41595),
            .I(N__41587));
    Span4Mux_v I__7960 (
            .O(N__41592),
            .I(N__41587));
    Span4Mux_h I__7959 (
            .O(N__41587),
            .I(N__41584));
    Odrv4 I__7958 (
            .O(N__41584),
            .I(\c0.n21813 ));
    CascadeMux I__7957 (
            .O(N__41581),
            .I(N__41578));
    InMux I__7956 (
            .O(N__41578),
            .I(N__41574));
    InMux I__7955 (
            .O(N__41577),
            .I(N__41571));
    LocalMux I__7954 (
            .O(N__41574),
            .I(N__41568));
    LocalMux I__7953 (
            .O(N__41571),
            .I(data_in_frame_6_5));
    Odrv12 I__7952 (
            .O(N__41568),
            .I(data_in_frame_6_5));
    InMux I__7951 (
            .O(N__41563),
            .I(N__41560));
    LocalMux I__7950 (
            .O(N__41560),
            .I(N__41557));
    Span4Mux_h I__7949 (
            .O(N__41557),
            .I(N__41554));
    Span4Mux_v I__7948 (
            .O(N__41554),
            .I(N__41551));
    Odrv4 I__7947 (
            .O(N__41551),
            .I(\c0.tx.n23987 ));
    InMux I__7946 (
            .O(N__41548),
            .I(N__41541));
    InMux I__7945 (
            .O(N__41547),
            .I(N__41541));
    InMux I__7944 (
            .O(N__41546),
            .I(N__41538));
    LocalMux I__7943 (
            .O(N__41541),
            .I(N__41535));
    LocalMux I__7942 (
            .O(N__41538),
            .I(N__41531));
    Span4Mux_h I__7941 (
            .O(N__41535),
            .I(N__41528));
    InMux I__7940 (
            .O(N__41534),
            .I(N__41525));
    Span12Mux_h I__7939 (
            .O(N__41531),
            .I(N__41522));
    Span4Mux_v I__7938 (
            .O(N__41528),
            .I(N__41519));
    LocalMux I__7937 (
            .O(N__41525),
            .I(\c0.tx.r_Clock_Count_6 ));
    Odrv12 I__7936 (
            .O(N__41522),
            .I(\c0.tx.r_Clock_Count_6 ));
    Odrv4 I__7935 (
            .O(N__41519),
            .I(\c0.tx.r_Clock_Count_6 ));
    InMux I__7934 (
            .O(N__41512),
            .I(N__41509));
    LocalMux I__7933 (
            .O(N__41509),
            .I(N__41506));
    Span4Mux_v I__7932 (
            .O(N__41506),
            .I(N__41503));
    Span4Mux_h I__7931 (
            .O(N__41503),
            .I(N__41500));
    Odrv4 I__7930 (
            .O(N__41500),
            .I(n313));
    CascadeMux I__7929 (
            .O(N__41497),
            .I(N__41493));
    CascadeMux I__7928 (
            .O(N__41496),
            .I(N__41487));
    InMux I__7927 (
            .O(N__41493),
            .I(N__41479));
    InMux I__7926 (
            .O(N__41492),
            .I(N__41479));
    InMux I__7925 (
            .O(N__41491),
            .I(N__41476));
    InMux I__7924 (
            .O(N__41490),
            .I(N__41471));
    InMux I__7923 (
            .O(N__41487),
            .I(N__41471));
    InMux I__7922 (
            .O(N__41486),
            .I(N__41468));
    InMux I__7921 (
            .O(N__41485),
            .I(N__41462));
    InMux I__7920 (
            .O(N__41484),
            .I(N__41462));
    LocalMux I__7919 (
            .O(N__41479),
            .I(N__41459));
    LocalMux I__7918 (
            .O(N__41476),
            .I(N__41451));
    LocalMux I__7917 (
            .O(N__41471),
            .I(N__41446));
    LocalMux I__7916 (
            .O(N__41468),
            .I(N__41446));
    CascadeMux I__7915 (
            .O(N__41467),
            .I(N__41440));
    LocalMux I__7914 (
            .O(N__41462),
            .I(N__41437));
    Span4Mux_h I__7913 (
            .O(N__41459),
            .I(N__41434));
    InMux I__7912 (
            .O(N__41458),
            .I(N__41429));
    InMux I__7911 (
            .O(N__41457),
            .I(N__41429));
    InMux I__7910 (
            .O(N__41456),
            .I(N__41422));
    InMux I__7909 (
            .O(N__41455),
            .I(N__41422));
    InMux I__7908 (
            .O(N__41454),
            .I(N__41422));
    Span4Mux_h I__7907 (
            .O(N__41451),
            .I(N__41419));
    Span4Mux_v I__7906 (
            .O(N__41446),
            .I(N__41416));
    InMux I__7905 (
            .O(N__41445),
            .I(N__41413));
    InMux I__7904 (
            .O(N__41444),
            .I(N__41406));
    InMux I__7903 (
            .O(N__41443),
            .I(N__41406));
    InMux I__7902 (
            .O(N__41440),
            .I(N__41406));
    Span4Mux_v I__7901 (
            .O(N__41437),
            .I(N__41399));
    Span4Mux_v I__7900 (
            .O(N__41434),
            .I(N__41399));
    LocalMux I__7899 (
            .O(N__41429),
            .I(N__41399));
    LocalMux I__7898 (
            .O(N__41422),
            .I(r_SM_Main_2_adj_4549));
    Odrv4 I__7897 (
            .O(N__41419),
            .I(r_SM_Main_2_adj_4549));
    Odrv4 I__7896 (
            .O(N__41416),
            .I(r_SM_Main_2_adj_4549));
    LocalMux I__7895 (
            .O(N__41413),
            .I(r_SM_Main_2_adj_4549));
    LocalMux I__7894 (
            .O(N__41406),
            .I(r_SM_Main_2_adj_4549));
    Odrv4 I__7893 (
            .O(N__41399),
            .I(r_SM_Main_2_adj_4549));
    InMux I__7892 (
            .O(N__41386),
            .I(N__41383));
    LocalMux I__7891 (
            .O(N__41383),
            .I(N__41379));
    InMux I__7890 (
            .O(N__41382),
            .I(N__41370));
    Span4Mux_h I__7889 (
            .O(N__41379),
            .I(N__41367));
    InMux I__7888 (
            .O(N__41378),
            .I(N__41362));
    InMux I__7887 (
            .O(N__41377),
            .I(N__41362));
    InMux I__7886 (
            .O(N__41376),
            .I(N__41353));
    InMux I__7885 (
            .O(N__41375),
            .I(N__41353));
    InMux I__7884 (
            .O(N__41374),
            .I(N__41353));
    InMux I__7883 (
            .O(N__41373),
            .I(N__41353));
    LocalMux I__7882 (
            .O(N__41370),
            .I(n8));
    Odrv4 I__7881 (
            .O(N__41367),
            .I(n8));
    LocalMux I__7880 (
            .O(N__41362),
            .I(n8));
    LocalMux I__7879 (
            .O(N__41353),
            .I(n8));
    InMux I__7878 (
            .O(N__41344),
            .I(N__41339));
    InMux I__7877 (
            .O(N__41343),
            .I(N__41334));
    InMux I__7876 (
            .O(N__41342),
            .I(N__41334));
    LocalMux I__7875 (
            .O(N__41339),
            .I(N__41331));
    LocalMux I__7874 (
            .O(N__41334),
            .I(N__41328));
    Span4Mux_v I__7873 (
            .O(N__41331),
            .I(N__41324));
    Span4Mux_h I__7872 (
            .O(N__41328),
            .I(N__41321));
    InMux I__7871 (
            .O(N__41327),
            .I(N__41318));
    Span4Mux_h I__7870 (
            .O(N__41324),
            .I(N__41315));
    Span4Mux_v I__7869 (
            .O(N__41321),
            .I(N__41312));
    LocalMux I__7868 (
            .O(N__41318),
            .I(r_Clock_Count_8));
    Odrv4 I__7867 (
            .O(N__41315),
            .I(r_Clock_Count_8));
    Odrv4 I__7866 (
            .O(N__41312),
            .I(r_Clock_Count_8));
    InMux I__7865 (
            .O(N__41305),
            .I(N__41302));
    LocalMux I__7864 (
            .O(N__41302),
            .I(N__41299));
    Span4Mux_h I__7863 (
            .O(N__41299),
            .I(N__41296));
    Odrv4 I__7862 (
            .O(N__41296),
            .I(n2253));
    InMux I__7861 (
            .O(N__41293),
            .I(N__41290));
    LocalMux I__7860 (
            .O(N__41290),
            .I(N__41287));
    Span12Mux_h I__7859 (
            .O(N__41287),
            .I(N__41284));
    Odrv12 I__7858 (
            .O(N__41284),
            .I(\c0.n21816 ));
    CascadeMux I__7857 (
            .O(N__41281),
            .I(\c0.n21740_cascade_ ));
    InMux I__7856 (
            .O(N__41278),
            .I(N__41274));
    CascadeMux I__7855 (
            .O(N__41277),
            .I(N__41271));
    LocalMux I__7854 (
            .O(N__41274),
            .I(N__41268));
    InMux I__7853 (
            .O(N__41271),
            .I(N__41265));
    Span4Mux_v I__7852 (
            .O(N__41268),
            .I(N__41262));
    LocalMux I__7851 (
            .O(N__41265),
            .I(\c0.data_in_frame_20_6 ));
    Odrv4 I__7850 (
            .O(N__41262),
            .I(\c0.data_in_frame_20_6 ));
    CascadeMux I__7849 (
            .O(N__41257),
            .I(n21744_cascade_));
    InMux I__7848 (
            .O(N__41254),
            .I(N__41250));
    InMux I__7847 (
            .O(N__41253),
            .I(N__41247));
    LocalMux I__7846 (
            .O(N__41250),
            .I(N__41244));
    LocalMux I__7845 (
            .O(N__41247),
            .I(data_in_frame_6_3));
    Odrv12 I__7844 (
            .O(N__41244),
            .I(data_in_frame_6_3));
    InMux I__7843 (
            .O(N__41239),
            .I(N__41236));
    LocalMux I__7842 (
            .O(N__41236),
            .I(N__41233));
    Span4Mux_h I__7841 (
            .O(N__41233),
            .I(N__41230));
    Odrv4 I__7840 (
            .O(N__41230),
            .I(\c0.n25_adj_4408 ));
    CascadeMux I__7839 (
            .O(N__41227),
            .I(N__41224));
    InMux I__7838 (
            .O(N__41224),
            .I(N__41221));
    LocalMux I__7837 (
            .O(N__41221),
            .I(N__41218));
    Odrv4 I__7836 (
            .O(N__41218),
            .I(\c0.n23648 ));
    InMux I__7835 (
            .O(N__41215),
            .I(N__41212));
    LocalMux I__7834 (
            .O(N__41212),
            .I(\c0.n16_adj_4401 ));
    InMux I__7833 (
            .O(N__41209),
            .I(N__41205));
    InMux I__7832 (
            .O(N__41208),
            .I(N__41202));
    LocalMux I__7831 (
            .O(N__41205),
            .I(\c0.n21893 ));
    LocalMux I__7830 (
            .O(N__41202),
            .I(\c0.n21893 ));
    InMux I__7829 (
            .O(N__41197),
            .I(N__41194));
    LocalMux I__7828 (
            .O(N__41194),
            .I(N__41191));
    Odrv12 I__7827 (
            .O(N__41191),
            .I(\c0.n44_adj_4409 ));
    CascadeMux I__7826 (
            .O(N__41188),
            .I(\c0.n6_adj_4393_cascade_ ));
    CascadeMux I__7825 (
            .O(N__41185),
            .I(\c0.n13086_cascade_ ));
    CascadeMux I__7824 (
            .O(N__41182),
            .I(\c0.n21986_cascade_ ));
    InMux I__7823 (
            .O(N__41179),
            .I(N__41173));
    InMux I__7822 (
            .O(N__41178),
            .I(N__41173));
    LocalMux I__7821 (
            .O(N__41173),
            .I(data_in_frame_6_0));
    CascadeMux I__7820 (
            .O(N__41170),
            .I(\c0.n38_adj_4407_cascade_ ));
    InMux I__7819 (
            .O(N__41167),
            .I(N__41164));
    LocalMux I__7818 (
            .O(N__41164),
            .I(\c0.n23836 ));
    CascadeMux I__7817 (
            .O(N__41161),
            .I(\c0.n43_adj_4410_cascade_ ));
    CascadeMux I__7816 (
            .O(N__41158),
            .I(\c0.n22443_cascade_ ));
    CascadeMux I__7815 (
            .O(N__41155),
            .I(N__41152));
    InMux I__7814 (
            .O(N__41152),
            .I(N__41148));
    InMux I__7813 (
            .O(N__41151),
            .I(N__41143));
    LocalMux I__7812 (
            .O(N__41148),
            .I(N__41140));
    InMux I__7811 (
            .O(N__41147),
            .I(N__41135));
    InMux I__7810 (
            .O(N__41146),
            .I(N__41135));
    LocalMux I__7809 (
            .O(N__41143),
            .I(N__41132));
    Span4Mux_h I__7808 (
            .O(N__41140),
            .I(N__41129));
    LocalMux I__7807 (
            .O(N__41135),
            .I(\c0.FRAME_MATCHER_state_30 ));
    Odrv4 I__7806 (
            .O(N__41132),
            .I(\c0.FRAME_MATCHER_state_30 ));
    Odrv4 I__7805 (
            .O(N__41129),
            .I(\c0.FRAME_MATCHER_state_30 ));
    SRMux I__7804 (
            .O(N__41122),
            .I(N__41119));
    LocalMux I__7803 (
            .O(N__41119),
            .I(N__41116));
    Span4Mux_h I__7802 (
            .O(N__41116),
            .I(N__41113));
    Span4Mux_h I__7801 (
            .O(N__41113),
            .I(N__41110));
    Odrv4 I__7800 (
            .O(N__41110),
            .I(\c0.n8_adj_4396 ));
    CascadeMux I__7799 (
            .O(N__41107),
            .I(\c0.n21737_cascade_ ));
    CascadeMux I__7798 (
            .O(N__41104),
            .I(N__41101));
    InMux I__7797 (
            .O(N__41101),
            .I(N__41096));
    InMux I__7796 (
            .O(N__41100),
            .I(N__41093));
    InMux I__7795 (
            .O(N__41099),
            .I(N__41090));
    LocalMux I__7794 (
            .O(N__41096),
            .I(N__41087));
    LocalMux I__7793 (
            .O(N__41093),
            .I(N__41084));
    LocalMux I__7792 (
            .O(N__41090),
            .I(N__41076));
    Sp12to4 I__7791 (
            .O(N__41087),
            .I(N__41076));
    Sp12to4 I__7790 (
            .O(N__41084),
            .I(N__41076));
    InMux I__7789 (
            .O(N__41083),
            .I(N__41073));
    Span12Mux_v I__7788 (
            .O(N__41076),
            .I(N__41070));
    LocalMux I__7787 (
            .O(N__41073),
            .I(\c0.FRAME_MATCHER_state_6 ));
    Odrv12 I__7786 (
            .O(N__41070),
            .I(\c0.FRAME_MATCHER_state_6 ));
    SRMux I__7785 (
            .O(N__41065),
            .I(N__41062));
    LocalMux I__7784 (
            .O(N__41062),
            .I(N__41059));
    Span12Mux_v I__7783 (
            .O(N__41059),
            .I(N__41056));
    Odrv12 I__7782 (
            .O(N__41056),
            .I(\c0.n21340 ));
    InMux I__7781 (
            .O(N__41053),
            .I(N__41049));
    CascadeMux I__7780 (
            .O(N__41052),
            .I(N__41045));
    LocalMux I__7779 (
            .O(N__41049),
            .I(N__41042));
    InMux I__7778 (
            .O(N__41048),
            .I(N__41038));
    InMux I__7777 (
            .O(N__41045),
            .I(N__41035));
    Span4Mux_v I__7776 (
            .O(N__41042),
            .I(N__41032));
    InMux I__7775 (
            .O(N__41041),
            .I(N__41029));
    LocalMux I__7774 (
            .O(N__41038),
            .I(\c0.FRAME_MATCHER_state_19 ));
    LocalMux I__7773 (
            .O(N__41035),
            .I(\c0.FRAME_MATCHER_state_19 ));
    Odrv4 I__7772 (
            .O(N__41032),
            .I(\c0.FRAME_MATCHER_state_19 ));
    LocalMux I__7771 (
            .O(N__41029),
            .I(\c0.FRAME_MATCHER_state_19 ));
    SRMux I__7770 (
            .O(N__41020),
            .I(N__41017));
    LocalMux I__7769 (
            .O(N__41017),
            .I(N__41014));
    Odrv12 I__7768 (
            .O(N__41014),
            .I(\c0.n8_adj_4398 ));
    CascadeMux I__7767 (
            .O(N__41011),
            .I(N__41008));
    InMux I__7766 (
            .O(N__41008),
            .I(N__41004));
    InMux I__7765 (
            .O(N__41007),
            .I(N__41000));
    LocalMux I__7764 (
            .O(N__41004),
            .I(N__40997));
    InMux I__7763 (
            .O(N__41003),
            .I(N__40993));
    LocalMux I__7762 (
            .O(N__41000),
            .I(N__40990));
    Span4Mux_v I__7761 (
            .O(N__40997),
            .I(N__40987));
    InMux I__7760 (
            .O(N__40996),
            .I(N__40984));
    LocalMux I__7759 (
            .O(N__40993),
            .I(N__40981));
    Span4Mux_h I__7758 (
            .O(N__40990),
            .I(N__40978));
    Span4Mux_h I__7757 (
            .O(N__40987),
            .I(N__40975));
    LocalMux I__7756 (
            .O(N__40984),
            .I(\c0.FRAME_MATCHER_state_5 ));
    Odrv12 I__7755 (
            .O(N__40981),
            .I(\c0.FRAME_MATCHER_state_5 ));
    Odrv4 I__7754 (
            .O(N__40978),
            .I(\c0.FRAME_MATCHER_state_5 ));
    Odrv4 I__7753 (
            .O(N__40975),
            .I(\c0.FRAME_MATCHER_state_5 ));
    SRMux I__7752 (
            .O(N__40966),
            .I(N__40963));
    LocalMux I__7751 (
            .O(N__40963),
            .I(N__40960));
    Span4Mux_h I__7750 (
            .O(N__40960),
            .I(N__40957));
    Odrv4 I__7749 (
            .O(N__40957),
            .I(\c0.n21338 ));
    CEMux I__7748 (
            .O(N__40954),
            .I(N__40947));
    CEMux I__7747 (
            .O(N__40953),
            .I(N__40941));
    CEMux I__7746 (
            .O(N__40952),
            .I(N__40938));
    CEMux I__7745 (
            .O(N__40951),
            .I(N__40935));
    CEMux I__7744 (
            .O(N__40950),
            .I(N__40931));
    LocalMux I__7743 (
            .O(N__40947),
            .I(N__40928));
    CEMux I__7742 (
            .O(N__40946),
            .I(N__40924));
    CEMux I__7741 (
            .O(N__40945),
            .I(N__40921));
    CEMux I__7740 (
            .O(N__40944),
            .I(N__40918));
    LocalMux I__7739 (
            .O(N__40941),
            .I(N__40915));
    LocalMux I__7738 (
            .O(N__40938),
            .I(N__40912));
    LocalMux I__7737 (
            .O(N__40935),
            .I(N__40909));
    SRMux I__7736 (
            .O(N__40934),
            .I(N__40906));
    LocalMux I__7735 (
            .O(N__40931),
            .I(N__40903));
    Span4Mux_v I__7734 (
            .O(N__40928),
            .I(N__40900));
    SRMux I__7733 (
            .O(N__40927),
            .I(N__40897));
    LocalMux I__7732 (
            .O(N__40924),
            .I(N__40894));
    LocalMux I__7731 (
            .O(N__40921),
            .I(N__40891));
    LocalMux I__7730 (
            .O(N__40918),
            .I(N__40886));
    Span4Mux_v I__7729 (
            .O(N__40915),
            .I(N__40886));
    Span4Mux_h I__7728 (
            .O(N__40912),
            .I(N__40883));
    Span4Mux_v I__7727 (
            .O(N__40909),
            .I(N__40880));
    LocalMux I__7726 (
            .O(N__40906),
            .I(N__40877));
    Span4Mux_h I__7725 (
            .O(N__40903),
            .I(N__40874));
    Span4Mux_v I__7724 (
            .O(N__40900),
            .I(N__40871));
    LocalMux I__7723 (
            .O(N__40897),
            .I(N__40868));
    Span4Mux_h I__7722 (
            .O(N__40894),
            .I(N__40865));
    Span4Mux_v I__7721 (
            .O(N__40891),
            .I(N__40858));
    Span4Mux_h I__7720 (
            .O(N__40886),
            .I(N__40858));
    Span4Mux_v I__7719 (
            .O(N__40883),
            .I(N__40858));
    Span4Mux_v I__7718 (
            .O(N__40880),
            .I(N__40855));
    Span4Mux_h I__7717 (
            .O(N__40877),
            .I(N__40852));
    Span4Mux_v I__7716 (
            .O(N__40874),
            .I(N__40849));
    Span4Mux_h I__7715 (
            .O(N__40871),
            .I(N__40846));
    Span4Mux_h I__7714 (
            .O(N__40868),
            .I(N__40843));
    Sp12to4 I__7713 (
            .O(N__40865),
            .I(N__40840));
    Span4Mux_v I__7712 (
            .O(N__40858),
            .I(N__40837));
    Span4Mux_h I__7711 (
            .O(N__40855),
            .I(N__40834));
    Span4Mux_h I__7710 (
            .O(N__40852),
            .I(N__40829));
    Span4Mux_v I__7709 (
            .O(N__40849),
            .I(N__40829));
    Span4Mux_v I__7708 (
            .O(N__40846),
            .I(N__40826));
    Sp12to4 I__7707 (
            .O(N__40843),
            .I(N__40821));
    Span12Mux_v I__7706 (
            .O(N__40840),
            .I(N__40821));
    Span4Mux_v I__7705 (
            .O(N__40837),
            .I(N__40818));
    Odrv4 I__7704 (
            .O(N__40834),
            .I(\c0.n8107 ));
    Odrv4 I__7703 (
            .O(N__40829),
            .I(\c0.n8107 ));
    Odrv4 I__7702 (
            .O(N__40826),
            .I(\c0.n8107 ));
    Odrv12 I__7701 (
            .O(N__40821),
            .I(\c0.n8107 ));
    Odrv4 I__7700 (
            .O(N__40818),
            .I(\c0.n8107 ));
    InMux I__7699 (
            .O(N__40807),
            .I(N__40804));
    LocalMux I__7698 (
            .O(N__40804),
            .I(N__40801));
    Odrv4 I__7697 (
            .O(N__40801),
            .I(\c0.n49 ));
    CascadeMux I__7696 (
            .O(N__40798),
            .I(N__40795));
    InMux I__7695 (
            .O(N__40795),
            .I(N__40792));
    LocalMux I__7694 (
            .O(N__40792),
            .I(N__40789));
    Span4Mux_v I__7693 (
            .O(N__40789),
            .I(N__40786));
    Odrv4 I__7692 (
            .O(N__40786),
            .I(\c0.n50 ));
    InMux I__7691 (
            .O(N__40783),
            .I(N__40780));
    LocalMux I__7690 (
            .O(N__40780),
            .I(\c0.n54 ));
    SRMux I__7689 (
            .O(N__40777),
            .I(N__40770));
    InMux I__7688 (
            .O(N__40776),
            .I(N__40770));
    InMux I__7687 (
            .O(N__40775),
            .I(N__40767));
    LocalMux I__7686 (
            .O(N__40770),
            .I(N__40764));
    LocalMux I__7685 (
            .O(N__40767),
            .I(N__40761));
    Span12Mux_v I__7684 (
            .O(N__40764),
            .I(N__40758));
    Span4Mux_v I__7683 (
            .O(N__40761),
            .I(N__40755));
    Odrv12 I__7682 (
            .O(N__40758),
            .I(\c0.n22665 ));
    Odrv4 I__7681 (
            .O(N__40755),
            .I(\c0.n22665 ));
    CascadeMux I__7680 (
            .O(N__40750),
            .I(N__40746));
    InMux I__7679 (
            .O(N__40749),
            .I(N__40741));
    InMux I__7678 (
            .O(N__40746),
            .I(N__40738));
    InMux I__7677 (
            .O(N__40745),
            .I(N__40735));
    CascadeMux I__7676 (
            .O(N__40744),
            .I(N__40731));
    LocalMux I__7675 (
            .O(N__40741),
            .I(N__40728));
    LocalMux I__7674 (
            .O(N__40738),
            .I(N__40725));
    LocalMux I__7673 (
            .O(N__40735),
            .I(N__40722));
    InMux I__7672 (
            .O(N__40734),
            .I(N__40717));
    InMux I__7671 (
            .O(N__40731),
            .I(N__40717));
    Span4Mux_v I__7670 (
            .O(N__40728),
            .I(N__40714));
    Odrv4 I__7669 (
            .O(N__40725),
            .I(\c0.n3239 ));
    Odrv4 I__7668 (
            .O(N__40722),
            .I(\c0.n3239 ));
    LocalMux I__7667 (
            .O(N__40717),
            .I(\c0.n3239 ));
    Odrv4 I__7666 (
            .O(N__40714),
            .I(\c0.n3239 ));
    CascadeMux I__7665 (
            .O(N__40705),
            .I(\c0.n63_adj_4293_cascade_ ));
    InMux I__7664 (
            .O(N__40702),
            .I(N__40698));
    InMux I__7663 (
            .O(N__40701),
            .I(N__40695));
    LocalMux I__7662 (
            .O(N__40698),
            .I(N__40690));
    LocalMux I__7661 (
            .O(N__40695),
            .I(N__40690));
    Odrv4 I__7660 (
            .O(N__40690),
            .I(\c0.n13020 ));
    InMux I__7659 (
            .O(N__40687),
            .I(N__40684));
    LocalMux I__7658 (
            .O(N__40684),
            .I(N__40681));
    Span4Mux_h I__7657 (
            .O(N__40681),
            .I(N__40678));
    Odrv4 I__7656 (
            .O(N__40678),
            .I(\c0.n4_adj_4345 ));
    CascadeMux I__7655 (
            .O(N__40675),
            .I(\c0.n84_cascade_ ));
    InMux I__7654 (
            .O(N__40672),
            .I(N__40667));
    InMux I__7653 (
            .O(N__40671),
            .I(N__40662));
    InMux I__7652 (
            .O(N__40670),
            .I(N__40662));
    LocalMux I__7651 (
            .O(N__40667),
            .I(\c0.n12990 ));
    LocalMux I__7650 (
            .O(N__40662),
            .I(\c0.n12990 ));
    InMux I__7649 (
            .O(N__40657),
            .I(N__40654));
    LocalMux I__7648 (
            .O(N__40654),
            .I(N__40649));
    InMux I__7647 (
            .O(N__40653),
            .I(N__40644));
    InMux I__7646 (
            .O(N__40652),
            .I(N__40644));
    Span12Mux_v I__7645 (
            .O(N__40649),
            .I(N__40641));
    LocalMux I__7644 (
            .O(N__40644),
            .I(N__40638));
    Odrv12 I__7643 (
            .O(N__40641),
            .I(\c0.n7_adj_4344 ));
    Odrv4 I__7642 (
            .O(N__40638),
            .I(\c0.n7_adj_4344 ));
    InMux I__7641 (
            .O(N__40633),
            .I(N__40630));
    LocalMux I__7640 (
            .O(N__40630),
            .I(N__40625));
    InMux I__7639 (
            .O(N__40629),
            .I(N__40618));
    InMux I__7638 (
            .O(N__40628),
            .I(N__40618));
    Span4Mux_v I__7637 (
            .O(N__40625),
            .I(N__40615));
    InMux I__7636 (
            .O(N__40624),
            .I(N__40610));
    InMux I__7635 (
            .O(N__40623),
            .I(N__40610));
    LocalMux I__7634 (
            .O(N__40618),
            .I(N__40607));
    Odrv4 I__7633 (
            .O(N__40615),
            .I(\c0.n12967 ));
    LocalMux I__7632 (
            .O(N__40610),
            .I(\c0.n12967 ));
    Odrv4 I__7631 (
            .O(N__40607),
            .I(\c0.n12967 ));
    InMux I__7630 (
            .O(N__40600),
            .I(N__40592));
    InMux I__7629 (
            .O(N__40599),
            .I(N__40589));
    CascadeMux I__7628 (
            .O(N__40598),
            .I(N__40586));
    CascadeMux I__7627 (
            .O(N__40597),
            .I(N__40582));
    InMux I__7626 (
            .O(N__40596),
            .I(N__40577));
    InMux I__7625 (
            .O(N__40595),
            .I(N__40577));
    LocalMux I__7624 (
            .O(N__40592),
            .I(N__40572));
    LocalMux I__7623 (
            .O(N__40589),
            .I(N__40569));
    InMux I__7622 (
            .O(N__40586),
            .I(N__40562));
    InMux I__7621 (
            .O(N__40585),
            .I(N__40562));
    InMux I__7620 (
            .O(N__40582),
            .I(N__40562));
    LocalMux I__7619 (
            .O(N__40577),
            .I(N__40559));
    InMux I__7618 (
            .O(N__40576),
            .I(N__40556));
    InMux I__7617 (
            .O(N__40575),
            .I(N__40553));
    Odrv12 I__7616 (
            .O(N__40572),
            .I(\c0.FRAME_MATCHER_state_0 ));
    Odrv4 I__7615 (
            .O(N__40569),
            .I(\c0.FRAME_MATCHER_state_0 ));
    LocalMux I__7614 (
            .O(N__40562),
            .I(\c0.FRAME_MATCHER_state_0 ));
    Odrv4 I__7613 (
            .O(N__40559),
            .I(\c0.FRAME_MATCHER_state_0 ));
    LocalMux I__7612 (
            .O(N__40556),
            .I(\c0.FRAME_MATCHER_state_0 ));
    LocalMux I__7611 (
            .O(N__40553),
            .I(\c0.FRAME_MATCHER_state_0 ));
    CascadeMux I__7610 (
            .O(N__40540),
            .I(N__40536));
    InMux I__7609 (
            .O(N__40539),
            .I(N__40528));
    InMux I__7608 (
            .O(N__40536),
            .I(N__40528));
    InMux I__7607 (
            .O(N__40535),
            .I(N__40528));
    LocalMux I__7606 (
            .O(N__40528),
            .I(N__40524));
    InMux I__7605 (
            .O(N__40527),
            .I(N__40521));
    Span4Mux_h I__7604 (
            .O(N__40524),
            .I(N__40516));
    LocalMux I__7603 (
            .O(N__40521),
            .I(N__40516));
    Odrv4 I__7602 (
            .O(N__40516),
            .I(\c0.n12996 ));
    InMux I__7601 (
            .O(N__40513),
            .I(N__40509));
    CascadeMux I__7600 (
            .O(N__40512),
            .I(N__40506));
    LocalMux I__7599 (
            .O(N__40509),
            .I(N__40502));
    InMux I__7598 (
            .O(N__40506),
            .I(N__40497));
    InMux I__7597 (
            .O(N__40505),
            .I(N__40497));
    Odrv4 I__7596 (
            .O(N__40502),
            .I(\c0.n4_adj_4419 ));
    LocalMux I__7595 (
            .O(N__40497),
            .I(\c0.n4_adj_4419 ));
    CascadeMux I__7594 (
            .O(N__40492),
            .I(\c0.data_out_frame_0__7__N_2568_cascade_ ));
    CascadeMux I__7593 (
            .O(N__40489),
            .I(\c0.n1220_cascade_ ));
    InMux I__7592 (
            .O(N__40486),
            .I(N__40483));
    LocalMux I__7591 (
            .O(N__40483),
            .I(N__40480));
    Span12Mux_v I__7590 (
            .O(N__40480),
            .I(N__40477));
    Odrv12 I__7589 (
            .O(N__40477),
            .I(\c0.n4_adj_4373 ));
    CascadeMux I__7588 (
            .O(N__40474),
            .I(\c0.n5024_cascade_ ));
    InMux I__7587 (
            .O(N__40471),
            .I(N__40468));
    LocalMux I__7586 (
            .O(N__40468),
            .I(N__40465));
    Span4Mux_h I__7585 (
            .O(N__40465),
            .I(N__40462));
    Odrv4 I__7584 (
            .O(N__40462),
            .I(\c0.n21773 ));
    CascadeMux I__7583 (
            .O(N__40459),
            .I(\c0.n21773_cascade_ ));
    InMux I__7582 (
            .O(N__40456),
            .I(N__40448));
    InMux I__7581 (
            .O(N__40455),
            .I(N__40448));
    InMux I__7580 (
            .O(N__40454),
            .I(N__40440));
    InMux I__7579 (
            .O(N__40453),
            .I(N__40440));
    LocalMux I__7578 (
            .O(N__40448),
            .I(N__40437));
    InMux I__7577 (
            .O(N__40447),
            .I(N__40430));
    InMux I__7576 (
            .O(N__40446),
            .I(N__40430));
    InMux I__7575 (
            .O(N__40445),
            .I(N__40430));
    LocalMux I__7574 (
            .O(N__40440),
            .I(\c0.data_out_frame_29_7_N_1483_1 ));
    Odrv4 I__7573 (
            .O(N__40437),
            .I(\c0.data_out_frame_29_7_N_1483_1 ));
    LocalMux I__7572 (
            .O(N__40430),
            .I(\c0.data_out_frame_29_7_N_1483_1 ));
    CascadeMux I__7571 (
            .O(N__40423),
            .I(\c0.n4_adj_4328_cascade_ ));
    InMux I__7570 (
            .O(N__40420),
            .I(N__40415));
    InMux I__7569 (
            .O(N__40419),
            .I(N__40412));
    InMux I__7568 (
            .O(N__40418),
            .I(N__40409));
    LocalMux I__7567 (
            .O(N__40415),
            .I(\c0.data_out_frame_0__7__N_2568 ));
    LocalMux I__7566 (
            .O(N__40412),
            .I(\c0.data_out_frame_0__7__N_2568 ));
    LocalMux I__7565 (
            .O(N__40409),
            .I(\c0.data_out_frame_0__7__N_2568 ));
    InMux I__7564 (
            .O(N__40402),
            .I(N__40396));
    InMux I__7563 (
            .O(N__40401),
            .I(N__40396));
    LocalMux I__7562 (
            .O(N__40396),
            .I(\c0.FRAME_MATCHER_state_1 ));
    InMux I__7561 (
            .O(N__40393),
            .I(N__40390));
    LocalMux I__7560 (
            .O(N__40390),
            .I(N__40387));
    Span4Mux_h I__7559 (
            .O(N__40387),
            .I(N__40384));
    Odrv4 I__7558 (
            .O(N__40384),
            .I(\c0.n4_adj_4391 ));
    CascadeMux I__7557 (
            .O(N__40381),
            .I(N__40378));
    InMux I__7556 (
            .O(N__40378),
            .I(N__40375));
    LocalMux I__7555 (
            .O(N__40375),
            .I(N__40372));
    Odrv12 I__7554 (
            .O(N__40372),
            .I(\c0.n38_adj_4390 ));
    InMux I__7553 (
            .O(N__40369),
            .I(N__40363));
    InMux I__7552 (
            .O(N__40368),
            .I(N__40360));
    CascadeMux I__7551 (
            .O(N__40367),
            .I(N__40356));
    CascadeMux I__7550 (
            .O(N__40366),
            .I(N__40352));
    LocalMux I__7549 (
            .O(N__40363),
            .I(N__40349));
    LocalMux I__7548 (
            .O(N__40360),
            .I(N__40346));
    InMux I__7547 (
            .O(N__40359),
            .I(N__40343));
    InMux I__7546 (
            .O(N__40356),
            .I(N__40340));
    InMux I__7545 (
            .O(N__40355),
            .I(N__40337));
    InMux I__7544 (
            .O(N__40352),
            .I(N__40334));
    Span4Mux_v I__7543 (
            .O(N__40349),
            .I(N__40331));
    Span4Mux_h I__7542 (
            .O(N__40346),
            .I(N__40328));
    LocalMux I__7541 (
            .O(N__40343),
            .I(N__40325));
    LocalMux I__7540 (
            .O(N__40340),
            .I(encoder0_position_23));
    LocalMux I__7539 (
            .O(N__40337),
            .I(encoder0_position_23));
    LocalMux I__7538 (
            .O(N__40334),
            .I(encoder0_position_23));
    Odrv4 I__7537 (
            .O(N__40331),
            .I(encoder0_position_23));
    Odrv4 I__7536 (
            .O(N__40328),
            .I(encoder0_position_23));
    Odrv12 I__7535 (
            .O(N__40325),
            .I(encoder0_position_23));
    CascadeMux I__7534 (
            .O(N__40312),
            .I(N__40309));
    InMux I__7533 (
            .O(N__40309),
            .I(N__40306));
    LocalMux I__7532 (
            .O(N__40306),
            .I(N__40301));
    InMux I__7531 (
            .O(N__40305),
            .I(N__40298));
    InMux I__7530 (
            .O(N__40304),
            .I(N__40295));
    Span4Mux_h I__7529 (
            .O(N__40301),
            .I(N__40291));
    LocalMux I__7528 (
            .O(N__40298),
            .I(N__40288));
    LocalMux I__7527 (
            .O(N__40295),
            .I(N__40285));
    CascadeMux I__7526 (
            .O(N__40294),
            .I(N__40281));
    Span4Mux_h I__7525 (
            .O(N__40291),
            .I(N__40276));
    Span4Mux_h I__7524 (
            .O(N__40288),
            .I(N__40276));
    Span4Mux_v I__7523 (
            .O(N__40285),
            .I(N__40273));
    InMux I__7522 (
            .O(N__40284),
            .I(N__40268));
    InMux I__7521 (
            .O(N__40281),
            .I(N__40268));
    Odrv4 I__7520 (
            .O(N__40276),
            .I(encoder0_position_8));
    Odrv4 I__7519 (
            .O(N__40273),
            .I(encoder0_position_8));
    LocalMux I__7518 (
            .O(N__40268),
            .I(encoder0_position_8));
    InMux I__7517 (
            .O(N__40261),
            .I(N__40258));
    LocalMux I__7516 (
            .O(N__40258),
            .I(N__40254));
    InMux I__7515 (
            .O(N__40257),
            .I(N__40251));
    Span4Mux_v I__7514 (
            .O(N__40254),
            .I(N__40246));
    LocalMux I__7513 (
            .O(N__40251),
            .I(N__40246));
    Odrv4 I__7512 (
            .O(N__40246),
            .I(\c0.n22032 ));
    InMux I__7511 (
            .O(N__40243),
            .I(N__40238));
    InMux I__7510 (
            .O(N__40242),
            .I(N__40233));
    InMux I__7509 (
            .O(N__40241),
            .I(N__40233));
    LocalMux I__7508 (
            .O(N__40238),
            .I(N__40229));
    LocalMux I__7507 (
            .O(N__40233),
            .I(N__40226));
    InMux I__7506 (
            .O(N__40232),
            .I(N__40223));
    Span4Mux_v I__7505 (
            .O(N__40229),
            .I(N__40218));
    Span4Mux_h I__7504 (
            .O(N__40226),
            .I(N__40218));
    LocalMux I__7503 (
            .O(N__40223),
            .I(data_in_3_0));
    Odrv4 I__7502 (
            .O(N__40218),
            .I(data_in_3_0));
    InMux I__7501 (
            .O(N__40213),
            .I(N__40210));
    LocalMux I__7500 (
            .O(N__40210),
            .I(N__40205));
    InMux I__7499 (
            .O(N__40209),
            .I(N__40202));
    InMux I__7498 (
            .O(N__40208),
            .I(N__40199));
    Span4Mux_v I__7497 (
            .O(N__40205),
            .I(N__40195));
    LocalMux I__7496 (
            .O(N__40202),
            .I(N__40192));
    LocalMux I__7495 (
            .O(N__40199),
            .I(N__40189));
    InMux I__7494 (
            .O(N__40198),
            .I(N__40186));
    Span4Mux_h I__7493 (
            .O(N__40195),
            .I(N__40179));
    Span4Mux_v I__7492 (
            .O(N__40192),
            .I(N__40179));
    Span4Mux_v I__7491 (
            .O(N__40189),
            .I(N__40179));
    LocalMux I__7490 (
            .O(N__40186),
            .I(control_mode_5));
    Odrv4 I__7489 (
            .O(N__40179),
            .I(control_mode_5));
    CascadeMux I__7488 (
            .O(N__40174),
            .I(\c0.n23215_cascade_ ));
    InMux I__7487 (
            .O(N__40171),
            .I(N__40166));
    InMux I__7486 (
            .O(N__40170),
            .I(N__40163));
    InMux I__7485 (
            .O(N__40169),
            .I(N__40160));
    LocalMux I__7484 (
            .O(N__40166),
            .I(N__40154));
    LocalMux I__7483 (
            .O(N__40163),
            .I(N__40151));
    LocalMux I__7482 (
            .O(N__40160),
            .I(N__40146));
    InMux I__7481 (
            .O(N__40159),
            .I(N__40143));
    InMux I__7480 (
            .O(N__40158),
            .I(N__40138));
    InMux I__7479 (
            .O(N__40157),
            .I(N__40138));
    Span4Mux_v I__7478 (
            .O(N__40154),
            .I(N__40133));
    Span4Mux_h I__7477 (
            .O(N__40151),
            .I(N__40133));
    InMux I__7476 (
            .O(N__40150),
            .I(N__40128));
    InMux I__7475 (
            .O(N__40149),
            .I(N__40128));
    Span4Mux_h I__7474 (
            .O(N__40146),
            .I(N__40125));
    LocalMux I__7473 (
            .O(N__40143),
            .I(N__40120));
    LocalMux I__7472 (
            .O(N__40138),
            .I(N__40120));
    Span4Mux_h I__7471 (
            .O(N__40133),
            .I(N__40115));
    LocalMux I__7470 (
            .O(N__40128),
            .I(N__40115));
    Span4Mux_h I__7469 (
            .O(N__40125),
            .I(N__40110));
    Span4Mux_v I__7468 (
            .O(N__40120),
            .I(N__40107));
    Span4Mux_h I__7467 (
            .O(N__40115),
            .I(N__40104));
    InMux I__7466 (
            .O(N__40114),
            .I(N__40099));
    InMux I__7465 (
            .O(N__40113),
            .I(N__40099));
    Odrv4 I__7464 (
            .O(N__40110),
            .I(data_out_frame_29_7_N_1483_2));
    Odrv4 I__7463 (
            .O(N__40107),
            .I(data_out_frame_29_7_N_1483_2));
    Odrv4 I__7462 (
            .O(N__40104),
            .I(data_out_frame_29_7_N_1483_2));
    LocalMux I__7461 (
            .O(N__40099),
            .I(data_out_frame_29_7_N_1483_2));
    InMux I__7460 (
            .O(N__40090),
            .I(N__40087));
    LocalMux I__7459 (
            .O(N__40087),
            .I(\c0.n6_adj_4338 ));
    CascadeMux I__7458 (
            .O(N__40084),
            .I(\c0.n17602_cascade_ ));
    InMux I__7457 (
            .O(N__40081),
            .I(N__40078));
    LocalMux I__7456 (
            .O(N__40078),
            .I(\c0.n8_adj_4417 ));
    InMux I__7455 (
            .O(N__40075),
            .I(N__40072));
    LocalMux I__7454 (
            .O(N__40072),
            .I(N__40069));
    Span4Mux_h I__7453 (
            .O(N__40069),
            .I(N__40066));
    Odrv4 I__7452 (
            .O(N__40066),
            .I(n2245));
    InMux I__7451 (
            .O(N__40063),
            .I(N__40060));
    LocalMux I__7450 (
            .O(N__40060),
            .I(N__40053));
    InMux I__7449 (
            .O(N__40059),
            .I(N__40050));
    InMux I__7448 (
            .O(N__40058),
            .I(N__40047));
    InMux I__7447 (
            .O(N__40057),
            .I(N__40044));
    InMux I__7446 (
            .O(N__40056),
            .I(N__40041));
    Span4Mux_v I__7445 (
            .O(N__40053),
            .I(N__40036));
    LocalMux I__7444 (
            .O(N__40050),
            .I(N__40033));
    LocalMux I__7443 (
            .O(N__40047),
            .I(N__40028));
    LocalMux I__7442 (
            .O(N__40044),
            .I(N__40028));
    LocalMux I__7441 (
            .O(N__40041),
            .I(N__40025));
    InMux I__7440 (
            .O(N__40040),
            .I(N__40022));
    InMux I__7439 (
            .O(N__40039),
            .I(N__40019));
    Span4Mux_h I__7438 (
            .O(N__40036),
            .I(N__40014));
    Span4Mux_v I__7437 (
            .O(N__40033),
            .I(N__40014));
    Span4Mux_v I__7436 (
            .O(N__40028),
            .I(N__40011));
    Span12Mux_h I__7435 (
            .O(N__40025),
            .I(N__40008));
    LocalMux I__7434 (
            .O(N__40022),
            .I(N__40005));
    LocalMux I__7433 (
            .O(N__40019),
            .I(encoder0_position_26));
    Odrv4 I__7432 (
            .O(N__40014),
            .I(encoder0_position_26));
    Odrv4 I__7431 (
            .O(N__40011),
            .I(encoder0_position_26));
    Odrv12 I__7430 (
            .O(N__40008),
            .I(encoder0_position_26));
    Odrv4 I__7429 (
            .O(N__40005),
            .I(encoder0_position_26));
    InMux I__7428 (
            .O(N__39994),
            .I(N__39991));
    LocalMux I__7427 (
            .O(N__39991),
            .I(N__39988));
    Span4Mux_v I__7426 (
            .O(N__39988),
            .I(N__39985));
    Sp12to4 I__7425 (
            .O(N__39985),
            .I(N__39982));
    Odrv12 I__7424 (
            .O(N__39982),
            .I(n2263));
    CascadeMux I__7423 (
            .O(N__39979),
            .I(N__39976));
    InMux I__7422 (
            .O(N__39976),
            .I(N__39971));
    InMux I__7421 (
            .O(N__39975),
            .I(N__39968));
    InMux I__7420 (
            .O(N__39974),
            .I(N__39963));
    LocalMux I__7419 (
            .O(N__39971),
            .I(N__39960));
    LocalMux I__7418 (
            .O(N__39968),
            .I(N__39957));
    InMux I__7417 (
            .O(N__39967),
            .I(N__39952));
    InMux I__7416 (
            .O(N__39966),
            .I(N__39952));
    LocalMux I__7415 (
            .O(N__39963),
            .I(encoder0_position_10));
    Odrv12 I__7414 (
            .O(N__39960),
            .I(encoder0_position_10));
    Odrv4 I__7413 (
            .O(N__39957),
            .I(encoder0_position_10));
    LocalMux I__7412 (
            .O(N__39952),
            .I(encoder0_position_10));
    CascadeMux I__7411 (
            .O(N__39943),
            .I(N__39940));
    InMux I__7410 (
            .O(N__39940),
            .I(N__39937));
    LocalMux I__7409 (
            .O(N__39937),
            .I(N__39934));
    Span4Mux_h I__7408 (
            .O(N__39934),
            .I(N__39930));
    InMux I__7407 (
            .O(N__39933),
            .I(N__39927));
    Span4Mux_h I__7406 (
            .O(N__39930),
            .I(N__39924));
    LocalMux I__7405 (
            .O(N__39927),
            .I(data_out_frame_8_2));
    Odrv4 I__7404 (
            .O(N__39924),
            .I(data_out_frame_8_2));
    InMux I__7403 (
            .O(N__39919),
            .I(N__39916));
    LocalMux I__7402 (
            .O(N__39916),
            .I(N__39913));
    Span4Mux_h I__7401 (
            .O(N__39913),
            .I(N__39910));
    Odrv4 I__7400 (
            .O(N__39910),
            .I(n2246));
    CascadeMux I__7399 (
            .O(N__39907),
            .I(N__39904));
    InMux I__7398 (
            .O(N__39904),
            .I(N__39899));
    InMux I__7397 (
            .O(N__39903),
            .I(N__39895));
    CascadeMux I__7396 (
            .O(N__39902),
            .I(N__39890));
    LocalMux I__7395 (
            .O(N__39899),
            .I(N__39886));
    InMux I__7394 (
            .O(N__39898),
            .I(N__39883));
    LocalMux I__7393 (
            .O(N__39895),
            .I(N__39880));
    InMux I__7392 (
            .O(N__39894),
            .I(N__39875));
    InMux I__7391 (
            .O(N__39893),
            .I(N__39875));
    InMux I__7390 (
            .O(N__39890),
            .I(N__39872));
    InMux I__7389 (
            .O(N__39889),
            .I(N__39869));
    Span4Mux_h I__7388 (
            .O(N__39886),
            .I(N__39866));
    LocalMux I__7387 (
            .O(N__39883),
            .I(N__39863));
    Span4Mux_v I__7386 (
            .O(N__39880),
            .I(N__39858));
    LocalMux I__7385 (
            .O(N__39875),
            .I(N__39858));
    LocalMux I__7384 (
            .O(N__39872),
            .I(encoder0_position_25));
    LocalMux I__7383 (
            .O(N__39869),
            .I(encoder0_position_25));
    Odrv4 I__7382 (
            .O(N__39866),
            .I(encoder0_position_25));
    Odrv12 I__7381 (
            .O(N__39863),
            .I(encoder0_position_25));
    Odrv4 I__7380 (
            .O(N__39858),
            .I(encoder0_position_25));
    InMux I__7379 (
            .O(N__39847),
            .I(N__39841));
    InMux I__7378 (
            .O(N__39846),
            .I(N__39841));
    LocalMux I__7377 (
            .O(N__39841),
            .I(data_out_frame_7_6));
    InMux I__7376 (
            .O(N__39838),
            .I(N__39829));
    InMux I__7375 (
            .O(N__39837),
            .I(N__39826));
    InMux I__7374 (
            .O(N__39836),
            .I(N__39823));
    InMux I__7373 (
            .O(N__39835),
            .I(N__39819));
    InMux I__7372 (
            .O(N__39834),
            .I(N__39811));
    InMux I__7371 (
            .O(N__39833),
            .I(N__39808));
    InMux I__7370 (
            .O(N__39832),
            .I(N__39801));
    LocalMux I__7369 (
            .O(N__39829),
            .I(N__39796));
    LocalMux I__7368 (
            .O(N__39826),
            .I(N__39791));
    LocalMux I__7367 (
            .O(N__39823),
            .I(N__39791));
    InMux I__7366 (
            .O(N__39822),
            .I(N__39788));
    LocalMux I__7365 (
            .O(N__39819),
            .I(N__39785));
    InMux I__7364 (
            .O(N__39818),
            .I(N__39782));
    InMux I__7363 (
            .O(N__39817),
            .I(N__39768));
    InMux I__7362 (
            .O(N__39816),
            .I(N__39763));
    InMux I__7361 (
            .O(N__39815),
            .I(N__39763));
    InMux I__7360 (
            .O(N__39814),
            .I(N__39760));
    LocalMux I__7359 (
            .O(N__39811),
            .I(N__39751));
    LocalMux I__7358 (
            .O(N__39808),
            .I(N__39751));
    InMux I__7357 (
            .O(N__39807),
            .I(N__39744));
    InMux I__7356 (
            .O(N__39806),
            .I(N__39744));
    InMux I__7355 (
            .O(N__39805),
            .I(N__39741));
    InMux I__7354 (
            .O(N__39804),
            .I(N__39738));
    LocalMux I__7353 (
            .O(N__39801),
            .I(N__39735));
    InMux I__7352 (
            .O(N__39800),
            .I(N__39727));
    InMux I__7351 (
            .O(N__39799),
            .I(N__39727));
    Span4Mux_v I__7350 (
            .O(N__39796),
            .I(N__39721));
    Span4Mux_v I__7349 (
            .O(N__39791),
            .I(N__39721));
    LocalMux I__7348 (
            .O(N__39788),
            .I(N__39715));
    Span4Mux_h I__7347 (
            .O(N__39785),
            .I(N__39715));
    LocalMux I__7346 (
            .O(N__39782),
            .I(N__39712));
    InMux I__7345 (
            .O(N__39781),
            .I(N__39709));
    InMux I__7344 (
            .O(N__39780),
            .I(N__39702));
    InMux I__7343 (
            .O(N__39779),
            .I(N__39702));
    InMux I__7342 (
            .O(N__39778),
            .I(N__39702));
    InMux I__7341 (
            .O(N__39777),
            .I(N__39697));
    InMux I__7340 (
            .O(N__39776),
            .I(N__39690));
    InMux I__7339 (
            .O(N__39775),
            .I(N__39690));
    InMux I__7338 (
            .O(N__39774),
            .I(N__39690));
    InMux I__7337 (
            .O(N__39773),
            .I(N__39687));
    InMux I__7336 (
            .O(N__39772),
            .I(N__39682));
    InMux I__7335 (
            .O(N__39771),
            .I(N__39682));
    LocalMux I__7334 (
            .O(N__39768),
            .I(N__39679));
    LocalMux I__7333 (
            .O(N__39763),
            .I(N__39676));
    LocalMux I__7332 (
            .O(N__39760),
            .I(N__39673));
    InMux I__7331 (
            .O(N__39759),
            .I(N__39668));
    InMux I__7330 (
            .O(N__39758),
            .I(N__39668));
    InMux I__7329 (
            .O(N__39757),
            .I(N__39663));
    InMux I__7328 (
            .O(N__39756),
            .I(N__39663));
    Span4Mux_v I__7327 (
            .O(N__39751),
            .I(N__39660));
    InMux I__7326 (
            .O(N__39750),
            .I(N__39655));
    InMux I__7325 (
            .O(N__39749),
            .I(N__39655));
    LocalMux I__7324 (
            .O(N__39744),
            .I(N__39650));
    LocalMux I__7323 (
            .O(N__39741),
            .I(N__39650));
    LocalMux I__7322 (
            .O(N__39738),
            .I(N__39647));
    Span4Mux_h I__7321 (
            .O(N__39735),
            .I(N__39644));
    InMux I__7320 (
            .O(N__39734),
            .I(N__39639));
    InMux I__7319 (
            .O(N__39733),
            .I(N__39639));
    InMux I__7318 (
            .O(N__39732),
            .I(N__39636));
    LocalMux I__7317 (
            .O(N__39727),
            .I(N__39633));
    InMux I__7316 (
            .O(N__39726),
            .I(N__39630));
    Sp12to4 I__7315 (
            .O(N__39721),
            .I(N__39627));
    CascadeMux I__7314 (
            .O(N__39720),
            .I(N__39623));
    Span4Mux_v I__7313 (
            .O(N__39715),
            .I(N__39616));
    Span4Mux_h I__7312 (
            .O(N__39712),
            .I(N__39616));
    LocalMux I__7311 (
            .O(N__39709),
            .I(N__39616));
    LocalMux I__7310 (
            .O(N__39702),
            .I(N__39613));
    InMux I__7309 (
            .O(N__39701),
            .I(N__39608));
    InMux I__7308 (
            .O(N__39700),
            .I(N__39608));
    LocalMux I__7307 (
            .O(N__39697),
            .I(N__39603));
    LocalMux I__7306 (
            .O(N__39690),
            .I(N__39603));
    LocalMux I__7305 (
            .O(N__39687),
            .I(N__39598));
    LocalMux I__7304 (
            .O(N__39682),
            .I(N__39598));
    Span4Mux_v I__7303 (
            .O(N__39679),
            .I(N__39591));
    Span4Mux_v I__7302 (
            .O(N__39676),
            .I(N__39591));
    Span4Mux_v I__7301 (
            .O(N__39673),
            .I(N__39591));
    LocalMux I__7300 (
            .O(N__39668),
            .I(N__39586));
    LocalMux I__7299 (
            .O(N__39663),
            .I(N__39586));
    Span4Mux_h I__7298 (
            .O(N__39660),
            .I(N__39583));
    LocalMux I__7297 (
            .O(N__39655),
            .I(N__39574));
    Span4Mux_v I__7296 (
            .O(N__39650),
            .I(N__39574));
    Span4Mux_v I__7295 (
            .O(N__39647),
            .I(N__39574));
    Span4Mux_h I__7294 (
            .O(N__39644),
            .I(N__39574));
    LocalMux I__7293 (
            .O(N__39639),
            .I(N__39569));
    LocalMux I__7292 (
            .O(N__39636),
            .I(N__39569));
    Span4Mux_v I__7291 (
            .O(N__39633),
            .I(N__39564));
    LocalMux I__7290 (
            .O(N__39630),
            .I(N__39564));
    Span12Mux_h I__7289 (
            .O(N__39627),
            .I(N__39561));
    InMux I__7288 (
            .O(N__39626),
            .I(N__39558));
    InMux I__7287 (
            .O(N__39623),
            .I(N__39555));
    Span4Mux_h I__7286 (
            .O(N__39616),
            .I(N__39552));
    Span4Mux_v I__7285 (
            .O(N__39613),
            .I(N__39541));
    LocalMux I__7284 (
            .O(N__39608),
            .I(N__39541));
    Span4Mux_v I__7283 (
            .O(N__39603),
            .I(N__39541));
    Span4Mux_v I__7282 (
            .O(N__39598),
            .I(N__39541));
    Span4Mux_h I__7281 (
            .O(N__39591),
            .I(N__39541));
    Span4Mux_h I__7280 (
            .O(N__39586),
            .I(N__39534));
    Span4Mux_v I__7279 (
            .O(N__39583),
            .I(N__39534));
    Span4Mux_h I__7278 (
            .O(N__39574),
            .I(N__39534));
    Span12Mux_v I__7277 (
            .O(N__39569),
            .I(N__39525));
    Sp12to4 I__7276 (
            .O(N__39564),
            .I(N__39525));
    Span12Mux_v I__7275 (
            .O(N__39561),
            .I(N__39525));
    LocalMux I__7274 (
            .O(N__39558),
            .I(N__39525));
    LocalMux I__7273 (
            .O(N__39555),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__7272 (
            .O(N__39552),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__7271 (
            .O(N__39541),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__7270 (
            .O(N__39534),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv12 I__7269 (
            .O(N__39525),
            .I(\c0.byte_transmit_counter_0 ));
    InMux I__7268 (
            .O(N__39514),
            .I(N__39511));
    LocalMux I__7267 (
            .O(N__39511),
            .I(N__39508));
    Span4Mux_v I__7266 (
            .O(N__39508),
            .I(N__39505));
    Span4Mux_h I__7265 (
            .O(N__39505),
            .I(N__39502));
    Odrv4 I__7264 (
            .O(N__39502),
            .I(\c0.n5_adj_4350 ));
    InMux I__7263 (
            .O(N__39499),
            .I(N__39496));
    LocalMux I__7262 (
            .O(N__39496),
            .I(N__39492));
    InMux I__7261 (
            .O(N__39495),
            .I(N__39489));
    Span4Mux_v I__7260 (
            .O(N__39492),
            .I(N__39481));
    LocalMux I__7259 (
            .O(N__39489),
            .I(N__39481));
    InMux I__7258 (
            .O(N__39488),
            .I(N__39478));
    InMux I__7257 (
            .O(N__39487),
            .I(N__39472));
    InMux I__7256 (
            .O(N__39486),
            .I(N__39469));
    Span4Mux_h I__7255 (
            .O(N__39481),
            .I(N__39466));
    LocalMux I__7254 (
            .O(N__39478),
            .I(N__39463));
    InMux I__7253 (
            .O(N__39477),
            .I(N__39458));
    InMux I__7252 (
            .O(N__39476),
            .I(N__39458));
    InMux I__7251 (
            .O(N__39475),
            .I(N__39455));
    LocalMux I__7250 (
            .O(N__39472),
            .I(N__39452));
    LocalMux I__7249 (
            .O(N__39469),
            .I(N__39447));
    Span4Mux_v I__7248 (
            .O(N__39466),
            .I(N__39447));
    Span12Mux_h I__7247 (
            .O(N__39463),
            .I(N__39440));
    LocalMux I__7246 (
            .O(N__39458),
            .I(N__39440));
    LocalMux I__7245 (
            .O(N__39455),
            .I(N__39440));
    Odrv12 I__7244 (
            .O(N__39452),
            .I(control_mode_2));
    Odrv4 I__7243 (
            .O(N__39447),
            .I(control_mode_2));
    Odrv12 I__7242 (
            .O(N__39440),
            .I(control_mode_2));
    CascadeMux I__7241 (
            .O(N__39433),
            .I(\c0.n6_adj_4315_cascade_ ));
    InMux I__7240 (
            .O(N__39430),
            .I(N__39427));
    LocalMux I__7239 (
            .O(N__39427),
            .I(N__39423));
    InMux I__7238 (
            .O(N__39426),
            .I(N__39420));
    Span4Mux_h I__7237 (
            .O(N__39423),
            .I(N__39417));
    LocalMux I__7236 (
            .O(N__39420),
            .I(N__39414));
    Span4Mux_v I__7235 (
            .O(N__39417),
            .I(N__39411));
    Span4Mux_v I__7234 (
            .O(N__39414),
            .I(N__39408));
    Odrv4 I__7233 (
            .O(N__39411),
            .I(\c0.n20171 ));
    Odrv4 I__7232 (
            .O(N__39408),
            .I(\c0.n20171 ));
    InMux I__7231 (
            .O(N__39403),
            .I(N__39400));
    LocalMux I__7230 (
            .O(N__39400),
            .I(\c0.data_out_frame_29__7__N_847 ));
    CascadeMux I__7229 (
            .O(N__39397),
            .I(\c0.data_out_frame_29__7__N_847_cascade_ ));
    CascadeMux I__7228 (
            .O(N__39394),
            .I(N__39387));
    CascadeMux I__7227 (
            .O(N__39393),
            .I(N__39384));
    CascadeMux I__7226 (
            .O(N__39392),
            .I(N__39381));
    CascadeMux I__7225 (
            .O(N__39391),
            .I(N__39378));
    CascadeMux I__7224 (
            .O(N__39390),
            .I(N__39375));
    InMux I__7223 (
            .O(N__39387),
            .I(N__39372));
    InMux I__7222 (
            .O(N__39384),
            .I(N__39367));
    InMux I__7221 (
            .O(N__39381),
            .I(N__39367));
    InMux I__7220 (
            .O(N__39378),
            .I(N__39364));
    InMux I__7219 (
            .O(N__39375),
            .I(N__39361));
    LocalMux I__7218 (
            .O(N__39372),
            .I(N__39355));
    LocalMux I__7217 (
            .O(N__39367),
            .I(N__39355));
    LocalMux I__7216 (
            .O(N__39364),
            .I(N__39350));
    LocalMux I__7215 (
            .O(N__39361),
            .I(N__39350));
    InMux I__7214 (
            .O(N__39360),
            .I(N__39347));
    Odrv4 I__7213 (
            .O(N__39355),
            .I(encoder0_position_11));
    Odrv12 I__7212 (
            .O(N__39350),
            .I(encoder0_position_11));
    LocalMux I__7211 (
            .O(N__39347),
            .I(encoder0_position_11));
    InMux I__7210 (
            .O(N__39340),
            .I(N__39337));
    LocalMux I__7209 (
            .O(N__39337),
            .I(\c0.n10_adj_4332 ));
    CascadeMux I__7208 (
            .O(N__39334),
            .I(N__39331));
    InMux I__7207 (
            .O(N__39331),
            .I(N__39328));
    LocalMux I__7206 (
            .O(N__39328),
            .I(N__39325));
    Span4Mux_h I__7205 (
            .O(N__39325),
            .I(N__39321));
    InMux I__7204 (
            .O(N__39324),
            .I(N__39314));
    Span4Mux_h I__7203 (
            .O(N__39321),
            .I(N__39311));
    InMux I__7202 (
            .O(N__39320),
            .I(N__39308));
    InMux I__7201 (
            .O(N__39319),
            .I(N__39301));
    InMux I__7200 (
            .O(N__39318),
            .I(N__39301));
    InMux I__7199 (
            .O(N__39317),
            .I(N__39301));
    LocalMux I__7198 (
            .O(N__39314),
            .I(encoder0_position_24));
    Odrv4 I__7197 (
            .O(N__39311),
            .I(encoder0_position_24));
    LocalMux I__7196 (
            .O(N__39308),
            .I(encoder0_position_24));
    LocalMux I__7195 (
            .O(N__39301),
            .I(encoder0_position_24));
    InMux I__7194 (
            .O(N__39292),
            .I(N__39289));
    LocalMux I__7193 (
            .O(N__39289),
            .I(N__39285));
    InMux I__7192 (
            .O(N__39288),
            .I(N__39282));
    Span12Mux_v I__7191 (
            .O(N__39285),
            .I(N__39279));
    LocalMux I__7190 (
            .O(N__39282),
            .I(\c0.n21931 ));
    Odrv12 I__7189 (
            .O(N__39279),
            .I(\c0.n21931 ));
    InMux I__7188 (
            .O(N__39274),
            .I(N__39270));
    InMux I__7187 (
            .O(N__39273),
            .I(N__39265));
    LocalMux I__7186 (
            .O(N__39270),
            .I(N__39261));
    InMux I__7185 (
            .O(N__39269),
            .I(N__39258));
    InMux I__7184 (
            .O(N__39268),
            .I(N__39255));
    LocalMux I__7183 (
            .O(N__39265),
            .I(N__39252));
    InMux I__7182 (
            .O(N__39264),
            .I(N__39249));
    Span4Mux_h I__7181 (
            .O(N__39261),
            .I(N__39243));
    LocalMux I__7180 (
            .O(N__39258),
            .I(N__39243));
    LocalMux I__7179 (
            .O(N__39255),
            .I(N__39236));
    Span4Mux_v I__7178 (
            .O(N__39252),
            .I(N__39236));
    LocalMux I__7177 (
            .O(N__39249),
            .I(N__39236));
    InMux I__7176 (
            .O(N__39248),
            .I(N__39233));
    Span4Mux_v I__7175 (
            .O(N__39243),
            .I(N__39230));
    Span4Mux_h I__7174 (
            .O(N__39236),
            .I(N__39225));
    LocalMux I__7173 (
            .O(N__39233),
            .I(N__39225));
    Odrv4 I__7172 (
            .O(N__39230),
            .I(\c0.r_SM_Main_2_N_3755_0 ));
    Odrv4 I__7171 (
            .O(N__39225),
            .I(\c0.r_SM_Main_2_N_3755_0 ));
    CEMux I__7170 (
            .O(N__39220),
            .I(N__39217));
    LocalMux I__7169 (
            .O(N__39217),
            .I(N__39214));
    Span4Mux_h I__7168 (
            .O(N__39214),
            .I(N__39211));
    Span4Mux_h I__7167 (
            .O(N__39211),
            .I(N__39208));
    Odrv4 I__7166 (
            .O(N__39208),
            .I(\c0.n14322 ));
    CascadeMux I__7165 (
            .O(N__39205),
            .I(\c0.n14322_cascade_ ));
    SRMux I__7164 (
            .O(N__39202),
            .I(N__39199));
    LocalMux I__7163 (
            .O(N__39199),
            .I(N__39196));
    Span12Mux_s8_h I__7162 (
            .O(N__39196),
            .I(N__39193));
    Odrv12 I__7161 (
            .O(N__39193),
            .I(\c0.n14871 ));
    CascadeMux I__7160 (
            .O(N__39190),
            .I(N__39186));
    InMux I__7159 (
            .O(N__39189),
            .I(N__39183));
    InMux I__7158 (
            .O(N__39186),
            .I(N__39180));
    LocalMux I__7157 (
            .O(N__39183),
            .I(N__39177));
    LocalMux I__7156 (
            .O(N__39180),
            .I(N__39174));
    Span4Mux_h I__7155 (
            .O(N__39177),
            .I(N__39171));
    Odrv12 I__7154 (
            .O(N__39174),
            .I(\c0.tx_transmit_N_3651 ));
    Odrv4 I__7153 (
            .O(N__39171),
            .I(\c0.tx_transmit_N_3651 ));
    InMux I__7152 (
            .O(N__39166),
            .I(N__39163));
    LocalMux I__7151 (
            .O(N__39163),
            .I(\c0.n23975 ));
    InMux I__7150 (
            .O(N__39160),
            .I(N__39157));
    LocalMux I__7149 (
            .O(N__39157),
            .I(N__39154));
    Span4Mux_v I__7148 (
            .O(N__39154),
            .I(N__39151));
    Odrv4 I__7147 (
            .O(N__39151),
            .I(\c0.n18_adj_4403 ));
    InMux I__7146 (
            .O(N__39148),
            .I(N__39145));
    LocalMux I__7145 (
            .O(N__39145),
            .I(N__39142));
    Odrv12 I__7144 (
            .O(N__39142),
            .I(\c0.n20875 ));
    InMux I__7143 (
            .O(N__39139),
            .I(N__39135));
    InMux I__7142 (
            .O(N__39138),
            .I(N__39132));
    LocalMux I__7141 (
            .O(N__39135),
            .I(\c0.n17602 ));
    LocalMux I__7140 (
            .O(N__39132),
            .I(\c0.n17602 ));
    InMux I__7139 (
            .O(N__39127),
            .I(N__39124));
    LocalMux I__7138 (
            .O(N__39124),
            .I(N__39121));
    Span4Mux_v I__7137 (
            .O(N__39121),
            .I(N__39118));
    Odrv4 I__7136 (
            .O(N__39118),
            .I(n2255));
    InMux I__7135 (
            .O(N__39115),
            .I(N__39111));
    CascadeMux I__7134 (
            .O(N__39114),
            .I(N__39108));
    LocalMux I__7133 (
            .O(N__39111),
            .I(N__39105));
    InMux I__7132 (
            .O(N__39108),
            .I(N__39102));
    Span4Mux_v I__7131 (
            .O(N__39105),
            .I(N__39098));
    LocalMux I__7130 (
            .O(N__39102),
            .I(N__39095));
    InMux I__7129 (
            .O(N__39101),
            .I(N__39092));
    Span4Mux_h I__7128 (
            .O(N__39098),
            .I(N__39086));
    Span4Mux_h I__7127 (
            .O(N__39095),
            .I(N__39081));
    LocalMux I__7126 (
            .O(N__39092),
            .I(N__39081));
    InMux I__7125 (
            .O(N__39091),
            .I(N__39078));
    InMux I__7124 (
            .O(N__39090),
            .I(N__39073));
    InMux I__7123 (
            .O(N__39089),
            .I(N__39073));
    Odrv4 I__7122 (
            .O(N__39086),
            .I(encoder0_position_16));
    Odrv4 I__7121 (
            .O(N__39081),
            .I(encoder0_position_16));
    LocalMux I__7120 (
            .O(N__39078),
            .I(encoder0_position_16));
    LocalMux I__7119 (
            .O(N__39073),
            .I(encoder0_position_16));
    InMux I__7118 (
            .O(N__39064),
            .I(N__39061));
    LocalMux I__7117 (
            .O(N__39061),
            .I(N__39057));
    InMux I__7116 (
            .O(N__39060),
            .I(N__39053));
    Span4Mux_h I__7115 (
            .O(N__39057),
            .I(N__39050));
    InMux I__7114 (
            .O(N__39056),
            .I(N__39047));
    LocalMux I__7113 (
            .O(N__39053),
            .I(\c0.n22408 ));
    Odrv4 I__7112 (
            .O(N__39050),
            .I(\c0.n22408 ));
    LocalMux I__7111 (
            .O(N__39047),
            .I(\c0.n22408 ));
    InMux I__7110 (
            .O(N__39040),
            .I(N__39037));
    LocalMux I__7109 (
            .O(N__39037),
            .I(N__39032));
    InMux I__7108 (
            .O(N__39036),
            .I(N__39029));
    InMux I__7107 (
            .O(N__39035),
            .I(N__39026));
    Span4Mux_h I__7106 (
            .O(N__39032),
            .I(N__39023));
    LocalMux I__7105 (
            .O(N__39029),
            .I(N__39020));
    LocalMux I__7104 (
            .O(N__39026),
            .I(N__39017));
    Span4Mux_v I__7103 (
            .O(N__39023),
            .I(N__39009));
    Span4Mux_v I__7102 (
            .O(N__39020),
            .I(N__39009));
    Span4Mux_h I__7101 (
            .O(N__39017),
            .I(N__39006));
    InMux I__7100 (
            .O(N__39016),
            .I(N__39001));
    InMux I__7099 (
            .O(N__39015),
            .I(N__39001));
    InMux I__7098 (
            .O(N__39014),
            .I(N__38998));
    Odrv4 I__7097 (
            .O(N__39009),
            .I(encoder0_position_4));
    Odrv4 I__7096 (
            .O(N__39006),
            .I(encoder0_position_4));
    LocalMux I__7095 (
            .O(N__39001),
            .I(encoder0_position_4));
    LocalMux I__7094 (
            .O(N__38998),
            .I(encoder0_position_4));
    CascadeMux I__7093 (
            .O(N__38989),
            .I(\c0.n22227_cascade_ ));
    InMux I__7092 (
            .O(N__38986),
            .I(N__38982));
    InMux I__7091 (
            .O(N__38985),
            .I(N__38979));
    LocalMux I__7090 (
            .O(N__38982),
            .I(N__38976));
    LocalMux I__7089 (
            .O(N__38979),
            .I(\c0.n22128 ));
    Odrv4 I__7088 (
            .O(N__38976),
            .I(\c0.n22128 ));
    CascadeMux I__7087 (
            .O(N__38971),
            .I(N__38968));
    InMux I__7086 (
            .O(N__38968),
            .I(N__38958));
    InMux I__7085 (
            .O(N__38967),
            .I(N__38958));
    InMux I__7084 (
            .O(N__38966),
            .I(N__38958));
    InMux I__7083 (
            .O(N__38965),
            .I(N__38955));
    LocalMux I__7082 (
            .O(N__38958),
            .I(N__38950));
    LocalMux I__7081 (
            .O(N__38955),
            .I(N__38950));
    Span4Mux_h I__7080 (
            .O(N__38950),
            .I(N__38947));
    Span4Mux_v I__7079 (
            .O(N__38947),
            .I(N__38944));
    Odrv4 I__7078 (
            .O(N__38944),
            .I(\c0.n10444 ));
    CascadeMux I__7077 (
            .O(N__38941),
            .I(N__38938));
    InMux I__7076 (
            .O(N__38938),
            .I(N__38935));
    LocalMux I__7075 (
            .O(N__38935),
            .I(N__38931));
    CascadeMux I__7074 (
            .O(N__38934),
            .I(N__38928));
    Span4Mux_h I__7073 (
            .O(N__38931),
            .I(N__38925));
    InMux I__7072 (
            .O(N__38928),
            .I(N__38922));
    Span4Mux_v I__7071 (
            .O(N__38925),
            .I(N__38917));
    LocalMux I__7070 (
            .O(N__38922),
            .I(N__38917));
    Span4Mux_h I__7069 (
            .O(N__38917),
            .I(N__38911));
    InMux I__7068 (
            .O(N__38916),
            .I(N__38906));
    InMux I__7067 (
            .O(N__38915),
            .I(N__38906));
    InMux I__7066 (
            .O(N__38914),
            .I(N__38902));
    Span4Mux_h I__7065 (
            .O(N__38911),
            .I(N__38897));
    LocalMux I__7064 (
            .O(N__38906),
            .I(N__38897));
    InMux I__7063 (
            .O(N__38905),
            .I(N__38894));
    LocalMux I__7062 (
            .O(N__38902),
            .I(encoder1_position_20));
    Odrv4 I__7061 (
            .O(N__38897),
            .I(encoder1_position_20));
    LocalMux I__7060 (
            .O(N__38894),
            .I(encoder1_position_20));
    CascadeMux I__7059 (
            .O(N__38887),
            .I(N__38884));
    InMux I__7058 (
            .O(N__38884),
            .I(N__38881));
    LocalMux I__7057 (
            .O(N__38881),
            .I(N__38878));
    Odrv12 I__7056 (
            .O(N__38878),
            .I(\c0.n6_adj_4312 ));
    InMux I__7055 (
            .O(N__38875),
            .I(N__38871));
    InMux I__7054 (
            .O(N__38874),
            .I(N__38866));
    LocalMux I__7053 (
            .O(N__38871),
            .I(N__38863));
    InMux I__7052 (
            .O(N__38870),
            .I(N__38860));
    InMux I__7051 (
            .O(N__38869),
            .I(N__38856));
    LocalMux I__7050 (
            .O(N__38866),
            .I(N__38851));
    Span4Mux_h I__7049 (
            .O(N__38863),
            .I(N__38851));
    LocalMux I__7048 (
            .O(N__38860),
            .I(N__38848));
    InMux I__7047 (
            .O(N__38859),
            .I(N__38844));
    LocalMux I__7046 (
            .O(N__38856),
            .I(N__38841));
    Span4Mux_h I__7045 (
            .O(N__38851),
            .I(N__38838));
    Span12Mux_h I__7044 (
            .O(N__38848),
            .I(N__38835));
    InMux I__7043 (
            .O(N__38847),
            .I(N__38832));
    LocalMux I__7042 (
            .O(N__38844),
            .I(encoder0_position_12));
    Odrv4 I__7041 (
            .O(N__38841),
            .I(encoder0_position_12));
    Odrv4 I__7040 (
            .O(N__38838),
            .I(encoder0_position_12));
    Odrv12 I__7039 (
            .O(N__38835),
            .I(encoder0_position_12));
    LocalMux I__7038 (
            .O(N__38832),
            .I(encoder0_position_12));
    InMux I__7037 (
            .O(N__38821),
            .I(N__38818));
    LocalMux I__7036 (
            .O(N__38818),
            .I(N__38815));
    Odrv4 I__7035 (
            .O(N__38815),
            .I(\c0.n22477 ));
    CascadeMux I__7034 (
            .O(N__38812),
            .I(\c0.n22477_cascade_ ));
    InMux I__7033 (
            .O(N__38809),
            .I(N__38806));
    LocalMux I__7032 (
            .O(N__38806),
            .I(N__38803));
    Odrv4 I__7031 (
            .O(N__38803),
            .I(\c0.n6_adj_4333 ));
    InMux I__7030 (
            .O(N__38800),
            .I(N__38797));
    LocalMux I__7029 (
            .O(N__38797),
            .I(N__38794));
    Span4Mux_h I__7028 (
            .O(N__38794),
            .I(N__38791));
    Span4Mux_h I__7027 (
            .O(N__38791),
            .I(N__38788));
    Odrv4 I__7026 (
            .O(N__38788),
            .I(n2243));
    CascadeMux I__7025 (
            .O(N__38785),
            .I(N__38780));
    InMux I__7024 (
            .O(N__38784),
            .I(N__38777));
    InMux I__7023 (
            .O(N__38783),
            .I(N__38774));
    InMux I__7022 (
            .O(N__38780),
            .I(N__38768));
    LocalMux I__7021 (
            .O(N__38777),
            .I(N__38765));
    LocalMux I__7020 (
            .O(N__38774),
            .I(N__38762));
    InMux I__7019 (
            .O(N__38773),
            .I(N__38757));
    InMux I__7018 (
            .O(N__38772),
            .I(N__38757));
    InMux I__7017 (
            .O(N__38771),
            .I(N__38753));
    LocalMux I__7016 (
            .O(N__38768),
            .I(N__38750));
    Span4Mux_h I__7015 (
            .O(N__38765),
            .I(N__38745));
    Span4Mux_h I__7014 (
            .O(N__38762),
            .I(N__38745));
    LocalMux I__7013 (
            .O(N__38757),
            .I(N__38742));
    InMux I__7012 (
            .O(N__38756),
            .I(N__38739));
    LocalMux I__7011 (
            .O(N__38753),
            .I(encoder0_position_28));
    Odrv4 I__7010 (
            .O(N__38750),
            .I(encoder0_position_28));
    Odrv4 I__7009 (
            .O(N__38745),
            .I(encoder0_position_28));
    Odrv4 I__7008 (
            .O(N__38742),
            .I(encoder0_position_28));
    LocalMux I__7007 (
            .O(N__38739),
            .I(encoder0_position_28));
    CascadeMux I__7006 (
            .O(N__38728),
            .I(N__38725));
    InMux I__7005 (
            .O(N__38725),
            .I(N__38719));
    InMux I__7004 (
            .O(N__38724),
            .I(N__38716));
    CascadeMux I__7003 (
            .O(N__38723),
            .I(N__38711));
    InMux I__7002 (
            .O(N__38722),
            .I(N__38708));
    LocalMux I__7001 (
            .O(N__38719),
            .I(N__38705));
    LocalMux I__7000 (
            .O(N__38716),
            .I(N__38702));
    InMux I__6999 (
            .O(N__38715),
            .I(N__38697));
    InMux I__6998 (
            .O(N__38714),
            .I(N__38697));
    InMux I__6997 (
            .O(N__38711),
            .I(N__38694));
    LocalMux I__6996 (
            .O(N__38708),
            .I(N__38687));
    Span4Mux_h I__6995 (
            .O(N__38705),
            .I(N__38687));
    Span4Mux_h I__6994 (
            .O(N__38702),
            .I(N__38687));
    LocalMux I__6993 (
            .O(N__38697),
            .I(N__38684));
    LocalMux I__6992 (
            .O(N__38694),
            .I(encoder0_position_9));
    Odrv4 I__6991 (
            .O(N__38687),
            .I(encoder0_position_9));
    Odrv4 I__6990 (
            .O(N__38684),
            .I(encoder0_position_9));
    InMux I__6989 (
            .O(N__38677),
            .I(N__38671));
    InMux I__6988 (
            .O(N__38676),
            .I(N__38671));
    LocalMux I__6987 (
            .O(N__38671),
            .I(\c0.n22427 ));
    CascadeMux I__6986 (
            .O(N__38668),
            .I(N__38663));
    InMux I__6985 (
            .O(N__38667),
            .I(N__38659));
    InMux I__6984 (
            .O(N__38666),
            .I(N__38656));
    InMux I__6983 (
            .O(N__38663),
            .I(N__38653));
    CascadeMux I__6982 (
            .O(N__38662),
            .I(N__38649));
    LocalMux I__6981 (
            .O(N__38659),
            .I(N__38645));
    LocalMux I__6980 (
            .O(N__38656),
            .I(N__38642));
    LocalMux I__6979 (
            .O(N__38653),
            .I(N__38639));
    InMux I__6978 (
            .O(N__38652),
            .I(N__38636));
    InMux I__6977 (
            .O(N__38649),
            .I(N__38633));
    InMux I__6976 (
            .O(N__38648),
            .I(N__38630));
    Span4Mux_h I__6975 (
            .O(N__38645),
            .I(N__38627));
    Span4Mux_h I__6974 (
            .O(N__38642),
            .I(N__38622));
    Span4Mux_h I__6973 (
            .O(N__38639),
            .I(N__38622));
    LocalMux I__6972 (
            .O(N__38636),
            .I(encoder0_position_19));
    LocalMux I__6971 (
            .O(N__38633),
            .I(encoder0_position_19));
    LocalMux I__6970 (
            .O(N__38630),
            .I(encoder0_position_19));
    Odrv4 I__6969 (
            .O(N__38627),
            .I(encoder0_position_19));
    Odrv4 I__6968 (
            .O(N__38622),
            .I(encoder0_position_19));
    CascadeMux I__6967 (
            .O(N__38611),
            .I(N__38607));
    InMux I__6966 (
            .O(N__38610),
            .I(N__38602));
    InMux I__6965 (
            .O(N__38607),
            .I(N__38602));
    LocalMux I__6964 (
            .O(N__38602),
            .I(\c0.n21885 ));
    InMux I__6963 (
            .O(N__38599),
            .I(N__38596));
    LocalMux I__6962 (
            .O(N__38596),
            .I(\c0.n22200 ));
    CascadeMux I__6961 (
            .O(N__38593),
            .I(\c0.n22200_cascade_ ));
    InMux I__6960 (
            .O(N__38590),
            .I(N__38587));
    LocalMux I__6959 (
            .O(N__38587),
            .I(N__38583));
    InMux I__6958 (
            .O(N__38586),
            .I(N__38580));
    Span4Mux_h I__6957 (
            .O(N__38583),
            .I(N__38576));
    LocalMux I__6956 (
            .O(N__38580),
            .I(N__38573));
    InMux I__6955 (
            .O(N__38579),
            .I(N__38570));
    Odrv4 I__6954 (
            .O(N__38576),
            .I(\c0.n21970 ));
    Odrv12 I__6953 (
            .O(N__38573),
            .I(\c0.n21970 ));
    LocalMux I__6952 (
            .O(N__38570),
            .I(\c0.n21970 ));
    InMux I__6951 (
            .O(N__38563),
            .I(N__38560));
    LocalMux I__6950 (
            .O(N__38560),
            .I(N__38557));
    Span4Mux_h I__6949 (
            .O(N__38557),
            .I(N__38553));
    InMux I__6948 (
            .O(N__38556),
            .I(N__38550));
    Odrv4 I__6947 (
            .O(N__38553),
            .I(\c0.n13705 ));
    LocalMux I__6946 (
            .O(N__38550),
            .I(\c0.n13705 ));
    InMux I__6945 (
            .O(N__38545),
            .I(N__38542));
    LocalMux I__6944 (
            .O(N__38542),
            .I(N__38539));
    Odrv12 I__6943 (
            .O(N__38539),
            .I(n2259));
    InMux I__6942 (
            .O(N__38536),
            .I(N__38533));
    LocalMux I__6941 (
            .O(N__38533),
            .I(N__38530));
    Span4Mux_v I__6940 (
            .O(N__38530),
            .I(N__38527));
    Odrv4 I__6939 (
            .O(N__38527),
            .I(n2267));
    InMux I__6938 (
            .O(N__38524),
            .I(N__38521));
    LocalMux I__6937 (
            .O(N__38521),
            .I(N__38518));
    Odrv4 I__6936 (
            .O(N__38518),
            .I(n2261));
    InMux I__6935 (
            .O(N__38515),
            .I(N__38512));
    LocalMux I__6934 (
            .O(N__38512),
            .I(N__38509));
    Odrv12 I__6933 (
            .O(N__38509),
            .I(\c0.n21908 ));
    InMux I__6932 (
            .O(N__38506),
            .I(N__38493));
    InMux I__6931 (
            .O(N__38505),
            .I(N__38488));
    InMux I__6930 (
            .O(N__38504),
            .I(N__38485));
    InMux I__6929 (
            .O(N__38503),
            .I(N__38482));
    InMux I__6928 (
            .O(N__38502),
            .I(N__38473));
    InMux I__6927 (
            .O(N__38501),
            .I(N__38473));
    InMux I__6926 (
            .O(N__38500),
            .I(N__38473));
    InMux I__6925 (
            .O(N__38499),
            .I(N__38473));
    InMux I__6924 (
            .O(N__38498),
            .I(N__38470));
    InMux I__6923 (
            .O(N__38497),
            .I(N__38467));
    CascadeMux I__6922 (
            .O(N__38496),
            .I(N__38462));
    LocalMux I__6921 (
            .O(N__38493),
            .I(N__38454));
    InMux I__6920 (
            .O(N__38492),
            .I(N__38449));
    InMux I__6919 (
            .O(N__38491),
            .I(N__38449));
    LocalMux I__6918 (
            .O(N__38488),
            .I(N__38446));
    LocalMux I__6917 (
            .O(N__38485),
            .I(N__38443));
    LocalMux I__6916 (
            .O(N__38482),
            .I(N__38434));
    LocalMux I__6915 (
            .O(N__38473),
            .I(N__38434));
    LocalMux I__6914 (
            .O(N__38470),
            .I(N__38434));
    LocalMux I__6913 (
            .O(N__38467),
            .I(N__38434));
    InMux I__6912 (
            .O(N__38466),
            .I(N__38431));
    InMux I__6911 (
            .O(N__38465),
            .I(N__38424));
    InMux I__6910 (
            .O(N__38462),
            .I(N__38424));
    InMux I__6909 (
            .O(N__38461),
            .I(N__38424));
    InMux I__6908 (
            .O(N__38460),
            .I(N__38419));
    InMux I__6907 (
            .O(N__38459),
            .I(N__38419));
    InMux I__6906 (
            .O(N__38458),
            .I(N__38416));
    InMux I__6905 (
            .O(N__38457),
            .I(N__38413));
    Span4Mux_h I__6904 (
            .O(N__38454),
            .I(N__38405));
    LocalMux I__6903 (
            .O(N__38449),
            .I(N__38405));
    Span4Mux_v I__6902 (
            .O(N__38446),
            .I(N__38402));
    Span4Mux_v I__6901 (
            .O(N__38443),
            .I(N__38397));
    Span4Mux_v I__6900 (
            .O(N__38434),
            .I(N__38397));
    LocalMux I__6899 (
            .O(N__38431),
            .I(N__38388));
    LocalMux I__6898 (
            .O(N__38424),
            .I(N__38388));
    LocalMux I__6897 (
            .O(N__38419),
            .I(N__38388));
    LocalMux I__6896 (
            .O(N__38416),
            .I(N__38383));
    LocalMux I__6895 (
            .O(N__38413),
            .I(N__38383));
    InMux I__6894 (
            .O(N__38412),
            .I(N__38378));
    InMux I__6893 (
            .O(N__38411),
            .I(N__38378));
    CascadeMux I__6892 (
            .O(N__38410),
            .I(N__38374));
    Span4Mux_v I__6891 (
            .O(N__38405),
            .I(N__38367));
    Span4Mux_h I__6890 (
            .O(N__38402),
            .I(N__38367));
    Span4Mux_h I__6889 (
            .O(N__38397),
            .I(N__38367));
    InMux I__6888 (
            .O(N__38396),
            .I(N__38364));
    InMux I__6887 (
            .O(N__38395),
            .I(N__38361));
    Span12Mux_v I__6886 (
            .O(N__38388),
            .I(N__38353));
    Span4Mux_v I__6885 (
            .O(N__38383),
            .I(N__38348));
    LocalMux I__6884 (
            .O(N__38378),
            .I(N__38348));
    InMux I__6883 (
            .O(N__38377),
            .I(N__38343));
    InMux I__6882 (
            .O(N__38374),
            .I(N__38343));
    Sp12to4 I__6881 (
            .O(N__38367),
            .I(N__38336));
    LocalMux I__6880 (
            .O(N__38364),
            .I(N__38336));
    LocalMux I__6879 (
            .O(N__38361),
            .I(N__38336));
    InMux I__6878 (
            .O(N__38360),
            .I(N__38327));
    InMux I__6877 (
            .O(N__38359),
            .I(N__38327));
    InMux I__6876 (
            .O(N__38358),
            .I(N__38327));
    InMux I__6875 (
            .O(N__38357),
            .I(N__38327));
    InMux I__6874 (
            .O(N__38356),
            .I(N__38324));
    Odrv12 I__6873 (
            .O(N__38353),
            .I(count_enable_adj_4544));
    Odrv4 I__6872 (
            .O(N__38348),
            .I(count_enable_adj_4544));
    LocalMux I__6871 (
            .O(N__38343),
            .I(count_enable_adj_4544));
    Odrv12 I__6870 (
            .O(N__38336),
            .I(count_enable_adj_4544));
    LocalMux I__6869 (
            .O(N__38327),
            .I(count_enable_adj_4544));
    LocalMux I__6868 (
            .O(N__38324),
            .I(count_enable_adj_4544));
    InMux I__6867 (
            .O(N__38311),
            .I(N__38308));
    LocalMux I__6866 (
            .O(N__38308),
            .I(N__38305));
    Span4Mux_h I__6865 (
            .O(N__38305),
            .I(N__38302));
    Span4Mux_h I__6864 (
            .O(N__38302),
            .I(N__38299));
    Odrv4 I__6863 (
            .O(N__38299),
            .I(n2185));
    InMux I__6862 (
            .O(N__38296),
            .I(N__38291));
    InMux I__6861 (
            .O(N__38295),
            .I(N__38288));
    InMux I__6860 (
            .O(N__38294),
            .I(N__38285));
    LocalMux I__6859 (
            .O(N__38291),
            .I(N__38282));
    LocalMux I__6858 (
            .O(N__38288),
            .I(N__38279));
    LocalMux I__6857 (
            .O(N__38285),
            .I(N__38276));
    Span4Mux_v I__6856 (
            .O(N__38282),
            .I(N__38273));
    Span4Mux_v I__6855 (
            .O(N__38279),
            .I(N__38270));
    Span4Mux_h I__6854 (
            .O(N__38276),
            .I(N__38267));
    Sp12to4 I__6853 (
            .O(N__38273),
            .I(N__38264));
    Odrv4 I__6852 (
            .O(N__38270),
            .I(\c0.n13839 ));
    Odrv4 I__6851 (
            .O(N__38267),
            .I(\c0.n13839 ));
    Odrv12 I__6850 (
            .O(N__38264),
            .I(\c0.n13839 ));
    InMux I__6849 (
            .O(N__38257),
            .I(N__38254));
    LocalMux I__6848 (
            .O(N__38254),
            .I(N__38251));
    Odrv4 I__6847 (
            .O(N__38251),
            .I(\c0.n22015 ));
    CascadeMux I__6846 (
            .O(N__38248),
            .I(N__38239));
    InMux I__6845 (
            .O(N__38247),
            .I(N__38236));
    InMux I__6844 (
            .O(N__38246),
            .I(N__38233));
    CascadeMux I__6843 (
            .O(N__38245),
            .I(N__38230));
    InMux I__6842 (
            .O(N__38244),
            .I(N__38227));
    InMux I__6841 (
            .O(N__38243),
            .I(N__38222));
    InMux I__6840 (
            .O(N__38242),
            .I(N__38222));
    InMux I__6839 (
            .O(N__38239),
            .I(N__38218));
    LocalMux I__6838 (
            .O(N__38236),
            .I(N__38215));
    LocalMux I__6837 (
            .O(N__38233),
            .I(N__38212));
    InMux I__6836 (
            .O(N__38230),
            .I(N__38209));
    LocalMux I__6835 (
            .O(N__38227),
            .I(N__38204));
    LocalMux I__6834 (
            .O(N__38222),
            .I(N__38204));
    InMux I__6833 (
            .O(N__38221),
            .I(N__38201));
    LocalMux I__6832 (
            .O(N__38218),
            .I(N__38196));
    Span4Mux_v I__6831 (
            .O(N__38215),
            .I(N__38196));
    Span4Mux_h I__6830 (
            .O(N__38212),
            .I(N__38193));
    LocalMux I__6829 (
            .O(N__38209),
            .I(N__38188));
    Span4Mux_h I__6828 (
            .O(N__38204),
            .I(N__38188));
    LocalMux I__6827 (
            .O(N__38201),
            .I(encoder0_position_29));
    Odrv4 I__6826 (
            .O(N__38196),
            .I(encoder0_position_29));
    Odrv4 I__6825 (
            .O(N__38193),
            .I(encoder0_position_29));
    Odrv4 I__6824 (
            .O(N__38188),
            .I(encoder0_position_29));
    InMux I__6823 (
            .O(N__38179),
            .I(N__38176));
    LocalMux I__6822 (
            .O(N__38176),
            .I(N__38173));
    Span4Mux_h I__6821 (
            .O(N__38173),
            .I(N__38170));
    Odrv4 I__6820 (
            .O(N__38170),
            .I(\c0.data_out_frame_29__7__N_856 ));
    InMux I__6819 (
            .O(N__38167),
            .I(N__38164));
    LocalMux I__6818 (
            .O(N__38164),
            .I(N__38160));
    InMux I__6817 (
            .O(N__38163),
            .I(N__38157));
    Span4Mux_h I__6816 (
            .O(N__38160),
            .I(N__38154));
    LocalMux I__6815 (
            .O(N__38157),
            .I(\c0.n22382 ));
    Odrv4 I__6814 (
            .O(N__38154),
            .I(\c0.n22382 ));
    CascadeMux I__6813 (
            .O(N__38149),
            .I(N__38146));
    InMux I__6812 (
            .O(N__38146),
            .I(N__38143));
    LocalMux I__6811 (
            .O(N__38143),
            .I(N__38140));
    Odrv4 I__6810 (
            .O(N__38140),
            .I(\c0.n6_adj_4311 ));
    InMux I__6809 (
            .O(N__38137),
            .I(N__38134));
    LocalMux I__6808 (
            .O(N__38134),
            .I(\c0.n14_adj_4400 ));
    CascadeMux I__6807 (
            .O(N__38131),
            .I(\c0.n17600_cascade_ ));
    InMux I__6806 (
            .O(N__38128),
            .I(N__38122));
    InMux I__6805 (
            .O(N__38127),
            .I(N__38122));
    LocalMux I__6804 (
            .O(N__38122),
            .I(\c0.data_in_frame_10_4 ));
    SRMux I__6803 (
            .O(N__38119),
            .I(N__38116));
    LocalMux I__6802 (
            .O(N__38116),
            .I(N__38113));
    Odrv12 I__6801 (
            .O(N__38113),
            .I(\c0.n21342 ));
    InMux I__6800 (
            .O(N__38110),
            .I(N__38104));
    InMux I__6799 (
            .O(N__38109),
            .I(N__38101));
    InMux I__6798 (
            .O(N__38108),
            .I(N__38098));
    InMux I__6797 (
            .O(N__38107),
            .I(N__38095));
    LocalMux I__6796 (
            .O(N__38104),
            .I(N__38088));
    LocalMux I__6795 (
            .O(N__38101),
            .I(N__38088));
    LocalMux I__6794 (
            .O(N__38098),
            .I(N__38088));
    LocalMux I__6793 (
            .O(N__38095),
            .I(\c0.FRAME_MATCHER_state_11 ));
    Odrv12 I__6792 (
            .O(N__38088),
            .I(\c0.FRAME_MATCHER_state_11 ));
    SRMux I__6791 (
            .O(N__38083),
            .I(N__38080));
    LocalMux I__6790 (
            .O(N__38080),
            .I(N__38077));
    Span4Mux_h I__6789 (
            .O(N__38077),
            .I(N__38074));
    Odrv4 I__6788 (
            .O(N__38074),
            .I(\c0.n21350 ));
    CascadeMux I__6787 (
            .O(N__38071),
            .I(N__38067));
    CascadeMux I__6786 (
            .O(N__38070),
            .I(N__38064));
    InMux I__6785 (
            .O(N__38067),
            .I(N__38060));
    InMux I__6784 (
            .O(N__38064),
            .I(N__38056));
    InMux I__6783 (
            .O(N__38063),
            .I(N__38053));
    LocalMux I__6782 (
            .O(N__38060),
            .I(N__38050));
    InMux I__6781 (
            .O(N__38059),
            .I(N__38047));
    LocalMux I__6780 (
            .O(N__38056),
            .I(N__38043));
    LocalMux I__6779 (
            .O(N__38053),
            .I(N__38040));
    Span4Mux_v I__6778 (
            .O(N__38050),
            .I(N__38035));
    LocalMux I__6777 (
            .O(N__38047),
            .I(N__38035));
    InMux I__6776 (
            .O(N__38046),
            .I(N__38032));
    Span4Mux_h I__6775 (
            .O(N__38043),
            .I(N__38025));
    Span4Mux_v I__6774 (
            .O(N__38040),
            .I(N__38025));
    Span4Mux_v I__6773 (
            .O(N__38035),
            .I(N__38025));
    LocalMux I__6772 (
            .O(N__38032),
            .I(encoder1_position_13));
    Odrv4 I__6771 (
            .O(N__38025),
            .I(encoder1_position_13));
    InMux I__6770 (
            .O(N__38020),
            .I(N__38017));
    LocalMux I__6769 (
            .O(N__38017),
            .I(N__38014));
    Span4Mux_v I__6768 (
            .O(N__38014),
            .I(N__38011));
    Span4Mux_h I__6767 (
            .O(N__38011),
            .I(N__38008));
    Span4Mux_h I__6766 (
            .O(N__38008),
            .I(N__38004));
    InMux I__6765 (
            .O(N__38007),
            .I(N__38001));
    Span4Mux_v I__6764 (
            .O(N__38004),
            .I(N__37998));
    LocalMux I__6763 (
            .O(N__38001),
            .I(data_out_frame_12_5));
    Odrv4 I__6762 (
            .O(N__37998),
            .I(data_out_frame_12_5));
    InMux I__6761 (
            .O(N__37993),
            .I(N__37990));
    LocalMux I__6760 (
            .O(N__37990),
            .I(N__37987));
    Odrv4 I__6759 (
            .O(N__37987),
            .I(\c0.n14_adj_4364 ));
    InMux I__6758 (
            .O(N__37984),
            .I(N__37981));
    LocalMux I__6757 (
            .O(N__37981),
            .I(\c0.n13 ));
    CascadeMux I__6756 (
            .O(N__37978),
            .I(\c0.n13_adj_4366_cascade_ ));
    InMux I__6755 (
            .O(N__37975),
            .I(N__37972));
    LocalMux I__6754 (
            .O(N__37972),
            .I(\c0.n14_adj_4365 ));
    InMux I__6753 (
            .O(N__37969),
            .I(N__37966));
    LocalMux I__6752 (
            .O(N__37966),
            .I(N__37963));
    Span4Mux_v I__6751 (
            .O(N__37963),
            .I(N__37960));
    Odrv4 I__6750 (
            .O(N__37960),
            .I(\c0.n20_adj_4482 ));
    CascadeMux I__6749 (
            .O(N__37957),
            .I(\c0.n21_adj_4480_cascade_ ));
    InMux I__6748 (
            .O(N__37954),
            .I(N__37951));
    LocalMux I__6747 (
            .O(N__37951),
            .I(N__37948));
    Odrv4 I__6746 (
            .O(N__37948),
            .I(\c0.n19_adj_4481 ));
    InMux I__6745 (
            .O(N__37945),
            .I(N__37941));
    CascadeMux I__6744 (
            .O(N__37944),
            .I(N__37937));
    LocalMux I__6743 (
            .O(N__37941),
            .I(N__37934));
    InMux I__6742 (
            .O(N__37940),
            .I(N__37931));
    InMux I__6741 (
            .O(N__37937),
            .I(N__37928));
    Span12Mux_h I__6740 (
            .O(N__37934),
            .I(N__37921));
    LocalMux I__6739 (
            .O(N__37931),
            .I(N__37921));
    LocalMux I__6738 (
            .O(N__37928),
            .I(N__37921));
    Odrv12 I__6737 (
            .O(N__37921),
            .I(\c0.n14789 ));
    CascadeMux I__6736 (
            .O(N__37918),
            .I(N__37915));
    InMux I__6735 (
            .O(N__37915),
            .I(N__37910));
    InMux I__6734 (
            .O(N__37914),
            .I(N__37907));
    InMux I__6733 (
            .O(N__37913),
            .I(N__37904));
    LocalMux I__6732 (
            .O(N__37910),
            .I(N__37896));
    LocalMux I__6731 (
            .O(N__37907),
            .I(N__37896));
    LocalMux I__6730 (
            .O(N__37904),
            .I(N__37896));
    InMux I__6729 (
            .O(N__37903),
            .I(N__37893));
    Span4Mux_v I__6728 (
            .O(N__37896),
            .I(N__37890));
    LocalMux I__6727 (
            .O(N__37893),
            .I(\c0.FRAME_MATCHER_state_18 ));
    Odrv4 I__6726 (
            .O(N__37890),
            .I(\c0.FRAME_MATCHER_state_18 ));
    CascadeMux I__6725 (
            .O(N__37885),
            .I(N__37882));
    InMux I__6724 (
            .O(N__37882),
            .I(N__37877));
    InMux I__6723 (
            .O(N__37881),
            .I(N__37873));
    InMux I__6722 (
            .O(N__37880),
            .I(N__37870));
    LocalMux I__6721 (
            .O(N__37877),
            .I(N__37867));
    InMux I__6720 (
            .O(N__37876),
            .I(N__37864));
    LocalMux I__6719 (
            .O(N__37873),
            .I(N__37857));
    LocalMux I__6718 (
            .O(N__37870),
            .I(N__37857));
    Span4Mux_v I__6717 (
            .O(N__37867),
            .I(N__37857));
    LocalMux I__6716 (
            .O(N__37864),
            .I(\c0.FRAME_MATCHER_state_16 ));
    Odrv4 I__6715 (
            .O(N__37857),
            .I(\c0.FRAME_MATCHER_state_16 ));
    InMux I__6714 (
            .O(N__37852),
            .I(N__37849));
    LocalMux I__6713 (
            .O(N__37849),
            .I(N__37843));
    InMux I__6712 (
            .O(N__37848),
            .I(N__37840));
    InMux I__6711 (
            .O(N__37847),
            .I(N__37837));
    InMux I__6710 (
            .O(N__37846),
            .I(N__37834));
    Span4Mux_h I__6709 (
            .O(N__37843),
            .I(N__37831));
    LocalMux I__6708 (
            .O(N__37840),
            .I(N__37828));
    LocalMux I__6707 (
            .O(N__37837),
            .I(\c0.FRAME_MATCHER_state_17 ));
    LocalMux I__6706 (
            .O(N__37834),
            .I(\c0.FRAME_MATCHER_state_17 ));
    Odrv4 I__6705 (
            .O(N__37831),
            .I(\c0.FRAME_MATCHER_state_17 ));
    Odrv4 I__6704 (
            .O(N__37828),
            .I(\c0.FRAME_MATCHER_state_17 ));
    InMux I__6703 (
            .O(N__37819),
            .I(N__37815));
    InMux I__6702 (
            .O(N__37818),
            .I(N__37812));
    LocalMux I__6701 (
            .O(N__37815),
            .I(N__37807));
    LocalMux I__6700 (
            .O(N__37812),
            .I(N__37807));
    Odrv4 I__6699 (
            .O(N__37807),
            .I(\c0.n21682 ));
    InMux I__6698 (
            .O(N__37804),
            .I(N__37800));
    CascadeMux I__6697 (
            .O(N__37803),
            .I(N__37796));
    LocalMux I__6696 (
            .O(N__37800),
            .I(N__37793));
    InMux I__6695 (
            .O(N__37799),
            .I(N__37790));
    InMux I__6694 (
            .O(N__37796),
            .I(N__37786));
    Span4Mux_h I__6693 (
            .O(N__37793),
            .I(N__37783));
    LocalMux I__6692 (
            .O(N__37790),
            .I(N__37780));
    InMux I__6691 (
            .O(N__37789),
            .I(N__37777));
    LocalMux I__6690 (
            .O(N__37786),
            .I(N__37774));
    Span4Mux_h I__6689 (
            .O(N__37783),
            .I(N__37769));
    Span4Mux_h I__6688 (
            .O(N__37780),
            .I(N__37769));
    LocalMux I__6687 (
            .O(N__37777),
            .I(\c0.FRAME_MATCHER_state_4 ));
    Odrv12 I__6686 (
            .O(N__37774),
            .I(\c0.FRAME_MATCHER_state_4 ));
    Odrv4 I__6685 (
            .O(N__37769),
            .I(\c0.FRAME_MATCHER_state_4 ));
    InMux I__6684 (
            .O(N__37762),
            .I(N__37759));
    LocalMux I__6683 (
            .O(N__37759),
            .I(N__37756));
    Odrv4 I__6682 (
            .O(N__37756),
            .I(\c0.n47 ));
    InMux I__6681 (
            .O(N__37753),
            .I(N__37747));
    InMux I__6680 (
            .O(N__37752),
            .I(N__37744));
    InMux I__6679 (
            .O(N__37751),
            .I(N__37741));
    InMux I__6678 (
            .O(N__37750),
            .I(N__37738));
    LocalMux I__6677 (
            .O(N__37747),
            .I(N__37735));
    LocalMux I__6676 (
            .O(N__37744),
            .I(\c0.FRAME_MATCHER_state_25 ));
    LocalMux I__6675 (
            .O(N__37741),
            .I(\c0.FRAME_MATCHER_state_25 ));
    LocalMux I__6674 (
            .O(N__37738),
            .I(\c0.FRAME_MATCHER_state_25 ));
    Odrv4 I__6673 (
            .O(N__37735),
            .I(\c0.FRAME_MATCHER_state_25 ));
    SRMux I__6672 (
            .O(N__37726),
            .I(N__37723));
    LocalMux I__6671 (
            .O(N__37723),
            .I(N__37720));
    Odrv12 I__6670 (
            .O(N__37720),
            .I(\c0.n21374 ));
    InMux I__6669 (
            .O(N__37717),
            .I(N__37711));
    InMux I__6668 (
            .O(N__37716),
            .I(N__37708));
    InMux I__6667 (
            .O(N__37715),
            .I(N__37703));
    InMux I__6666 (
            .O(N__37714),
            .I(N__37703));
    LocalMux I__6665 (
            .O(N__37711),
            .I(N__37698));
    LocalMux I__6664 (
            .O(N__37708),
            .I(N__37698));
    LocalMux I__6663 (
            .O(N__37703),
            .I(\c0.FRAME_MATCHER_state_10 ));
    Odrv4 I__6662 (
            .O(N__37698),
            .I(\c0.FRAME_MATCHER_state_10 ));
    SRMux I__6661 (
            .O(N__37693),
            .I(N__37690));
    LocalMux I__6660 (
            .O(N__37690),
            .I(\c0.n21348 ));
    InMux I__6659 (
            .O(N__37687),
            .I(N__37681));
    InMux I__6658 (
            .O(N__37686),
            .I(N__37676));
    InMux I__6657 (
            .O(N__37685),
            .I(N__37676));
    InMux I__6656 (
            .O(N__37684),
            .I(N__37673));
    LocalMux I__6655 (
            .O(N__37681),
            .I(N__37668));
    LocalMux I__6654 (
            .O(N__37676),
            .I(N__37668));
    LocalMux I__6653 (
            .O(N__37673),
            .I(\c0.FRAME_MATCHER_state_7 ));
    Odrv4 I__6652 (
            .O(N__37668),
            .I(\c0.FRAME_MATCHER_state_7 ));
    CascadeMux I__6651 (
            .O(N__37663),
            .I(\c0.n48_cascade_ ));
    InMux I__6650 (
            .O(N__37660),
            .I(N__37657));
    LocalMux I__6649 (
            .O(N__37657),
            .I(\c0.n45_adj_4413 ));
    CascadeMux I__6648 (
            .O(N__37654),
            .I(N__37650));
    InMux I__6647 (
            .O(N__37653),
            .I(N__37645));
    InMux I__6646 (
            .O(N__37650),
            .I(N__37645));
    LocalMux I__6645 (
            .O(N__37645),
            .I(N__37642));
    Span4Mux_v I__6644 (
            .O(N__37642),
            .I(N__37637));
    InMux I__6643 (
            .O(N__37641),
            .I(N__37634));
    InMux I__6642 (
            .O(N__37640),
            .I(N__37631));
    Sp12to4 I__6641 (
            .O(N__37637),
            .I(N__37628));
    LocalMux I__6640 (
            .O(N__37634),
            .I(\c0.FRAME_MATCHER_state_23 ));
    LocalMux I__6639 (
            .O(N__37631),
            .I(\c0.FRAME_MATCHER_state_23 ));
    Odrv12 I__6638 (
            .O(N__37628),
            .I(\c0.FRAME_MATCHER_state_23 ));
    InMux I__6637 (
            .O(N__37621),
            .I(N__37617));
    InMux I__6636 (
            .O(N__37620),
            .I(N__37614));
    LocalMux I__6635 (
            .O(N__37617),
            .I(\c0.n14_adj_4316 ));
    LocalMux I__6634 (
            .O(N__37614),
            .I(\c0.n14_adj_4316 ));
    InMux I__6633 (
            .O(N__37609),
            .I(N__37606));
    LocalMux I__6632 (
            .O(N__37606),
            .I(N__37600));
    InMux I__6631 (
            .O(N__37605),
            .I(N__37593));
    InMux I__6630 (
            .O(N__37604),
            .I(N__37593));
    InMux I__6629 (
            .O(N__37603),
            .I(N__37593));
    Odrv4 I__6628 (
            .O(N__37600),
            .I(\c0.FRAME_MATCHER_state_24 ));
    LocalMux I__6627 (
            .O(N__37593),
            .I(\c0.FRAME_MATCHER_state_24 ));
    SRMux I__6626 (
            .O(N__37588),
            .I(N__37585));
    LocalMux I__6625 (
            .O(N__37585),
            .I(\c0.n21372 ));
    SRMux I__6624 (
            .O(N__37582),
            .I(N__37579));
    LocalMux I__6623 (
            .O(N__37579),
            .I(N__37576));
    Span4Mux_h I__6622 (
            .O(N__37576),
            .I(N__37573));
    Odrv4 I__6621 (
            .O(N__37573),
            .I(\c0.n21346 ));
    SRMux I__6620 (
            .O(N__37570),
            .I(N__37567));
    LocalMux I__6619 (
            .O(N__37567),
            .I(N__37564));
    Span4Mux_v I__6618 (
            .O(N__37564),
            .I(N__37561));
    Span4Mux_h I__6617 (
            .O(N__37561),
            .I(N__37558));
    Odrv4 I__6616 (
            .O(N__37558),
            .I(\c0.n21364 ));
    CascadeMux I__6615 (
            .O(N__37555),
            .I(N__37552));
    InMux I__6614 (
            .O(N__37552),
            .I(N__37546));
    InMux I__6613 (
            .O(N__37551),
            .I(N__37546));
    LocalMux I__6612 (
            .O(N__37546),
            .I(N__37542));
    InMux I__6611 (
            .O(N__37545),
            .I(N__37538));
    Span4Mux_v I__6610 (
            .O(N__37542),
            .I(N__37535));
    InMux I__6609 (
            .O(N__37541),
            .I(N__37532));
    LocalMux I__6608 (
            .O(N__37538),
            .I(\c0.FRAME_MATCHER_state_9 ));
    Odrv4 I__6607 (
            .O(N__37535),
            .I(\c0.FRAME_MATCHER_state_9 ));
    LocalMux I__6606 (
            .O(N__37532),
            .I(\c0.FRAME_MATCHER_state_9 ));
    InMux I__6605 (
            .O(N__37525),
            .I(N__37522));
    LocalMux I__6604 (
            .O(N__37522),
            .I(\c0.n46 ));
    CascadeMux I__6603 (
            .O(N__37519),
            .I(N__37516));
    InMux I__6602 (
            .O(N__37516),
            .I(N__37510));
    InMux I__6601 (
            .O(N__37515),
            .I(N__37503));
    InMux I__6600 (
            .O(N__37514),
            .I(N__37503));
    InMux I__6599 (
            .O(N__37513),
            .I(N__37503));
    LocalMux I__6598 (
            .O(N__37510),
            .I(N__37496));
    LocalMux I__6597 (
            .O(N__37503),
            .I(N__37496));
    InMux I__6596 (
            .O(N__37502),
            .I(N__37489));
    InMux I__6595 (
            .O(N__37501),
            .I(N__37489));
    Span4Mux_h I__6594 (
            .O(N__37496),
            .I(N__37486));
    InMux I__6593 (
            .O(N__37495),
            .I(N__37481));
    InMux I__6592 (
            .O(N__37494),
            .I(N__37481));
    LocalMux I__6591 (
            .O(N__37489),
            .I(\c0.n117 ));
    Odrv4 I__6590 (
            .O(N__37486),
            .I(\c0.n117 ));
    LocalMux I__6589 (
            .O(N__37481),
            .I(\c0.n117 ));
    InMux I__6588 (
            .O(N__37474),
            .I(N__37459));
    InMux I__6587 (
            .O(N__37473),
            .I(N__37459));
    InMux I__6586 (
            .O(N__37472),
            .I(N__37459));
    InMux I__6585 (
            .O(N__37471),
            .I(N__37459));
    InMux I__6584 (
            .O(N__37470),
            .I(N__37454));
    InMux I__6583 (
            .O(N__37469),
            .I(N__37454));
    InMux I__6582 (
            .O(N__37468),
            .I(N__37451));
    LocalMux I__6581 (
            .O(N__37459),
            .I(N__37446));
    LocalMux I__6580 (
            .O(N__37454),
            .I(N__37446));
    LocalMux I__6579 (
            .O(N__37451),
            .I(N__37443));
    Span4Mux_h I__6578 (
            .O(N__37446),
            .I(N__37440));
    Odrv4 I__6577 (
            .O(N__37443),
            .I(\c0.n63_adj_4301 ));
    Odrv4 I__6576 (
            .O(N__37440),
            .I(\c0.n63_adj_4301 ));
    CascadeMux I__6575 (
            .O(N__37435),
            .I(\c0.n16958_cascade_ ));
    CascadeMux I__6574 (
            .O(N__37432),
            .I(N__37425));
    InMux I__6573 (
            .O(N__37431),
            .I(N__37415));
    InMux I__6572 (
            .O(N__37430),
            .I(N__37415));
    InMux I__6571 (
            .O(N__37429),
            .I(N__37415));
    InMux I__6570 (
            .O(N__37428),
            .I(N__37415));
    InMux I__6569 (
            .O(N__37425),
            .I(N__37410));
    InMux I__6568 (
            .O(N__37424),
            .I(N__37410));
    LocalMux I__6567 (
            .O(N__37415),
            .I(N__37404));
    LocalMux I__6566 (
            .O(N__37410),
            .I(N__37404));
    InMux I__6565 (
            .O(N__37409),
            .I(N__37401));
    Span4Mux_h I__6564 (
            .O(N__37404),
            .I(N__37398));
    LocalMux I__6563 (
            .O(N__37401),
            .I(\c0.n63 ));
    Odrv4 I__6562 (
            .O(N__37398),
            .I(\c0.n63 ));
    CascadeMux I__6561 (
            .O(N__37393),
            .I(\c0.n22695_cascade_ ));
    CascadeMux I__6560 (
            .O(N__37390),
            .I(N__37385));
    InMux I__6559 (
            .O(N__37389),
            .I(N__37382));
    InMux I__6558 (
            .O(N__37388),
            .I(N__37377));
    InMux I__6557 (
            .O(N__37385),
            .I(N__37377));
    LocalMux I__6556 (
            .O(N__37382),
            .I(\c0.FRAME_MATCHER_state_2 ));
    LocalMux I__6555 (
            .O(N__37377),
            .I(\c0.FRAME_MATCHER_state_2 ));
    CascadeMux I__6554 (
            .O(N__37372),
            .I(N__37369));
    InMux I__6553 (
            .O(N__37369),
            .I(N__37366));
    LocalMux I__6552 (
            .O(N__37366),
            .I(N__37363));
    Odrv4 I__6551 (
            .O(N__37363),
            .I(\c0.n13_adj_4388 ));
    InMux I__6550 (
            .O(N__37360),
            .I(N__37357));
    LocalMux I__6549 (
            .O(N__37357),
            .I(N__37353));
    InMux I__6548 (
            .O(N__37356),
            .I(N__37350));
    Odrv4 I__6547 (
            .O(N__37353),
            .I(\c0.n9207 ));
    LocalMux I__6546 (
            .O(N__37350),
            .I(\c0.n9207 ));
    InMux I__6545 (
            .O(N__37345),
            .I(N__37342));
    LocalMux I__6544 (
            .O(N__37342),
            .I(\c0.n14_adj_4337 ));
    CascadeMux I__6543 (
            .O(N__37339),
            .I(\c0.n7_adj_4352_cascade_ ));
    InMux I__6542 (
            .O(N__37336),
            .I(N__37331));
    CascadeMux I__6541 (
            .O(N__37335),
            .I(N__37328));
    InMux I__6540 (
            .O(N__37334),
            .I(N__37325));
    LocalMux I__6539 (
            .O(N__37331),
            .I(N__37322));
    InMux I__6538 (
            .O(N__37328),
            .I(N__37319));
    LocalMux I__6537 (
            .O(N__37325),
            .I(N__37313));
    Span4Mux_h I__6536 (
            .O(N__37322),
            .I(N__37313));
    LocalMux I__6535 (
            .O(N__37319),
            .I(N__37310));
    InMux I__6534 (
            .O(N__37318),
            .I(N__37307));
    Sp12to4 I__6533 (
            .O(N__37313),
            .I(N__37302));
    Span12Mux_v I__6532 (
            .O(N__37310),
            .I(N__37302));
    LocalMux I__6531 (
            .O(N__37307),
            .I(\c0.FRAME_MATCHER_state_26 ));
    Odrv12 I__6530 (
            .O(N__37302),
            .I(\c0.FRAME_MATCHER_state_26 ));
    InMux I__6529 (
            .O(N__37297),
            .I(N__37294));
    LocalMux I__6528 (
            .O(N__37294),
            .I(N__37291));
    Odrv4 I__6527 (
            .O(N__37291),
            .I(\c0.n21789 ));
    CascadeMux I__6526 (
            .O(N__37288),
            .I(\c0.n12996_cascade_ ));
    CascadeMux I__6525 (
            .O(N__37285),
            .I(\c0.n13020_cascade_ ));
    CascadeMux I__6524 (
            .O(N__37282),
            .I(\c0.data_out_frame_29_7_N_1483_1_cascade_ ));
    InMux I__6523 (
            .O(N__37279),
            .I(N__37276));
    LocalMux I__6522 (
            .O(N__37276),
            .I(\c0.n6650 ));
    CascadeMux I__6521 (
            .O(N__37273),
            .I(\c0.n6650_cascade_ ));
    InMux I__6520 (
            .O(N__37270),
            .I(N__37267));
    LocalMux I__6519 (
            .O(N__37267),
            .I(\c0.n6_adj_4270 ));
    CascadeMux I__6518 (
            .O(N__37264),
            .I(N__37260));
    InMux I__6517 (
            .O(N__37263),
            .I(N__37257));
    InMux I__6516 (
            .O(N__37260),
            .I(N__37254));
    LocalMux I__6515 (
            .O(N__37257),
            .I(N__37251));
    LocalMux I__6514 (
            .O(N__37254),
            .I(N__37247));
    Span4Mux_h I__6513 (
            .O(N__37251),
            .I(N__37243));
    InMux I__6512 (
            .O(N__37250),
            .I(N__37240));
    Span4Mux_h I__6511 (
            .O(N__37247),
            .I(N__37237));
    InMux I__6510 (
            .O(N__37246),
            .I(N__37234));
    Span4Mux_h I__6509 (
            .O(N__37243),
            .I(N__37231));
    LocalMux I__6508 (
            .O(N__37240),
            .I(encoder1_position_17));
    Odrv4 I__6507 (
            .O(N__37237),
            .I(encoder1_position_17));
    LocalMux I__6506 (
            .O(N__37234),
            .I(encoder1_position_17));
    Odrv4 I__6505 (
            .O(N__37231),
            .I(encoder1_position_17));
    CascadeMux I__6504 (
            .O(N__37222),
            .I(N__37218));
    InMux I__6503 (
            .O(N__37221),
            .I(N__37215));
    InMux I__6502 (
            .O(N__37218),
            .I(N__37212));
    LocalMux I__6501 (
            .O(N__37215),
            .I(data_out_frame_11_1));
    LocalMux I__6500 (
            .O(N__37212),
            .I(data_out_frame_11_1));
    CascadeMux I__6499 (
            .O(N__37207),
            .I(\c0.n9_adj_4415_cascade_ ));
    InMux I__6498 (
            .O(N__37204),
            .I(N__37200));
    InMux I__6497 (
            .O(N__37203),
            .I(N__37197));
    LocalMux I__6496 (
            .O(N__37200),
            .I(N__37194));
    LocalMux I__6495 (
            .O(N__37197),
            .I(N__37190));
    Span4Mux_v I__6494 (
            .O(N__37194),
            .I(N__37187));
    InMux I__6493 (
            .O(N__37193),
            .I(N__37184));
    Span12Mux_h I__6492 (
            .O(N__37190),
            .I(N__37181));
    Sp12to4 I__6491 (
            .O(N__37187),
            .I(N__37176));
    LocalMux I__6490 (
            .O(N__37184),
            .I(N__37176));
    Odrv12 I__6489 (
            .O(N__37181),
            .I(n14252));
    Odrv12 I__6488 (
            .O(N__37176),
            .I(n14252));
    InMux I__6487 (
            .O(N__37171),
            .I(N__37167));
    InMux I__6486 (
            .O(N__37170),
            .I(N__37164));
    LocalMux I__6485 (
            .O(N__37167),
            .I(N__37161));
    LocalMux I__6484 (
            .O(N__37164),
            .I(N__37158));
    Span4Mux_h I__6483 (
            .O(N__37161),
            .I(N__37155));
    Span4Mux_v I__6482 (
            .O(N__37158),
            .I(N__37152));
    Odrv4 I__6481 (
            .O(N__37155),
            .I(\c0.n38_adj_4387 ));
    Odrv4 I__6480 (
            .O(N__37152),
            .I(\c0.n38_adj_4387 ));
    InMux I__6479 (
            .O(N__37147),
            .I(N__37143));
    CascadeMux I__6478 (
            .O(N__37146),
            .I(N__37139));
    LocalMux I__6477 (
            .O(N__37143),
            .I(N__37136));
    InMux I__6476 (
            .O(N__37142),
            .I(N__37132));
    InMux I__6475 (
            .O(N__37139),
            .I(N__37129));
    Span4Mux_h I__6474 (
            .O(N__37136),
            .I(N__37126));
    InMux I__6473 (
            .O(N__37135),
            .I(N__37123));
    LocalMux I__6472 (
            .O(N__37132),
            .I(N__37118));
    LocalMux I__6471 (
            .O(N__37129),
            .I(N__37118));
    Odrv4 I__6470 (
            .O(N__37126),
            .I(\c0.tx_active ));
    LocalMux I__6469 (
            .O(N__37123),
            .I(\c0.tx_active ));
    Odrv12 I__6468 (
            .O(N__37118),
            .I(\c0.tx_active ));
    InMux I__6467 (
            .O(N__37111),
            .I(N__37108));
    LocalMux I__6466 (
            .O(N__37108),
            .I(\c0.n22651 ));
    CascadeMux I__6465 (
            .O(N__37105),
            .I(n22661_cascade_));
    InMux I__6464 (
            .O(N__37102),
            .I(N__37099));
    LocalMux I__6463 (
            .O(N__37099),
            .I(N__37095));
    InMux I__6462 (
            .O(N__37098),
            .I(N__37092));
    Span4Mux_h I__6461 (
            .O(N__37095),
            .I(N__37089));
    LocalMux I__6460 (
            .O(N__37092),
            .I(data_out_frame_7_3));
    Odrv4 I__6459 (
            .O(N__37089),
            .I(data_out_frame_7_3));
    InMux I__6458 (
            .O(N__37084),
            .I(N__37080));
    InMux I__6457 (
            .O(N__37083),
            .I(N__37077));
    LocalMux I__6456 (
            .O(N__37080),
            .I(data_out_frame_6_1));
    LocalMux I__6455 (
            .O(N__37077),
            .I(data_out_frame_6_1));
    CascadeMux I__6454 (
            .O(N__37072),
            .I(N__37068));
    CascadeMux I__6453 (
            .O(N__37071),
            .I(N__37065));
    InMux I__6452 (
            .O(N__37068),
            .I(N__37062));
    InMux I__6451 (
            .O(N__37065),
            .I(N__37057));
    LocalMux I__6450 (
            .O(N__37062),
            .I(N__37054));
    InMux I__6449 (
            .O(N__37061),
            .I(N__37051));
    InMux I__6448 (
            .O(N__37060),
            .I(N__37048));
    LocalMux I__6447 (
            .O(N__37057),
            .I(N__37043));
    Span4Mux_v I__6446 (
            .O(N__37054),
            .I(N__37036));
    LocalMux I__6445 (
            .O(N__37051),
            .I(N__37036));
    LocalMux I__6444 (
            .O(N__37048),
            .I(N__37036));
    InMux I__6443 (
            .O(N__37047),
            .I(N__37033));
    InMux I__6442 (
            .O(N__37046),
            .I(N__37030));
    Span4Mux_v I__6441 (
            .O(N__37043),
            .I(N__37025));
    Span4Mux_h I__6440 (
            .O(N__37036),
            .I(N__37025));
    LocalMux I__6439 (
            .O(N__37033),
            .I(encoder0_position_0));
    LocalMux I__6438 (
            .O(N__37030),
            .I(encoder0_position_0));
    Odrv4 I__6437 (
            .O(N__37025),
            .I(encoder0_position_0));
    InMux I__6436 (
            .O(N__37018),
            .I(N__37015));
    LocalMux I__6435 (
            .O(N__37015),
            .I(N__37011));
    InMux I__6434 (
            .O(N__37014),
            .I(N__37008));
    Span4Mux_v I__6433 (
            .O(N__37011),
            .I(N__37005));
    LocalMux I__6432 (
            .O(N__37008),
            .I(data_out_frame_9_0));
    Odrv4 I__6431 (
            .O(N__37005),
            .I(data_out_frame_9_0));
    InMux I__6430 (
            .O(N__37000),
            .I(N__36997));
    LocalMux I__6429 (
            .O(N__36997),
            .I(n2242));
    InMux I__6428 (
            .O(N__36994),
            .I(N__36990));
    InMux I__6427 (
            .O(N__36993),
            .I(N__36987));
    LocalMux I__6426 (
            .O(N__36990),
            .I(N__36982));
    LocalMux I__6425 (
            .O(N__36987),
            .I(N__36979));
    InMux I__6424 (
            .O(N__36986),
            .I(N__36974));
    InMux I__6423 (
            .O(N__36985),
            .I(N__36974));
    Span12Mux_v I__6422 (
            .O(N__36982),
            .I(N__36971));
    Span4Mux_v I__6421 (
            .O(N__36979),
            .I(N__36968));
    LocalMux I__6420 (
            .O(N__36974),
            .I(data_in_3_6));
    Odrv12 I__6419 (
            .O(N__36971),
            .I(data_in_3_6));
    Odrv4 I__6418 (
            .O(N__36968),
            .I(data_in_3_6));
    CascadeMux I__6417 (
            .O(N__36961),
            .I(N__36957));
    InMux I__6416 (
            .O(N__36960),
            .I(N__36952));
    InMux I__6415 (
            .O(N__36957),
            .I(N__36952));
    LocalMux I__6414 (
            .O(N__36952),
            .I(N__36949));
    Span4Mux_h I__6413 (
            .O(N__36949),
            .I(N__36944));
    InMux I__6412 (
            .O(N__36948),
            .I(N__36941));
    InMux I__6411 (
            .O(N__36947),
            .I(N__36938));
    Span4Mux_v I__6410 (
            .O(N__36944),
            .I(N__36933));
    LocalMux I__6409 (
            .O(N__36941),
            .I(N__36933));
    LocalMux I__6408 (
            .O(N__36938),
            .I(data_in_2_6));
    Odrv4 I__6407 (
            .O(N__36933),
            .I(data_in_2_6));
    InMux I__6406 (
            .O(N__36928),
            .I(N__36925));
    LocalMux I__6405 (
            .O(N__36925),
            .I(N__36921));
    InMux I__6404 (
            .O(N__36924),
            .I(N__36918));
    Span12Mux_v I__6403 (
            .O(N__36921),
            .I(N__36915));
    LocalMux I__6402 (
            .O(N__36918),
            .I(data_out_frame_10_1));
    Odrv12 I__6401 (
            .O(N__36915),
            .I(data_out_frame_10_1));
    CascadeMux I__6400 (
            .O(N__36910),
            .I(N__36903));
    InMux I__6399 (
            .O(N__36909),
            .I(N__36891));
    InMux I__6398 (
            .O(N__36908),
            .I(N__36884));
    InMux I__6397 (
            .O(N__36907),
            .I(N__36877));
    InMux I__6396 (
            .O(N__36906),
            .I(N__36877));
    InMux I__6395 (
            .O(N__36903),
            .I(N__36874));
    InMux I__6394 (
            .O(N__36902),
            .I(N__36867));
    CascadeMux I__6393 (
            .O(N__36901),
            .I(N__36864));
    CascadeMux I__6392 (
            .O(N__36900),
            .I(N__36859));
    InMux I__6391 (
            .O(N__36899),
            .I(N__36854));
    InMux I__6390 (
            .O(N__36898),
            .I(N__36854));
    InMux I__6389 (
            .O(N__36897),
            .I(N__36849));
    InMux I__6388 (
            .O(N__36896),
            .I(N__36849));
    InMux I__6387 (
            .O(N__36895),
            .I(N__36844));
    InMux I__6386 (
            .O(N__36894),
            .I(N__36841));
    LocalMux I__6385 (
            .O(N__36891),
            .I(N__36838));
    InMux I__6384 (
            .O(N__36890),
            .I(N__36835));
    InMux I__6383 (
            .O(N__36889),
            .I(N__36830));
    InMux I__6382 (
            .O(N__36888),
            .I(N__36825));
    InMux I__6381 (
            .O(N__36887),
            .I(N__36825));
    LocalMux I__6380 (
            .O(N__36884),
            .I(N__36822));
    InMux I__6379 (
            .O(N__36883),
            .I(N__36819));
    InMux I__6378 (
            .O(N__36882),
            .I(N__36814));
    LocalMux I__6377 (
            .O(N__36877),
            .I(N__36809));
    LocalMux I__6376 (
            .O(N__36874),
            .I(N__36809));
    InMux I__6375 (
            .O(N__36873),
            .I(N__36800));
    InMux I__6374 (
            .O(N__36872),
            .I(N__36800));
    InMux I__6373 (
            .O(N__36871),
            .I(N__36800));
    InMux I__6372 (
            .O(N__36870),
            .I(N__36800));
    LocalMux I__6371 (
            .O(N__36867),
            .I(N__36797));
    InMux I__6370 (
            .O(N__36864),
            .I(N__36788));
    InMux I__6369 (
            .O(N__36863),
            .I(N__36788));
    InMux I__6368 (
            .O(N__36862),
            .I(N__36788));
    InMux I__6367 (
            .O(N__36859),
            .I(N__36788));
    LocalMux I__6366 (
            .O(N__36854),
            .I(N__36783));
    LocalMux I__6365 (
            .O(N__36849),
            .I(N__36783));
    InMux I__6364 (
            .O(N__36848),
            .I(N__36778));
    InMux I__6363 (
            .O(N__36847),
            .I(N__36778));
    LocalMux I__6362 (
            .O(N__36844),
            .I(N__36769));
    LocalMux I__6361 (
            .O(N__36841),
            .I(N__36769));
    Span4Mux_v I__6360 (
            .O(N__36838),
            .I(N__36769));
    LocalMux I__6359 (
            .O(N__36835),
            .I(N__36769));
    InMux I__6358 (
            .O(N__36834),
            .I(N__36766));
    CascadeMux I__6357 (
            .O(N__36833),
            .I(N__36762));
    LocalMux I__6356 (
            .O(N__36830),
            .I(N__36756));
    LocalMux I__6355 (
            .O(N__36825),
            .I(N__36749));
    Span4Mux_v I__6354 (
            .O(N__36822),
            .I(N__36749));
    LocalMux I__6353 (
            .O(N__36819),
            .I(N__36749));
    InMux I__6352 (
            .O(N__36818),
            .I(N__36746));
    CascadeMux I__6351 (
            .O(N__36817),
            .I(N__36743));
    LocalMux I__6350 (
            .O(N__36814),
            .I(N__36738));
    Span4Mux_v I__6349 (
            .O(N__36809),
            .I(N__36733));
    LocalMux I__6348 (
            .O(N__36800),
            .I(N__36733));
    Span4Mux_v I__6347 (
            .O(N__36797),
            .I(N__36728));
    LocalMux I__6346 (
            .O(N__36788),
            .I(N__36728));
    Span4Mux_v I__6345 (
            .O(N__36783),
            .I(N__36721));
    LocalMux I__6344 (
            .O(N__36778),
            .I(N__36721));
    Span4Mux_h I__6343 (
            .O(N__36769),
            .I(N__36721));
    LocalMux I__6342 (
            .O(N__36766),
            .I(N__36718));
    InMux I__6341 (
            .O(N__36765),
            .I(N__36715));
    InMux I__6340 (
            .O(N__36762),
            .I(N__36712));
    InMux I__6339 (
            .O(N__36761),
            .I(N__36705));
    InMux I__6338 (
            .O(N__36760),
            .I(N__36705));
    InMux I__6337 (
            .O(N__36759),
            .I(N__36705));
    Span4Mux_v I__6336 (
            .O(N__36756),
            .I(N__36698));
    Span4Mux_v I__6335 (
            .O(N__36749),
            .I(N__36698));
    LocalMux I__6334 (
            .O(N__36746),
            .I(N__36698));
    InMux I__6333 (
            .O(N__36743),
            .I(N__36695));
    InMux I__6332 (
            .O(N__36742),
            .I(N__36692));
    InMux I__6331 (
            .O(N__36741),
            .I(N__36689));
    Span4Mux_v I__6330 (
            .O(N__36738),
            .I(N__36682));
    Span4Mux_v I__6329 (
            .O(N__36733),
            .I(N__36682));
    Span4Mux_v I__6328 (
            .O(N__36728),
            .I(N__36682));
    Span4Mux_h I__6327 (
            .O(N__36721),
            .I(N__36679));
    Span4Mux_h I__6326 (
            .O(N__36718),
            .I(N__36676));
    LocalMux I__6325 (
            .O(N__36715),
            .I(N__36665));
    LocalMux I__6324 (
            .O(N__36712),
            .I(N__36665));
    LocalMux I__6323 (
            .O(N__36705),
            .I(N__36665));
    Sp12to4 I__6322 (
            .O(N__36698),
            .I(N__36665));
    LocalMux I__6321 (
            .O(N__36695),
            .I(N__36665));
    LocalMux I__6320 (
            .O(N__36692),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__6319 (
            .O(N__36689),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__6318 (
            .O(N__36682),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__6317 (
            .O(N__36679),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__6316 (
            .O(N__36676),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv12 I__6315 (
            .O(N__36665),
            .I(\c0.byte_transmit_counter_1 ));
    InMux I__6314 (
            .O(N__36652),
            .I(N__36649));
    LocalMux I__6313 (
            .O(N__36649),
            .I(\c0.n24183 ));
    InMux I__6312 (
            .O(N__36646),
            .I(N__36638));
    InMux I__6311 (
            .O(N__36645),
            .I(N__36638));
    InMux I__6310 (
            .O(N__36644),
            .I(N__36633));
    InMux I__6309 (
            .O(N__36643),
            .I(N__36633));
    LocalMux I__6308 (
            .O(N__36638),
            .I(N__36630));
    LocalMux I__6307 (
            .O(N__36633),
            .I(data_in_3_7));
    Odrv12 I__6306 (
            .O(N__36630),
            .I(data_in_3_7));
    InMux I__6305 (
            .O(N__36625),
            .I(N__36620));
    InMux I__6304 (
            .O(N__36624),
            .I(N__36617));
    InMux I__6303 (
            .O(N__36623),
            .I(N__36614));
    LocalMux I__6302 (
            .O(N__36620),
            .I(N__36611));
    LocalMux I__6301 (
            .O(N__36617),
            .I(N__36608));
    LocalMux I__6300 (
            .O(N__36614),
            .I(N__36605));
    Span4Mux_h I__6299 (
            .O(N__36611),
            .I(N__36600));
    Span4Mux_v I__6298 (
            .O(N__36608),
            .I(N__36600));
    Odrv4 I__6297 (
            .O(N__36605),
            .I(data_in_2_7));
    Odrv4 I__6296 (
            .O(N__36600),
            .I(data_in_2_7));
    InMux I__6295 (
            .O(N__36595),
            .I(N__36591));
    InMux I__6294 (
            .O(N__36594),
            .I(N__36588));
    LocalMux I__6293 (
            .O(N__36591),
            .I(N__36583));
    LocalMux I__6292 (
            .O(N__36588),
            .I(N__36580));
    InMux I__6291 (
            .O(N__36587),
            .I(N__36577));
    InMux I__6290 (
            .O(N__36586),
            .I(N__36574));
    Span4Mux_h I__6289 (
            .O(N__36583),
            .I(N__36571));
    Span4Mux_v I__6288 (
            .O(N__36580),
            .I(N__36566));
    LocalMux I__6287 (
            .O(N__36577),
            .I(N__36566));
    LocalMux I__6286 (
            .O(N__36574),
            .I(data_in_3_2));
    Odrv4 I__6285 (
            .O(N__36571),
            .I(data_in_3_2));
    Odrv4 I__6284 (
            .O(N__36566),
            .I(data_in_3_2));
    InMux I__6283 (
            .O(N__36559),
            .I(N__36553));
    InMux I__6282 (
            .O(N__36558),
            .I(N__36550));
    CascadeMux I__6281 (
            .O(N__36557),
            .I(N__36546));
    CascadeMux I__6280 (
            .O(N__36556),
            .I(N__36543));
    LocalMux I__6279 (
            .O(N__36553),
            .I(N__36540));
    LocalMux I__6278 (
            .O(N__36550),
            .I(N__36537));
    InMux I__6277 (
            .O(N__36549),
            .I(N__36532));
    InMux I__6276 (
            .O(N__36546),
            .I(N__36532));
    InMux I__6275 (
            .O(N__36543),
            .I(N__36527));
    Span4Mux_v I__6274 (
            .O(N__36540),
            .I(N__36522));
    Span4Mux_h I__6273 (
            .O(N__36537),
            .I(N__36522));
    LocalMux I__6272 (
            .O(N__36532),
            .I(N__36519));
    InMux I__6271 (
            .O(N__36531),
            .I(N__36514));
    InMux I__6270 (
            .O(N__36530),
            .I(N__36514));
    LocalMux I__6269 (
            .O(N__36527),
            .I(encoder0_position_17));
    Odrv4 I__6268 (
            .O(N__36522),
            .I(encoder0_position_17));
    Odrv4 I__6267 (
            .O(N__36519),
            .I(encoder0_position_17));
    LocalMux I__6266 (
            .O(N__36514),
            .I(encoder0_position_17));
    CascadeMux I__6265 (
            .O(N__36505),
            .I(N__36500));
    InMux I__6264 (
            .O(N__36504),
            .I(N__36496));
    CascadeMux I__6263 (
            .O(N__36503),
            .I(N__36492));
    InMux I__6262 (
            .O(N__36500),
            .I(N__36489));
    InMux I__6261 (
            .O(N__36499),
            .I(N__36486));
    LocalMux I__6260 (
            .O(N__36496),
            .I(N__36483));
    InMux I__6259 (
            .O(N__36495),
            .I(N__36480));
    InMux I__6258 (
            .O(N__36492),
            .I(N__36477));
    LocalMux I__6257 (
            .O(N__36489),
            .I(N__36472));
    LocalMux I__6256 (
            .O(N__36486),
            .I(N__36472));
    Span4Mux_h I__6255 (
            .O(N__36483),
            .I(N__36469));
    LocalMux I__6254 (
            .O(N__36480),
            .I(encoder1_position_28));
    LocalMux I__6253 (
            .O(N__36477),
            .I(encoder1_position_28));
    Odrv12 I__6252 (
            .O(N__36472),
            .I(encoder1_position_28));
    Odrv4 I__6251 (
            .O(N__36469),
            .I(encoder1_position_28));
    CascadeMux I__6250 (
            .O(N__36460),
            .I(N__36455));
    InMux I__6249 (
            .O(N__36459),
            .I(N__36451));
    InMux I__6248 (
            .O(N__36458),
            .I(N__36446));
    InMux I__6247 (
            .O(N__36455),
            .I(N__36446));
    InMux I__6246 (
            .O(N__36454),
            .I(N__36443));
    LocalMux I__6245 (
            .O(N__36451),
            .I(N__36440));
    LocalMux I__6244 (
            .O(N__36446),
            .I(N__36433));
    LocalMux I__6243 (
            .O(N__36443),
            .I(N__36433));
    Span4Mux_h I__6242 (
            .O(N__36440),
            .I(N__36433));
    Span4Mux_h I__6241 (
            .O(N__36433),
            .I(N__36430));
    Odrv4 I__6240 (
            .O(N__36430),
            .I(\c0.n13338 ));
    InMux I__6239 (
            .O(N__36427),
            .I(N__36422));
    InMux I__6238 (
            .O(N__36426),
            .I(N__36419));
    CascadeMux I__6237 (
            .O(N__36425),
            .I(N__36416));
    LocalMux I__6236 (
            .O(N__36422),
            .I(N__36413));
    LocalMux I__6235 (
            .O(N__36419),
            .I(N__36410));
    InMux I__6234 (
            .O(N__36416),
            .I(N__36407));
    Span4Mux_h I__6233 (
            .O(N__36413),
            .I(N__36403));
    Span4Mux_h I__6232 (
            .O(N__36410),
            .I(N__36398));
    LocalMux I__6231 (
            .O(N__36407),
            .I(N__36398));
    InMux I__6230 (
            .O(N__36406),
            .I(N__36395));
    Span4Mux_v I__6229 (
            .O(N__36403),
            .I(N__36392));
    Span4Mux_v I__6228 (
            .O(N__36398),
            .I(N__36389));
    LocalMux I__6227 (
            .O(N__36395),
            .I(data_in_2_5));
    Odrv4 I__6226 (
            .O(N__36392),
            .I(data_in_2_5));
    Odrv4 I__6225 (
            .O(N__36389),
            .I(data_in_2_5));
    InMux I__6224 (
            .O(N__36382),
            .I(N__36378));
    InMux I__6223 (
            .O(N__36381),
            .I(N__36374));
    LocalMux I__6222 (
            .O(N__36378),
            .I(N__36371));
    InMux I__6221 (
            .O(N__36377),
            .I(N__36368));
    LocalMux I__6220 (
            .O(N__36374),
            .I(N__36364));
    Span4Mux_h I__6219 (
            .O(N__36371),
            .I(N__36359));
    LocalMux I__6218 (
            .O(N__36368),
            .I(N__36359));
    InMux I__6217 (
            .O(N__36367),
            .I(N__36356));
    Span4Mux_v I__6216 (
            .O(N__36364),
            .I(N__36353));
    Span4Mux_v I__6215 (
            .O(N__36359),
            .I(N__36350));
    LocalMux I__6214 (
            .O(N__36356),
            .I(data_in_1_3));
    Odrv4 I__6213 (
            .O(N__36353),
            .I(data_in_1_3));
    Odrv4 I__6212 (
            .O(N__36350),
            .I(data_in_1_3));
    InMux I__6211 (
            .O(N__36343),
            .I(N__36340));
    LocalMux I__6210 (
            .O(N__36340),
            .I(N__36337));
    Span4Mux_h I__6209 (
            .O(N__36337),
            .I(N__36334));
    Odrv4 I__6208 (
            .O(N__36334),
            .I(\c0.n16_adj_4478 ));
    InMux I__6207 (
            .O(N__36331),
            .I(N__36328));
    LocalMux I__6206 (
            .O(N__36328),
            .I(N__36325));
    Span4Mux_h I__6205 (
            .O(N__36325),
            .I(N__36320));
    InMux I__6204 (
            .O(N__36324),
            .I(N__36315));
    InMux I__6203 (
            .O(N__36323),
            .I(N__36315));
    Odrv4 I__6202 (
            .O(N__36320),
            .I(data_in_1_1));
    LocalMux I__6201 (
            .O(N__36315),
            .I(data_in_1_1));
    CascadeMux I__6200 (
            .O(N__36310),
            .I(N__36307));
    InMux I__6199 (
            .O(N__36307),
            .I(N__36304));
    LocalMux I__6198 (
            .O(N__36304),
            .I(N__36301));
    Span4Mux_h I__6197 (
            .O(N__36301),
            .I(N__36296));
    InMux I__6196 (
            .O(N__36300),
            .I(N__36291));
    InMux I__6195 (
            .O(N__36299),
            .I(N__36291));
    Odrv4 I__6194 (
            .O(N__36296),
            .I(data_in_0_1));
    LocalMux I__6193 (
            .O(N__36291),
            .I(data_in_0_1));
    InMux I__6192 (
            .O(N__36286),
            .I(N__36282));
    InMux I__6191 (
            .O(N__36285),
            .I(N__36279));
    LocalMux I__6190 (
            .O(N__36282),
            .I(N__36276));
    LocalMux I__6189 (
            .O(N__36279),
            .I(data_out_frame_6_5));
    Odrv12 I__6188 (
            .O(N__36276),
            .I(data_out_frame_6_5));
    InMux I__6187 (
            .O(N__36271),
            .I(N__36268));
    LocalMux I__6186 (
            .O(N__36268),
            .I(n2256));
    CascadeMux I__6185 (
            .O(N__36265),
            .I(N__36262));
    InMux I__6184 (
            .O(N__36262),
            .I(N__36259));
    LocalMux I__6183 (
            .O(N__36259),
            .I(N__36253));
    InMux I__6182 (
            .O(N__36258),
            .I(N__36249));
    CascadeMux I__6181 (
            .O(N__36257),
            .I(N__36246));
    InMux I__6180 (
            .O(N__36256),
            .I(N__36243));
    Span4Mux_h I__6179 (
            .O(N__36253),
            .I(N__36240));
    InMux I__6178 (
            .O(N__36252),
            .I(N__36237));
    LocalMux I__6177 (
            .O(N__36249),
            .I(N__36234));
    InMux I__6176 (
            .O(N__36246),
            .I(N__36231));
    LocalMux I__6175 (
            .O(N__36243),
            .I(encoder0_position_15));
    Odrv4 I__6174 (
            .O(N__36240),
            .I(encoder0_position_15));
    LocalMux I__6173 (
            .O(N__36237),
            .I(encoder0_position_15));
    Odrv12 I__6172 (
            .O(N__36234),
            .I(encoder0_position_15));
    LocalMux I__6171 (
            .O(N__36231),
            .I(encoder0_position_15));
    InMux I__6170 (
            .O(N__36220),
            .I(N__36217));
    LocalMux I__6169 (
            .O(N__36217),
            .I(N__36213));
    CascadeMux I__6168 (
            .O(N__36216),
            .I(N__36210));
    Span4Mux_v I__6167 (
            .O(N__36213),
            .I(N__36207));
    InMux I__6166 (
            .O(N__36210),
            .I(N__36204));
    Span4Mux_h I__6165 (
            .O(N__36207),
            .I(N__36201));
    LocalMux I__6164 (
            .O(N__36204),
            .I(N__36198));
    Span4Mux_h I__6163 (
            .O(N__36201),
            .I(N__36193));
    Span4Mux_h I__6162 (
            .O(N__36198),
            .I(N__36190));
    InMux I__6161 (
            .O(N__36197),
            .I(N__36185));
    InMux I__6160 (
            .O(N__36196),
            .I(N__36185));
    Odrv4 I__6159 (
            .O(N__36193),
            .I(data_in_2_0));
    Odrv4 I__6158 (
            .O(N__36190),
            .I(data_in_2_0));
    LocalMux I__6157 (
            .O(N__36185),
            .I(data_in_2_0));
    InMux I__6156 (
            .O(N__36178),
            .I(N__36175));
    LocalMux I__6155 (
            .O(N__36175),
            .I(n2247));
    InMux I__6154 (
            .O(N__36172),
            .I(N__36169));
    LocalMux I__6153 (
            .O(N__36169),
            .I(n2265));
    InMux I__6152 (
            .O(N__36166),
            .I(N__36160));
    InMux I__6151 (
            .O(N__36165),
            .I(N__36160));
    LocalMux I__6150 (
            .O(N__36160),
            .I(N__36156));
    InMux I__6149 (
            .O(N__36159),
            .I(N__36151));
    Span4Mux_h I__6148 (
            .O(N__36156),
            .I(N__36148));
    InMux I__6147 (
            .O(N__36155),
            .I(N__36143));
    InMux I__6146 (
            .O(N__36154),
            .I(N__36143));
    LocalMux I__6145 (
            .O(N__36151),
            .I(encoder0_position_6));
    Odrv4 I__6144 (
            .O(N__36148),
            .I(encoder0_position_6));
    LocalMux I__6143 (
            .O(N__36143),
            .I(encoder0_position_6));
    CascadeMux I__6142 (
            .O(N__36136),
            .I(N__36133));
    InMux I__6141 (
            .O(N__36133),
            .I(N__36130));
    LocalMux I__6140 (
            .O(N__36130),
            .I(N__36127));
    Span4Mux_v I__6139 (
            .O(N__36127),
            .I(N__36124));
    Span4Mux_h I__6138 (
            .O(N__36124),
            .I(N__36118));
    InMux I__6137 (
            .O(N__36123),
            .I(N__36115));
    InMux I__6136 (
            .O(N__36122),
            .I(N__36112));
    InMux I__6135 (
            .O(N__36121),
            .I(N__36108));
    Span4Mux_h I__6134 (
            .O(N__36118),
            .I(N__36105));
    LocalMux I__6133 (
            .O(N__36115),
            .I(N__36100));
    LocalMux I__6132 (
            .O(N__36112),
            .I(N__36100));
    InMux I__6131 (
            .O(N__36111),
            .I(N__36097));
    LocalMux I__6130 (
            .O(N__36108),
            .I(encoder0_position_20));
    Odrv4 I__6129 (
            .O(N__36105),
            .I(encoder0_position_20));
    Odrv4 I__6128 (
            .O(N__36100),
            .I(encoder0_position_20));
    LocalMux I__6127 (
            .O(N__36097),
            .I(encoder0_position_20));
    InMux I__6126 (
            .O(N__36088),
            .I(N__36085));
    LocalMux I__6125 (
            .O(N__36085),
            .I(n2266));
    CascadeMux I__6124 (
            .O(N__36082),
            .I(N__36079));
    InMux I__6123 (
            .O(N__36079),
            .I(N__36075));
    CascadeMux I__6122 (
            .O(N__36078),
            .I(N__36072));
    LocalMux I__6121 (
            .O(N__36075),
            .I(N__36069));
    InMux I__6120 (
            .O(N__36072),
            .I(N__36066));
    Span4Mux_h I__6119 (
            .O(N__36069),
            .I(N__36063));
    LocalMux I__6118 (
            .O(N__36066),
            .I(N__36059));
    Span4Mux_h I__6117 (
            .O(N__36063),
            .I(N__36053));
    InMux I__6116 (
            .O(N__36062),
            .I(N__36050));
    Span4Mux_h I__6115 (
            .O(N__36059),
            .I(N__36047));
    InMux I__6114 (
            .O(N__36058),
            .I(N__36044));
    InMux I__6113 (
            .O(N__36057),
            .I(N__36039));
    InMux I__6112 (
            .O(N__36056),
            .I(N__36039));
    Odrv4 I__6111 (
            .O(N__36053),
            .I(encoder0_position_5));
    LocalMux I__6110 (
            .O(N__36050),
            .I(encoder0_position_5));
    Odrv4 I__6109 (
            .O(N__36047),
            .I(encoder0_position_5));
    LocalMux I__6108 (
            .O(N__36044),
            .I(encoder0_position_5));
    LocalMux I__6107 (
            .O(N__36039),
            .I(encoder0_position_5));
    InMux I__6106 (
            .O(N__36028),
            .I(N__36024));
    InMux I__6105 (
            .O(N__36027),
            .I(N__36021));
    LocalMux I__6104 (
            .O(N__36024),
            .I(N__36018));
    LocalMux I__6103 (
            .O(N__36021),
            .I(N__36015));
    Odrv12 I__6102 (
            .O(N__36018),
            .I(\c0.n21808 ));
    Odrv4 I__6101 (
            .O(N__36015),
            .I(\c0.n21808 ));
    InMux I__6100 (
            .O(N__36010),
            .I(N__36007));
    LocalMux I__6099 (
            .O(N__36007),
            .I(n2250));
    CascadeMux I__6098 (
            .O(N__36004),
            .I(N__36001));
    InMux I__6097 (
            .O(N__36001),
            .I(N__35998));
    LocalMux I__6096 (
            .O(N__35998),
            .I(N__35994));
    InMux I__6095 (
            .O(N__35997),
            .I(N__35990));
    Span4Mux_h I__6094 (
            .O(N__35994),
            .I(N__35986));
    CascadeMux I__6093 (
            .O(N__35993),
            .I(N__35983));
    LocalMux I__6092 (
            .O(N__35990),
            .I(N__35980));
    InMux I__6091 (
            .O(N__35989),
            .I(N__35976));
    Span4Mux_h I__6090 (
            .O(N__35986),
            .I(N__35973));
    InMux I__6089 (
            .O(N__35983),
            .I(N__35970));
    Span4Mux_h I__6088 (
            .O(N__35980),
            .I(N__35967));
    InMux I__6087 (
            .O(N__35979),
            .I(N__35964));
    LocalMux I__6086 (
            .O(N__35976),
            .I(encoder0_position_21));
    Odrv4 I__6085 (
            .O(N__35973),
            .I(encoder0_position_21));
    LocalMux I__6084 (
            .O(N__35970),
            .I(encoder0_position_21));
    Odrv4 I__6083 (
            .O(N__35967),
            .I(encoder0_position_21));
    LocalMux I__6082 (
            .O(N__35964),
            .I(encoder0_position_21));
    InMux I__6081 (
            .O(N__35953),
            .I(N__35950));
    LocalMux I__6080 (
            .O(N__35950),
            .I(n2262));
    InMux I__6079 (
            .O(N__35947),
            .I(N__35944));
    LocalMux I__6078 (
            .O(N__35944),
            .I(N__35941));
    Odrv12 I__6077 (
            .O(N__35941),
            .I(n2260));
    InMux I__6076 (
            .O(N__35938),
            .I(N__35935));
    LocalMux I__6075 (
            .O(N__35935),
            .I(n2254));
    InMux I__6074 (
            .O(N__35932),
            .I(N__35929));
    LocalMux I__6073 (
            .O(N__35929),
            .I(N__35925));
    InMux I__6072 (
            .O(N__35928),
            .I(N__35922));
    Span4Mux_h I__6071 (
            .O(N__35925),
            .I(N__35919));
    LocalMux I__6070 (
            .O(N__35922),
            .I(N__35916));
    Odrv4 I__6069 (
            .O(N__35919),
            .I(\c0.n10394 ));
    Odrv12 I__6068 (
            .O(N__35916),
            .I(\c0.n10394 ));
    InMux I__6067 (
            .O(N__35911),
            .I(N__35908));
    LocalMux I__6066 (
            .O(N__35908),
            .I(N__35905));
    Span4Mux_h I__6065 (
            .O(N__35905),
            .I(N__35902));
    Odrv4 I__6064 (
            .O(N__35902),
            .I(\c0.n20328 ));
    CascadeMux I__6063 (
            .O(N__35899),
            .I(N__35896));
    InMux I__6062 (
            .O(N__35896),
            .I(N__35892));
    InMux I__6061 (
            .O(N__35895),
            .I(N__35887));
    LocalMux I__6060 (
            .O(N__35892),
            .I(N__35884));
    InMux I__6059 (
            .O(N__35891),
            .I(N__35881));
    CascadeMux I__6058 (
            .O(N__35890),
            .I(N__35878));
    LocalMux I__6057 (
            .O(N__35887),
            .I(N__35874));
    Span4Mux_h I__6056 (
            .O(N__35884),
            .I(N__35869));
    LocalMux I__6055 (
            .O(N__35881),
            .I(N__35866));
    InMux I__6054 (
            .O(N__35878),
            .I(N__35861));
    InMux I__6053 (
            .O(N__35877),
            .I(N__35861));
    Span4Mux_h I__6052 (
            .O(N__35874),
            .I(N__35858));
    InMux I__6051 (
            .O(N__35873),
            .I(N__35853));
    InMux I__6050 (
            .O(N__35872),
            .I(N__35853));
    Odrv4 I__6049 (
            .O(N__35869),
            .I(encoder0_position_14));
    Odrv4 I__6048 (
            .O(N__35866),
            .I(encoder0_position_14));
    LocalMux I__6047 (
            .O(N__35861),
            .I(encoder0_position_14));
    Odrv4 I__6046 (
            .O(N__35858),
            .I(encoder0_position_14));
    LocalMux I__6045 (
            .O(N__35853),
            .I(encoder0_position_14));
    CascadeMux I__6044 (
            .O(N__35842),
            .I(\c0.n20328_cascade_ ));
    InMux I__6043 (
            .O(N__35839),
            .I(N__35836));
    LocalMux I__6042 (
            .O(N__35836),
            .I(N__35833));
    Span4Mux_h I__6041 (
            .O(N__35833),
            .I(N__35830));
    Odrv4 I__6040 (
            .O(N__35830),
            .I(\c0.n22367 ));
    CascadeMux I__6039 (
            .O(N__35827),
            .I(\c0.n22367_cascade_ ));
    InMux I__6038 (
            .O(N__35824),
            .I(N__35821));
    LocalMux I__6037 (
            .O(N__35821),
            .I(\c0.n23569 ));
    InMux I__6036 (
            .O(N__35818),
            .I(N__35815));
    LocalMux I__6035 (
            .O(N__35815),
            .I(n2271));
    InMux I__6034 (
            .O(N__35812),
            .I(N__35807));
    InMux I__6033 (
            .O(N__35811),
            .I(N__35804));
    InMux I__6032 (
            .O(N__35810),
            .I(N__35801));
    LocalMux I__6031 (
            .O(N__35807),
            .I(\c0.n10_adj_4331 ));
    LocalMux I__6030 (
            .O(N__35804),
            .I(\c0.n10_adj_4331 ));
    LocalMux I__6029 (
            .O(N__35801),
            .I(\c0.n10_adj_4331 ));
    CascadeMux I__6028 (
            .O(N__35794),
            .I(N__35791));
    InMux I__6027 (
            .O(N__35791),
            .I(N__35788));
    LocalMux I__6026 (
            .O(N__35788),
            .I(N__35784));
    InMux I__6025 (
            .O(N__35787),
            .I(N__35781));
    Odrv12 I__6024 (
            .O(N__35784),
            .I(\c0.n22230 ));
    LocalMux I__6023 (
            .O(N__35781),
            .I(\c0.n22230 ));
    CascadeMux I__6022 (
            .O(N__35776),
            .I(N__35773));
    InMux I__6021 (
            .O(N__35773),
            .I(N__35769));
    InMux I__6020 (
            .O(N__35772),
            .I(N__35766));
    LocalMux I__6019 (
            .O(N__35769),
            .I(N__35759));
    LocalMux I__6018 (
            .O(N__35766),
            .I(N__35756));
    InMux I__6017 (
            .O(N__35765),
            .I(N__35753));
    InMux I__6016 (
            .O(N__35764),
            .I(N__35750));
    InMux I__6015 (
            .O(N__35763),
            .I(N__35747));
    InMux I__6014 (
            .O(N__35762),
            .I(N__35744));
    Span4Mux_v I__6013 (
            .O(N__35759),
            .I(N__35739));
    Span4Mux_h I__6012 (
            .O(N__35756),
            .I(N__35739));
    LocalMux I__6011 (
            .O(N__35753),
            .I(encoder0_position_1));
    LocalMux I__6010 (
            .O(N__35750),
            .I(encoder0_position_1));
    LocalMux I__6009 (
            .O(N__35747),
            .I(encoder0_position_1));
    LocalMux I__6008 (
            .O(N__35744),
            .I(encoder0_position_1));
    Odrv4 I__6007 (
            .O(N__35739),
            .I(encoder0_position_1));
    CascadeMux I__6006 (
            .O(N__35728),
            .I(\c0.n22461_cascade_ ));
    InMux I__6005 (
            .O(N__35725),
            .I(N__35720));
    CascadeMux I__6004 (
            .O(N__35724),
            .I(N__35717));
    InMux I__6003 (
            .O(N__35723),
            .I(N__35714));
    LocalMux I__6002 (
            .O(N__35720),
            .I(N__35710));
    InMux I__6001 (
            .O(N__35717),
            .I(N__35707));
    LocalMux I__6000 (
            .O(N__35714),
            .I(N__35704));
    InMux I__5999 (
            .O(N__35713),
            .I(N__35698));
    Span12Mux_h I__5998 (
            .O(N__35710),
            .I(N__35695));
    LocalMux I__5997 (
            .O(N__35707),
            .I(N__35690));
    Span4Mux_h I__5996 (
            .O(N__35704),
            .I(N__35690));
    InMux I__5995 (
            .O(N__35703),
            .I(N__35687));
    InMux I__5994 (
            .O(N__35702),
            .I(N__35684));
    InMux I__5993 (
            .O(N__35701),
            .I(N__35681));
    LocalMux I__5992 (
            .O(N__35698),
            .I(encoder0_position_13));
    Odrv12 I__5991 (
            .O(N__35695),
            .I(encoder0_position_13));
    Odrv4 I__5990 (
            .O(N__35690),
            .I(encoder0_position_13));
    LocalMux I__5989 (
            .O(N__35687),
            .I(encoder0_position_13));
    LocalMux I__5988 (
            .O(N__35684),
            .I(encoder0_position_13));
    LocalMux I__5987 (
            .O(N__35681),
            .I(encoder0_position_13));
    InMux I__5986 (
            .O(N__35668),
            .I(N__35665));
    LocalMux I__5985 (
            .O(N__35665),
            .I(N__35662));
    Odrv4 I__5984 (
            .O(N__35662),
            .I(\c0.n20_adj_4318 ));
    CascadeMux I__5983 (
            .O(N__35659),
            .I(N__35656));
    InMux I__5982 (
            .O(N__35656),
            .I(N__35652));
    CascadeMux I__5981 (
            .O(N__35655),
            .I(N__35649));
    LocalMux I__5980 (
            .O(N__35652),
            .I(N__35646));
    InMux I__5979 (
            .O(N__35649),
            .I(N__35641));
    Span4Mux_h I__5978 (
            .O(N__35646),
            .I(N__35638));
    InMux I__5977 (
            .O(N__35645),
            .I(N__35635));
    InMux I__5976 (
            .O(N__35644),
            .I(N__35632));
    LocalMux I__5975 (
            .O(N__35641),
            .I(N__35629));
    Sp12to4 I__5974 (
            .O(N__35638),
            .I(N__35624));
    LocalMux I__5973 (
            .O(N__35635),
            .I(N__35624));
    LocalMux I__5972 (
            .O(N__35632),
            .I(N__35619));
    Span4Mux_h I__5971 (
            .O(N__35629),
            .I(N__35619));
    Odrv12 I__5970 (
            .O(N__35624),
            .I(encoder1_position_26));
    Odrv4 I__5969 (
            .O(N__35619),
            .I(encoder1_position_26));
    InMux I__5968 (
            .O(N__35614),
            .I(N__35611));
    LocalMux I__5967 (
            .O(N__35611),
            .I(N__35606));
    InMux I__5966 (
            .O(N__35610),
            .I(N__35600));
    InMux I__5965 (
            .O(N__35609),
            .I(N__35600));
    Span4Mux_v I__5964 (
            .O(N__35606),
            .I(N__35597));
    InMux I__5963 (
            .O(N__35605),
            .I(N__35594));
    LocalMux I__5962 (
            .O(N__35600),
            .I(N__35591));
    Span4Mux_h I__5961 (
            .O(N__35597),
            .I(N__35587));
    LocalMux I__5960 (
            .O(N__35594),
            .I(N__35582));
    Span4Mux_h I__5959 (
            .O(N__35591),
            .I(N__35582));
    InMux I__5958 (
            .O(N__35590),
            .I(N__35579));
    Odrv4 I__5957 (
            .O(N__35587),
            .I(\c0.n20236 ));
    Odrv4 I__5956 (
            .O(N__35582),
            .I(\c0.n20236 ));
    LocalMux I__5955 (
            .O(N__35579),
            .I(\c0.n20236 ));
    InMux I__5954 (
            .O(N__35572),
            .I(N__35569));
    LocalMux I__5953 (
            .O(N__35569),
            .I(N__35565));
    InMux I__5952 (
            .O(N__35568),
            .I(N__35562));
    Span4Mux_h I__5951 (
            .O(N__35565),
            .I(N__35559));
    LocalMux I__5950 (
            .O(N__35562),
            .I(N__35556));
    Span4Mux_v I__5949 (
            .O(N__35559),
            .I(N__35553));
    Span4Mux_v I__5948 (
            .O(N__35556),
            .I(N__35550));
    Odrv4 I__5947 (
            .O(N__35553),
            .I(\c0.n22449 ));
    Odrv4 I__5946 (
            .O(N__35550),
            .I(\c0.n22449 ));
    CascadeMux I__5945 (
            .O(N__35545),
            .I(N__35542));
    InMux I__5944 (
            .O(N__35542),
            .I(N__35539));
    LocalMux I__5943 (
            .O(N__35539),
            .I(\c0.n22474 ));
    InMux I__5942 (
            .O(N__35536),
            .I(N__35533));
    LocalMux I__5941 (
            .O(N__35533),
            .I(\c0.n22483 ));
    CascadeMux I__5940 (
            .O(N__35530),
            .I(N__35526));
    InMux I__5939 (
            .O(N__35529),
            .I(N__35523));
    InMux I__5938 (
            .O(N__35526),
            .I(N__35520));
    LocalMux I__5937 (
            .O(N__35523),
            .I(N__35514));
    LocalMux I__5936 (
            .O(N__35520),
            .I(N__35511));
    InMux I__5935 (
            .O(N__35519),
            .I(N__35508));
    InMux I__5934 (
            .O(N__35518),
            .I(N__35505));
    InMux I__5933 (
            .O(N__35517),
            .I(N__35502));
    Span4Mux_h I__5932 (
            .O(N__35514),
            .I(N__35499));
    Span4Mux_h I__5931 (
            .O(N__35511),
            .I(N__35496));
    LocalMux I__5930 (
            .O(N__35508),
            .I(N__35493));
    LocalMux I__5929 (
            .O(N__35505),
            .I(N__35486));
    LocalMux I__5928 (
            .O(N__35502),
            .I(N__35486));
    Span4Mux_v I__5927 (
            .O(N__35499),
            .I(N__35486));
    Odrv4 I__5926 (
            .O(N__35496),
            .I(encoder1_position_30));
    Odrv12 I__5925 (
            .O(N__35493),
            .I(encoder1_position_30));
    Odrv4 I__5924 (
            .O(N__35486),
            .I(encoder1_position_30));
    CascadeMux I__5923 (
            .O(N__35479),
            .I(\c0.n16_adj_4321_cascade_ ));
    CascadeMux I__5922 (
            .O(N__35476),
            .I(\c0.n18_adj_4322_cascade_ ));
    InMux I__5921 (
            .O(N__35473),
            .I(N__35470));
    LocalMux I__5920 (
            .O(N__35470),
            .I(N__35467));
    Span4Mux_h I__5919 (
            .O(N__35467),
            .I(N__35464));
    Odrv4 I__5918 (
            .O(N__35464),
            .I(\c0.n17_adj_4323 ));
    InMux I__5917 (
            .O(N__35461),
            .I(N__35458));
    LocalMux I__5916 (
            .O(N__35458),
            .I(N__35455));
    Span4Mux_v I__5915 (
            .O(N__35455),
            .I(N__35452));
    Odrv4 I__5914 (
            .O(N__35452),
            .I(\c0.n14_adj_4324 ));
    InMux I__5913 (
            .O(N__35449),
            .I(N__35446));
    LocalMux I__5912 (
            .O(N__35446),
            .I(N__35442));
    InMux I__5911 (
            .O(N__35445),
            .I(N__35439));
    Span12Mux_v I__5910 (
            .O(N__35442),
            .I(N__35434));
    LocalMux I__5909 (
            .O(N__35439),
            .I(N__35434));
    Odrv12 I__5908 (
            .O(N__35434),
            .I(\c0.n22376 ));
    InMux I__5907 (
            .O(N__35431),
            .I(N__35428));
    LocalMux I__5906 (
            .O(N__35428),
            .I(\c0.n13619 ));
    CascadeMux I__5905 (
            .O(N__35425),
            .I(\c0.n13619_cascade_ ));
    InMux I__5904 (
            .O(N__35422),
            .I(N__35419));
    LocalMux I__5903 (
            .O(N__35419),
            .I(N__35415));
    InMux I__5902 (
            .O(N__35418),
            .I(N__35412));
    Span4Mux_h I__5901 (
            .O(N__35415),
            .I(N__35409));
    LocalMux I__5900 (
            .O(N__35412),
            .I(\c0.n22412 ));
    Odrv4 I__5899 (
            .O(N__35409),
            .I(\c0.n22412 ));
    CascadeMux I__5898 (
            .O(N__35404),
            .I(\c0.n13524_cascade_ ));
    InMux I__5897 (
            .O(N__35401),
            .I(N__35398));
    LocalMux I__5896 (
            .O(N__35398),
            .I(\c0.n10_adj_4317 ));
    CascadeMux I__5895 (
            .O(N__35395),
            .I(N__35392));
    InMux I__5894 (
            .O(N__35392),
            .I(N__35387));
    InMux I__5893 (
            .O(N__35391),
            .I(N__35382));
    InMux I__5892 (
            .O(N__35390),
            .I(N__35378));
    LocalMux I__5891 (
            .O(N__35387),
            .I(N__35375));
    InMux I__5890 (
            .O(N__35386),
            .I(N__35370));
    InMux I__5889 (
            .O(N__35385),
            .I(N__35370));
    LocalMux I__5888 (
            .O(N__35382),
            .I(N__35366));
    InMux I__5887 (
            .O(N__35381),
            .I(N__35363));
    LocalMux I__5886 (
            .O(N__35378),
            .I(N__35360));
    Span4Mux_h I__5885 (
            .O(N__35375),
            .I(N__35355));
    LocalMux I__5884 (
            .O(N__35370),
            .I(N__35355));
    InMux I__5883 (
            .O(N__35369),
            .I(N__35352));
    Odrv4 I__5882 (
            .O(N__35366),
            .I(encoder1_position_8));
    LocalMux I__5881 (
            .O(N__35363),
            .I(encoder1_position_8));
    Odrv4 I__5880 (
            .O(N__35360),
            .I(encoder1_position_8));
    Odrv4 I__5879 (
            .O(N__35355),
            .I(encoder1_position_8));
    LocalMux I__5878 (
            .O(N__35352),
            .I(encoder1_position_8));
    InMux I__5877 (
            .O(N__35341),
            .I(N__35338));
    LocalMux I__5876 (
            .O(N__35338),
            .I(N__35335));
    Span4Mux_h I__5875 (
            .O(N__35335),
            .I(N__35331));
    InMux I__5874 (
            .O(N__35334),
            .I(N__35328));
    Span4Mux_h I__5873 (
            .O(N__35331),
            .I(N__35325));
    LocalMux I__5872 (
            .O(N__35328),
            .I(data_out_frame_12_0));
    Odrv4 I__5871 (
            .O(N__35325),
            .I(data_out_frame_12_0));
    CascadeMux I__5870 (
            .O(N__35320),
            .I(N__35317));
    InMux I__5869 (
            .O(N__35317),
            .I(N__35311));
    InMux I__5868 (
            .O(N__35316),
            .I(N__35311));
    LocalMux I__5867 (
            .O(N__35311),
            .I(N__35305));
    InMux I__5866 (
            .O(N__35310),
            .I(N__35300));
    InMux I__5865 (
            .O(N__35309),
            .I(N__35300));
    InMux I__5864 (
            .O(N__35308),
            .I(N__35297));
    Span4Mux_v I__5863 (
            .O(N__35305),
            .I(N__35294));
    LocalMux I__5862 (
            .O(N__35300),
            .I(N__35289));
    LocalMux I__5861 (
            .O(N__35297),
            .I(N__35289));
    Odrv4 I__5860 (
            .O(N__35294),
            .I(\c0.n13079 ));
    Odrv12 I__5859 (
            .O(N__35289),
            .I(\c0.n13079 ));
    InMux I__5858 (
            .O(N__35284),
            .I(N__35280));
    CascadeMux I__5857 (
            .O(N__35283),
            .I(N__35277));
    LocalMux I__5856 (
            .O(N__35280),
            .I(N__35274));
    InMux I__5855 (
            .O(N__35277),
            .I(N__35271));
    Span4Mux_v I__5854 (
            .O(N__35274),
            .I(N__35268));
    LocalMux I__5853 (
            .O(N__35271),
            .I(N__35265));
    Odrv4 I__5852 (
            .O(N__35268),
            .I(\c0.n22174 ));
    Odrv12 I__5851 (
            .O(N__35265),
            .I(\c0.n22174 ));
    CascadeMux I__5850 (
            .O(N__35260),
            .I(N__35257));
    InMux I__5849 (
            .O(N__35257),
            .I(N__35254));
    LocalMux I__5848 (
            .O(N__35254),
            .I(N__35249));
    InMux I__5847 (
            .O(N__35253),
            .I(N__35246));
    InMux I__5846 (
            .O(N__35252),
            .I(N__35242));
    Span4Mux_h I__5845 (
            .O(N__35249),
            .I(N__35239));
    LocalMux I__5844 (
            .O(N__35246),
            .I(N__35236));
    InMux I__5843 (
            .O(N__35245),
            .I(N__35233));
    LocalMux I__5842 (
            .O(N__35242),
            .I(N__35226));
    Sp12to4 I__5841 (
            .O(N__35239),
            .I(N__35226));
    Span12Mux_h I__5840 (
            .O(N__35236),
            .I(N__35226));
    LocalMux I__5839 (
            .O(N__35233),
            .I(data_in_3_5));
    Odrv12 I__5838 (
            .O(N__35226),
            .I(data_in_3_5));
    InMux I__5837 (
            .O(N__35221),
            .I(N__35217));
    InMux I__5836 (
            .O(N__35220),
            .I(N__35214));
    LocalMux I__5835 (
            .O(N__35217),
            .I(N__35210));
    LocalMux I__5834 (
            .O(N__35214),
            .I(N__35205));
    InMux I__5833 (
            .O(N__35213),
            .I(N__35202));
    Span12Mux_h I__5832 (
            .O(N__35210),
            .I(N__35197));
    InMux I__5831 (
            .O(N__35209),
            .I(N__35194));
    InMux I__5830 (
            .O(N__35208),
            .I(N__35191));
    Span4Mux_h I__5829 (
            .O(N__35205),
            .I(N__35186));
    LocalMux I__5828 (
            .O(N__35202),
            .I(N__35186));
    InMux I__5827 (
            .O(N__35201),
            .I(N__35181));
    InMux I__5826 (
            .O(N__35200),
            .I(N__35181));
    Odrv12 I__5825 (
            .O(N__35197),
            .I(encoder1_position_10));
    LocalMux I__5824 (
            .O(N__35194),
            .I(encoder1_position_10));
    LocalMux I__5823 (
            .O(N__35191),
            .I(encoder1_position_10));
    Odrv4 I__5822 (
            .O(N__35186),
            .I(encoder1_position_10));
    LocalMux I__5821 (
            .O(N__35181),
            .I(encoder1_position_10));
    InMux I__5820 (
            .O(N__35170),
            .I(N__35166));
    CascadeMux I__5819 (
            .O(N__35169),
            .I(N__35163));
    LocalMux I__5818 (
            .O(N__35166),
            .I(N__35160));
    InMux I__5817 (
            .O(N__35163),
            .I(N__35157));
    Span4Mux_v I__5816 (
            .O(N__35160),
            .I(N__35154));
    LocalMux I__5815 (
            .O(N__35157),
            .I(data_out_frame_12_2));
    Odrv4 I__5814 (
            .O(N__35154),
            .I(data_out_frame_12_2));
    InMux I__5813 (
            .O(N__35149),
            .I(N__35146));
    LocalMux I__5812 (
            .O(N__35146),
            .I(N__35143));
    Odrv12 I__5811 (
            .O(N__35143),
            .I(\c0.n21918 ));
    CascadeMux I__5810 (
            .O(N__35140),
            .I(N__35136));
    InMux I__5809 (
            .O(N__35139),
            .I(N__35131));
    InMux I__5808 (
            .O(N__35136),
            .I(N__35128));
    InMux I__5807 (
            .O(N__35135),
            .I(N__35123));
    InMux I__5806 (
            .O(N__35134),
            .I(N__35123));
    LocalMux I__5805 (
            .O(N__35131),
            .I(N__35117));
    LocalMux I__5804 (
            .O(N__35128),
            .I(N__35111));
    LocalMux I__5803 (
            .O(N__35123),
            .I(N__35111));
    InMux I__5802 (
            .O(N__35122),
            .I(N__35108));
    InMux I__5801 (
            .O(N__35121),
            .I(N__35103));
    InMux I__5800 (
            .O(N__35120),
            .I(N__35103));
    Span4Mux_v I__5799 (
            .O(N__35117),
            .I(N__35100));
    InMux I__5798 (
            .O(N__35116),
            .I(N__35097));
    Span4Mux_h I__5797 (
            .O(N__35111),
            .I(N__35094));
    LocalMux I__5796 (
            .O(N__35108),
            .I(N__35091));
    LocalMux I__5795 (
            .O(N__35103),
            .I(encoder1_position_4));
    Odrv4 I__5794 (
            .O(N__35100),
            .I(encoder1_position_4));
    LocalMux I__5793 (
            .O(N__35097),
            .I(encoder1_position_4));
    Odrv4 I__5792 (
            .O(N__35094),
            .I(encoder1_position_4));
    Odrv4 I__5791 (
            .O(N__35091),
            .I(encoder1_position_4));
    InMux I__5790 (
            .O(N__35080),
            .I(N__35076));
    InMux I__5789 (
            .O(N__35079),
            .I(N__35073));
    LocalMux I__5788 (
            .O(N__35076),
            .I(N__35070));
    LocalMux I__5787 (
            .O(N__35073),
            .I(data_out_frame_13_4));
    Odrv4 I__5786 (
            .O(N__35070),
            .I(data_out_frame_13_4));
    CascadeMux I__5785 (
            .O(N__35065),
            .I(N__35061));
    CascadeMux I__5784 (
            .O(N__35064),
            .I(N__35058));
    InMux I__5783 (
            .O(N__35061),
            .I(N__35054));
    InMux I__5782 (
            .O(N__35058),
            .I(N__35051));
    InMux I__5781 (
            .O(N__35057),
            .I(N__35048));
    LocalMux I__5780 (
            .O(N__35054),
            .I(N__35043));
    LocalMux I__5779 (
            .O(N__35051),
            .I(N__35043));
    LocalMux I__5778 (
            .O(N__35048),
            .I(N__35039));
    Span4Mux_h I__5777 (
            .O(N__35043),
            .I(N__35036));
    CascadeMux I__5776 (
            .O(N__35042),
            .I(N__35032));
    Span4Mux_h I__5775 (
            .O(N__35039),
            .I(N__35027));
    Span4Mux_h I__5774 (
            .O(N__35036),
            .I(N__35024));
    InMux I__5773 (
            .O(N__35035),
            .I(N__35021));
    InMux I__5772 (
            .O(N__35032),
            .I(N__35016));
    InMux I__5771 (
            .O(N__35031),
            .I(N__35016));
    InMux I__5770 (
            .O(N__35030),
            .I(N__35013));
    Odrv4 I__5769 (
            .O(N__35027),
            .I(encoder1_position_2));
    Odrv4 I__5768 (
            .O(N__35024),
            .I(encoder1_position_2));
    LocalMux I__5767 (
            .O(N__35021),
            .I(encoder1_position_2));
    LocalMux I__5766 (
            .O(N__35016),
            .I(encoder1_position_2));
    LocalMux I__5765 (
            .O(N__35013),
            .I(encoder1_position_2));
    InMux I__5764 (
            .O(N__35002),
            .I(N__34999));
    LocalMux I__5763 (
            .O(N__34999),
            .I(N__34995));
    InMux I__5762 (
            .O(N__34998),
            .I(N__34992));
    Span4Mux_h I__5761 (
            .O(N__34995),
            .I(N__34989));
    LocalMux I__5760 (
            .O(N__34992),
            .I(data_out_frame_13_2));
    Odrv4 I__5759 (
            .O(N__34989),
            .I(data_out_frame_13_2));
    CascadeMux I__5758 (
            .O(N__34984),
            .I(N__34981));
    InMux I__5757 (
            .O(N__34981),
            .I(N__34975));
    InMux I__5756 (
            .O(N__34980),
            .I(N__34972));
    InMux I__5755 (
            .O(N__34979),
            .I(N__34967));
    InMux I__5754 (
            .O(N__34978),
            .I(N__34967));
    LocalMux I__5753 (
            .O(N__34975),
            .I(N__34963));
    LocalMux I__5752 (
            .O(N__34972),
            .I(N__34958));
    LocalMux I__5751 (
            .O(N__34967),
            .I(N__34958));
    CascadeMux I__5750 (
            .O(N__34966),
            .I(N__34954));
    Span4Mux_v I__5749 (
            .O(N__34963),
            .I(N__34949));
    Span4Mux_h I__5748 (
            .O(N__34958),
            .I(N__34949));
    InMux I__5747 (
            .O(N__34957),
            .I(N__34946));
    InMux I__5746 (
            .O(N__34954),
            .I(N__34943));
    Span4Mux_h I__5745 (
            .O(N__34949),
            .I(N__34940));
    LocalMux I__5744 (
            .O(N__34946),
            .I(encoder1_position_6));
    LocalMux I__5743 (
            .O(N__34943),
            .I(encoder1_position_6));
    Odrv4 I__5742 (
            .O(N__34940),
            .I(encoder1_position_6));
    CascadeMux I__5741 (
            .O(N__34933),
            .I(N__34930));
    InMux I__5740 (
            .O(N__34930),
            .I(N__34922));
    CascadeMux I__5739 (
            .O(N__34929),
            .I(N__34919));
    InMux I__5738 (
            .O(N__34928),
            .I(N__34916));
    InMux I__5737 (
            .O(N__34927),
            .I(N__34913));
    InMux I__5736 (
            .O(N__34926),
            .I(N__34908));
    InMux I__5735 (
            .O(N__34925),
            .I(N__34908));
    LocalMux I__5734 (
            .O(N__34922),
            .I(N__34904));
    InMux I__5733 (
            .O(N__34919),
            .I(N__34901));
    LocalMux I__5732 (
            .O(N__34916),
            .I(N__34898));
    LocalMux I__5731 (
            .O(N__34913),
            .I(N__34893));
    LocalMux I__5730 (
            .O(N__34908),
            .I(N__34893));
    InMux I__5729 (
            .O(N__34907),
            .I(N__34890));
    Span4Mux_h I__5728 (
            .O(N__34904),
            .I(N__34887));
    LocalMux I__5727 (
            .O(N__34901),
            .I(N__34884));
    Span4Mux_v I__5726 (
            .O(N__34898),
            .I(N__34879));
    Span4Mux_h I__5725 (
            .O(N__34893),
            .I(N__34879));
    LocalMux I__5724 (
            .O(N__34890),
            .I(encoder1_position_7));
    Odrv4 I__5723 (
            .O(N__34887),
            .I(encoder1_position_7));
    Odrv12 I__5722 (
            .O(N__34884),
            .I(encoder1_position_7));
    Odrv4 I__5721 (
            .O(N__34879),
            .I(encoder1_position_7));
    InMux I__5720 (
            .O(N__34870),
            .I(N__34867));
    LocalMux I__5719 (
            .O(N__34867),
            .I(N__34864));
    Odrv4 I__5718 (
            .O(N__34864),
            .I(\c0.n21896 ));
    InMux I__5717 (
            .O(N__34861),
            .I(N__34858));
    LocalMux I__5716 (
            .O(N__34858),
            .I(N__34854));
    InMux I__5715 (
            .O(N__34857),
            .I(N__34851));
    Span4Mux_v I__5714 (
            .O(N__34854),
            .I(N__34845));
    LocalMux I__5713 (
            .O(N__34851),
            .I(N__34845));
    InMux I__5712 (
            .O(N__34850),
            .I(N__34842));
    Span4Mux_h I__5711 (
            .O(N__34845),
            .I(N__34839));
    LocalMux I__5710 (
            .O(N__34842),
            .I(\c0.n21998 ));
    Odrv4 I__5709 (
            .O(N__34839),
            .I(\c0.n21998 ));
    InMux I__5708 (
            .O(N__34834),
            .I(N__34831));
    LocalMux I__5707 (
            .O(N__34831),
            .I(\c0.n21852 ));
    InMux I__5706 (
            .O(N__34828),
            .I(N__34824));
    CascadeMux I__5705 (
            .O(N__34827),
            .I(N__34821));
    LocalMux I__5704 (
            .O(N__34824),
            .I(N__34818));
    InMux I__5703 (
            .O(N__34821),
            .I(N__34814));
    Span4Mux_h I__5702 (
            .O(N__34818),
            .I(N__34811));
    InMux I__5701 (
            .O(N__34817),
            .I(N__34808));
    LocalMux I__5700 (
            .O(N__34814),
            .I(\c0.n20249 ));
    Odrv4 I__5699 (
            .O(N__34811),
            .I(\c0.n20249 ));
    LocalMux I__5698 (
            .O(N__34808),
            .I(\c0.n20249 ));
    InMux I__5697 (
            .O(N__34801),
            .I(N__34798));
    LocalMux I__5696 (
            .O(N__34798),
            .I(N__34795));
    Span4Mux_v I__5695 (
            .O(N__34795),
            .I(N__34789));
    InMux I__5694 (
            .O(N__34794),
            .I(N__34784));
    InMux I__5693 (
            .O(N__34793),
            .I(N__34784));
    InMux I__5692 (
            .O(N__34792),
            .I(N__34781));
    Odrv4 I__5691 (
            .O(N__34789),
            .I(\c0.n21210 ));
    LocalMux I__5690 (
            .O(N__34784),
            .I(\c0.n21210 ));
    LocalMux I__5689 (
            .O(N__34781),
            .I(\c0.n21210 ));
    InMux I__5688 (
            .O(N__34774),
            .I(N__34771));
    LocalMux I__5687 (
            .O(N__34771),
            .I(\c0.n17_adj_4499 ));
    InMux I__5686 (
            .O(N__34768),
            .I(N__34765));
    LocalMux I__5685 (
            .O(N__34765),
            .I(N__34762));
    Odrv4 I__5684 (
            .O(N__34762),
            .I(\c0.data_out_frame_29_7 ));
    InMux I__5683 (
            .O(N__34759),
            .I(N__34756));
    LocalMux I__5682 (
            .O(N__34756),
            .I(\c0.data_out_frame_28_7 ));
    InMux I__5681 (
            .O(N__34753),
            .I(N__34750));
    LocalMux I__5680 (
            .O(N__34750),
            .I(N__34747));
    Span4Mux_h I__5679 (
            .O(N__34747),
            .I(N__34744));
    Span4Mux_h I__5678 (
            .O(N__34744),
            .I(N__34741));
    Span4Mux_v I__5677 (
            .O(N__34741),
            .I(N__34738));
    Odrv4 I__5676 (
            .O(N__34738),
            .I(\c0.n26_adj_4359 ));
    InMux I__5675 (
            .O(N__34735),
            .I(N__34732));
    LocalMux I__5674 (
            .O(N__34732),
            .I(N__34728));
    InMux I__5673 (
            .O(N__34731),
            .I(N__34725));
    Span4Mux_h I__5672 (
            .O(N__34728),
            .I(N__34722));
    LocalMux I__5671 (
            .O(N__34725),
            .I(data_out_frame_13_1));
    Odrv4 I__5670 (
            .O(N__34722),
            .I(data_out_frame_13_1));
    InMux I__5669 (
            .O(N__34717),
            .I(N__34714));
    LocalMux I__5668 (
            .O(N__34714),
            .I(N__34711));
    Span4Mux_h I__5667 (
            .O(N__34711),
            .I(N__34707));
    InMux I__5666 (
            .O(N__34710),
            .I(N__34704));
    Span4Mux_h I__5665 (
            .O(N__34707),
            .I(N__34701));
    LocalMux I__5664 (
            .O(N__34704),
            .I(data_out_frame_12_1));
    Odrv4 I__5663 (
            .O(N__34701),
            .I(data_out_frame_12_1));
    CascadeMux I__5662 (
            .O(N__34696),
            .I(N__34693));
    InMux I__5661 (
            .O(N__34693),
            .I(N__34690));
    LocalMux I__5660 (
            .O(N__34690),
            .I(N__34687));
    Span4Mux_v I__5659 (
            .O(N__34687),
            .I(N__34684));
    Span4Mux_h I__5658 (
            .O(N__34684),
            .I(N__34681));
    Span4Mux_v I__5657 (
            .O(N__34681),
            .I(N__34678));
    Odrv4 I__5656 (
            .O(N__34678),
            .I(\c0.n11_adj_4520 ));
    InMux I__5655 (
            .O(N__34675),
            .I(N__34672));
    LocalMux I__5654 (
            .O(N__34672),
            .I(N__34669));
    Span4Mux_v I__5653 (
            .O(N__34669),
            .I(N__34665));
    InMux I__5652 (
            .O(N__34668),
            .I(N__34662));
    Span4Mux_h I__5651 (
            .O(N__34665),
            .I(N__34659));
    LocalMux I__5650 (
            .O(N__34662),
            .I(data_out_frame_8_3));
    Odrv4 I__5649 (
            .O(N__34659),
            .I(data_out_frame_8_3));
    CascadeMux I__5648 (
            .O(N__34654),
            .I(N__34651));
    InMux I__5647 (
            .O(N__34651),
            .I(N__34648));
    LocalMux I__5646 (
            .O(N__34648),
            .I(N__34645));
    Span4Mux_v I__5645 (
            .O(N__34645),
            .I(N__34642));
    Span4Mux_h I__5644 (
            .O(N__34642),
            .I(N__34639));
    Odrv4 I__5643 (
            .O(N__34639),
            .I(\c0.n11_adj_4303 ));
    InMux I__5642 (
            .O(N__34636),
            .I(N__34632));
    InMux I__5641 (
            .O(N__34635),
            .I(N__34628));
    LocalMux I__5640 (
            .O(N__34632),
            .I(N__34624));
    InMux I__5639 (
            .O(N__34631),
            .I(N__34618));
    LocalMux I__5638 (
            .O(N__34628),
            .I(N__34615));
    InMux I__5637 (
            .O(N__34627),
            .I(N__34612));
    Span4Mux_h I__5636 (
            .O(N__34624),
            .I(N__34609));
    InMux I__5635 (
            .O(N__34623),
            .I(N__34602));
    InMux I__5634 (
            .O(N__34622),
            .I(N__34602));
    InMux I__5633 (
            .O(N__34621),
            .I(N__34602));
    LocalMux I__5632 (
            .O(N__34618),
            .I(N__34595));
    Span4Mux_v I__5631 (
            .O(N__34615),
            .I(N__34595));
    LocalMux I__5630 (
            .O(N__34612),
            .I(N__34595));
    Odrv4 I__5629 (
            .O(N__34609),
            .I(encoder1_position_12));
    LocalMux I__5628 (
            .O(N__34602),
            .I(encoder1_position_12));
    Odrv4 I__5627 (
            .O(N__34595),
            .I(encoder1_position_12));
    CascadeMux I__5626 (
            .O(N__34588),
            .I(N__34585));
    InMux I__5625 (
            .O(N__34585),
            .I(N__34579));
    InMux I__5624 (
            .O(N__34584),
            .I(N__34579));
    LocalMux I__5623 (
            .O(N__34579),
            .I(data_out_frame_12_4));
    InMux I__5622 (
            .O(N__34576),
            .I(N__34573));
    LocalMux I__5621 (
            .O(N__34573),
            .I(N__34570));
    Odrv4 I__5620 (
            .O(N__34570),
            .I(\c0.n44_adj_4412 ));
    InMux I__5619 (
            .O(N__34567),
            .I(N__34559));
    InMux I__5618 (
            .O(N__34566),
            .I(N__34559));
    InMux I__5617 (
            .O(N__34565),
            .I(N__34556));
    InMux I__5616 (
            .O(N__34564),
            .I(N__34553));
    LocalMux I__5615 (
            .O(N__34559),
            .I(N__34550));
    LocalMux I__5614 (
            .O(N__34556),
            .I(\c0.FRAME_MATCHER_state_14 ));
    LocalMux I__5613 (
            .O(N__34553),
            .I(\c0.FRAME_MATCHER_state_14 ));
    Odrv4 I__5612 (
            .O(N__34550),
            .I(\c0.FRAME_MATCHER_state_14 ));
    CascadeMux I__5611 (
            .O(N__34543),
            .I(N__34537));
    InMux I__5610 (
            .O(N__34542),
            .I(N__34534));
    InMux I__5609 (
            .O(N__34541),
            .I(N__34531));
    InMux I__5608 (
            .O(N__34540),
            .I(N__34526));
    InMux I__5607 (
            .O(N__34537),
            .I(N__34526));
    LocalMux I__5606 (
            .O(N__34534),
            .I(N__34523));
    LocalMux I__5605 (
            .O(N__34531),
            .I(\c0.FRAME_MATCHER_state_21 ));
    LocalMux I__5604 (
            .O(N__34526),
            .I(\c0.FRAME_MATCHER_state_21 ));
    Odrv12 I__5603 (
            .O(N__34523),
            .I(\c0.FRAME_MATCHER_state_21 ));
    SRMux I__5602 (
            .O(N__34516),
            .I(N__34513));
    LocalMux I__5601 (
            .O(N__34513),
            .I(N__34510));
    Span4Mux_h I__5600 (
            .O(N__34510),
            .I(N__34507));
    Odrv4 I__5599 (
            .O(N__34507),
            .I(\c0.n21368 ));
    InMux I__5598 (
            .O(N__34504),
            .I(N__34497));
    InMux I__5597 (
            .O(N__34503),
            .I(N__34497));
    InMux I__5596 (
            .O(N__34502),
            .I(N__34494));
    LocalMux I__5595 (
            .O(N__34497),
            .I(N__34491));
    LocalMux I__5594 (
            .O(N__34494),
            .I(\c0.FRAME_MATCHER_state_29 ));
    Odrv12 I__5593 (
            .O(N__34491),
            .I(\c0.FRAME_MATCHER_state_29 ));
    SRMux I__5592 (
            .O(N__34486),
            .I(N__34483));
    LocalMux I__5591 (
            .O(N__34483),
            .I(N__34480));
    Odrv12 I__5590 (
            .O(N__34480),
            .I(\c0.n21326 ));
    InMux I__5589 (
            .O(N__34477),
            .I(N__34473));
    InMux I__5588 (
            .O(N__34476),
            .I(N__34470));
    LocalMux I__5587 (
            .O(N__34473),
            .I(N__34467));
    LocalMux I__5586 (
            .O(N__34470),
            .I(N__34464));
    Span4Mux_v I__5585 (
            .O(N__34467),
            .I(N__34459));
    Span4Mux_v I__5584 (
            .O(N__34464),
            .I(N__34459));
    Odrv4 I__5583 (
            .O(N__34459),
            .I(\c0.n20658 ));
    InMux I__5582 (
            .O(N__34456),
            .I(N__34449));
    InMux I__5581 (
            .O(N__34455),
            .I(N__34446));
    InMux I__5580 (
            .O(N__34454),
            .I(N__34438));
    InMux I__5579 (
            .O(N__34453),
            .I(N__34438));
    InMux I__5578 (
            .O(N__34452),
            .I(N__34438));
    LocalMux I__5577 (
            .O(N__34449),
            .I(N__34433));
    LocalMux I__5576 (
            .O(N__34446),
            .I(N__34433));
    InMux I__5575 (
            .O(N__34445),
            .I(N__34430));
    LocalMux I__5574 (
            .O(N__34438),
            .I(N__34427));
    Span4Mux_v I__5573 (
            .O(N__34433),
            .I(N__34421));
    LocalMux I__5572 (
            .O(N__34430),
            .I(N__34421));
    Span4Mux_h I__5571 (
            .O(N__34427),
            .I(N__34418));
    InMux I__5570 (
            .O(N__34426),
            .I(N__34415));
    Span4Mux_h I__5569 (
            .O(N__34421),
            .I(N__34412));
    Span4Mux_v I__5568 (
            .O(N__34418),
            .I(N__34409));
    LocalMux I__5567 (
            .O(N__34415),
            .I(N__34406));
    Odrv4 I__5566 (
            .O(N__34412),
            .I(\c0.n21152 ));
    Odrv4 I__5565 (
            .O(N__34409),
            .I(\c0.n21152 ));
    Odrv12 I__5564 (
            .O(N__34406),
            .I(\c0.n21152 ));
    InMux I__5563 (
            .O(N__34399),
            .I(N__34395));
    CascadeMux I__5562 (
            .O(N__34398),
            .I(N__34392));
    LocalMux I__5561 (
            .O(N__34395),
            .I(N__34389));
    InMux I__5560 (
            .O(N__34392),
            .I(N__34383));
    Span4Mux_h I__5559 (
            .O(N__34389),
            .I(N__34380));
    InMux I__5558 (
            .O(N__34388),
            .I(N__34373));
    InMux I__5557 (
            .O(N__34387),
            .I(N__34373));
    InMux I__5556 (
            .O(N__34386),
            .I(N__34373));
    LocalMux I__5555 (
            .O(N__34383),
            .I(\c0.n21168 ));
    Odrv4 I__5554 (
            .O(N__34380),
            .I(\c0.n21168 ));
    LocalMux I__5553 (
            .O(N__34373),
            .I(\c0.n21168 ));
    InMux I__5552 (
            .O(N__34366),
            .I(N__34363));
    LocalMux I__5551 (
            .O(N__34363),
            .I(N__34359));
    InMux I__5550 (
            .O(N__34362),
            .I(N__34356));
    Span4Mux_h I__5549 (
            .O(N__34359),
            .I(N__34353));
    LocalMux I__5548 (
            .O(N__34356),
            .I(\c0.n12542 ));
    Odrv4 I__5547 (
            .O(N__34353),
            .I(\c0.n12542 ));
    InMux I__5546 (
            .O(N__34348),
            .I(N__34345));
    LocalMux I__5545 (
            .O(N__34345),
            .I(N__34340));
    InMux I__5544 (
            .O(N__34344),
            .I(N__34337));
    InMux I__5543 (
            .O(N__34343),
            .I(N__34334));
    Span4Mux_v I__5542 (
            .O(N__34340),
            .I(N__34329));
    LocalMux I__5541 (
            .O(N__34337),
            .I(N__34329));
    LocalMux I__5540 (
            .O(N__34334),
            .I(N__34326));
    Span4Mux_h I__5539 (
            .O(N__34329),
            .I(N__34323));
    Odrv4 I__5538 (
            .O(N__34326),
            .I(\c0.n20180 ));
    Odrv4 I__5537 (
            .O(N__34323),
            .I(\c0.n20180 ));
    InMux I__5536 (
            .O(N__34318),
            .I(N__34315));
    LocalMux I__5535 (
            .O(N__34315),
            .I(\c0.n23260 ));
    CascadeMux I__5534 (
            .O(N__34312),
            .I(\c0.n16_adj_4498_cascade_ ));
    InMux I__5533 (
            .O(N__34309),
            .I(N__34303));
    InMux I__5532 (
            .O(N__34308),
            .I(N__34303));
    LocalMux I__5531 (
            .O(N__34303),
            .I(N__34298));
    InMux I__5530 (
            .O(N__34302),
            .I(N__34295));
    InMux I__5529 (
            .O(N__34301),
            .I(N__34292));
    Span4Mux_h I__5528 (
            .O(N__34298),
            .I(N__34289));
    LocalMux I__5527 (
            .O(N__34295),
            .I(\c0.FRAME_MATCHER_state_22 ));
    LocalMux I__5526 (
            .O(N__34292),
            .I(\c0.FRAME_MATCHER_state_22 ));
    Odrv4 I__5525 (
            .O(N__34289),
            .I(\c0.FRAME_MATCHER_state_22 ));
    CascadeMux I__5524 (
            .O(N__34282),
            .I(\c0.n14457_cascade_ ));
    InMux I__5523 (
            .O(N__34279),
            .I(N__34274));
    InMux I__5522 (
            .O(N__34278),
            .I(N__34269));
    InMux I__5521 (
            .O(N__34277),
            .I(N__34269));
    LocalMux I__5520 (
            .O(N__34274),
            .I(\c0.FRAME_MATCHER_state_27 ));
    LocalMux I__5519 (
            .O(N__34269),
            .I(\c0.FRAME_MATCHER_state_27 ));
    SRMux I__5518 (
            .O(N__34264),
            .I(N__34261));
    LocalMux I__5517 (
            .O(N__34261),
            .I(N__34258));
    Span4Mux_h I__5516 (
            .O(N__34258),
            .I(N__34255));
    Odrv4 I__5515 (
            .O(N__34255),
            .I(\c0.n21330 ));
    CascadeMux I__5514 (
            .O(N__34252),
            .I(\c0.n30_adj_4411_cascade_ ));
    InMux I__5513 (
            .O(N__34249),
            .I(N__34241));
    InMux I__5512 (
            .O(N__34248),
            .I(N__34241));
    InMux I__5511 (
            .O(N__34247),
            .I(N__34238));
    InMux I__5510 (
            .O(N__34246),
            .I(N__34235));
    LocalMux I__5509 (
            .O(N__34241),
            .I(N__34232));
    LocalMux I__5508 (
            .O(N__34238),
            .I(N__34229));
    LocalMux I__5507 (
            .O(N__34235),
            .I(\c0.FRAME_MATCHER_state_8 ));
    Odrv4 I__5506 (
            .O(N__34232),
            .I(\c0.FRAME_MATCHER_state_8 ));
    Odrv4 I__5505 (
            .O(N__34229),
            .I(\c0.FRAME_MATCHER_state_8 ));
    SRMux I__5504 (
            .O(N__34222),
            .I(N__34219));
    LocalMux I__5503 (
            .O(N__34219),
            .I(N__34216));
    Span4Mux_h I__5502 (
            .O(N__34216),
            .I(N__34213));
    Odrv4 I__5501 (
            .O(N__34213),
            .I(\c0.n21344 ));
    SRMux I__5500 (
            .O(N__34210),
            .I(N__34207));
    LocalMux I__5499 (
            .O(N__34207),
            .I(N__34204));
    Span4Mux_h I__5498 (
            .O(N__34204),
            .I(N__34201));
    Odrv4 I__5497 (
            .O(N__34201),
            .I(\c0.n21336 ));
    InMux I__5496 (
            .O(N__34198),
            .I(N__34194));
    InMux I__5495 (
            .O(N__34197),
            .I(N__34189));
    LocalMux I__5494 (
            .O(N__34194),
            .I(N__34186));
    InMux I__5493 (
            .O(N__34193),
            .I(N__34183));
    InMux I__5492 (
            .O(N__34192),
            .I(N__34180));
    LocalMux I__5491 (
            .O(N__34189),
            .I(N__34177));
    Span4Mux_h I__5490 (
            .O(N__34186),
            .I(N__34172));
    LocalMux I__5489 (
            .O(N__34183),
            .I(N__34172));
    LocalMux I__5488 (
            .O(N__34180),
            .I(data_in_2_3));
    Odrv4 I__5487 (
            .O(N__34177),
            .I(data_in_2_3));
    Odrv4 I__5486 (
            .O(N__34172),
            .I(data_in_2_3));
    InMux I__5485 (
            .O(N__34165),
            .I(N__34161));
    InMux I__5484 (
            .O(N__34164),
            .I(N__34158));
    LocalMux I__5483 (
            .O(N__34161),
            .I(N__34153));
    LocalMux I__5482 (
            .O(N__34158),
            .I(N__34150));
    InMux I__5481 (
            .O(N__34157),
            .I(N__34147));
    InMux I__5480 (
            .O(N__34156),
            .I(N__34144));
    Span4Mux_v I__5479 (
            .O(N__34153),
            .I(N__34141));
    Odrv4 I__5478 (
            .O(N__34150),
            .I(data_in_2_1));
    LocalMux I__5477 (
            .O(N__34147),
            .I(data_in_2_1));
    LocalMux I__5476 (
            .O(N__34144),
            .I(data_in_2_1));
    Odrv4 I__5475 (
            .O(N__34141),
            .I(data_in_2_1));
    CascadeMux I__5474 (
            .O(N__34132),
            .I(\c0.n13_adj_4388_cascade_ ));
    InMux I__5473 (
            .O(N__34129),
            .I(N__34126));
    LocalMux I__5472 (
            .O(N__34126),
            .I(\c0.n23135 ));
    InMux I__5471 (
            .O(N__34123),
            .I(N__34120));
    LocalMux I__5470 (
            .O(N__34120),
            .I(N__34116));
    InMux I__5469 (
            .O(N__34119),
            .I(N__34113));
    Span4Mux_h I__5468 (
            .O(N__34116),
            .I(N__34110));
    LocalMux I__5467 (
            .O(N__34113),
            .I(\quad_counter0.b_delay_counter_14 ));
    Odrv4 I__5466 (
            .O(N__34110),
            .I(\quad_counter0.b_delay_counter_14 ));
    InMux I__5465 (
            .O(N__34105),
            .I(N__34102));
    LocalMux I__5464 (
            .O(N__34102),
            .I(N__34098));
    InMux I__5463 (
            .O(N__34101),
            .I(N__34095));
    Span4Mux_h I__5462 (
            .O(N__34098),
            .I(N__34092));
    LocalMux I__5461 (
            .O(N__34095),
            .I(\quad_counter0.b_delay_counter_7 ));
    Odrv4 I__5460 (
            .O(N__34092),
            .I(\quad_counter0.b_delay_counter_7 ));
    CascadeMux I__5459 (
            .O(N__34087),
            .I(N__34084));
    InMux I__5458 (
            .O(N__34084),
            .I(N__34081));
    LocalMux I__5457 (
            .O(N__34081),
            .I(N__34077));
    InMux I__5456 (
            .O(N__34080),
            .I(N__34074));
    Span4Mux_h I__5455 (
            .O(N__34077),
            .I(N__34071));
    LocalMux I__5454 (
            .O(N__34074),
            .I(\quad_counter0.b_delay_counter_12 ));
    Odrv4 I__5453 (
            .O(N__34071),
            .I(\quad_counter0.b_delay_counter_12 ));
    InMux I__5452 (
            .O(N__34066),
            .I(N__34063));
    LocalMux I__5451 (
            .O(N__34063),
            .I(N__34059));
    InMux I__5450 (
            .O(N__34062),
            .I(N__34056));
    Span4Mux_h I__5449 (
            .O(N__34059),
            .I(N__34053));
    LocalMux I__5448 (
            .O(N__34056),
            .I(\quad_counter0.b_delay_counter_15 ));
    Odrv4 I__5447 (
            .O(N__34053),
            .I(\quad_counter0.b_delay_counter_15 ));
    InMux I__5446 (
            .O(N__34048),
            .I(N__34045));
    LocalMux I__5445 (
            .O(N__34045),
            .I(N__34042));
    Span4Mux_h I__5444 (
            .O(N__34042),
            .I(N__34039));
    Odrv4 I__5443 (
            .O(N__34039),
            .I(\quad_counter0.n27_adj_4200 ));
    InMux I__5442 (
            .O(N__34036),
            .I(N__34033));
    LocalMux I__5441 (
            .O(N__34033),
            .I(\c0.n14457 ));
    InMux I__5440 (
            .O(N__34030),
            .I(N__34027));
    LocalMux I__5439 (
            .O(N__34027),
            .I(N__34024));
    Span4Mux_v I__5438 (
            .O(N__34024),
            .I(N__34020));
    InMux I__5437 (
            .O(N__34023),
            .I(N__34017));
    Span4Mux_h I__5436 (
            .O(N__34020),
            .I(N__34014));
    LocalMux I__5435 (
            .O(N__34017),
            .I(data_out_frame_8_0));
    Odrv4 I__5434 (
            .O(N__34014),
            .I(data_out_frame_8_0));
    CascadeMux I__5433 (
            .O(N__34009),
            .I(N__34006));
    InMux I__5432 (
            .O(N__34006),
            .I(N__34000));
    InMux I__5431 (
            .O(N__34005),
            .I(N__34000));
    LocalMux I__5430 (
            .O(N__34000),
            .I(data_out_frame_7_1));
    InMux I__5429 (
            .O(N__33997),
            .I(N__33994));
    LocalMux I__5428 (
            .O(N__33994),
            .I(\c0.n24093 ));
    CascadeMux I__5427 (
            .O(N__33991),
            .I(\c0.n5_adj_4518_cascade_ ));
    InMux I__5426 (
            .O(N__33988),
            .I(N__33985));
    LocalMux I__5425 (
            .O(N__33985),
            .I(N__33982));
    Span4Mux_h I__5424 (
            .O(N__33982),
            .I(N__33979));
    Odrv4 I__5423 (
            .O(N__33979),
            .I(\c0.n23862 ));
    InMux I__5422 (
            .O(N__33976),
            .I(N__33972));
    CascadeMux I__5421 (
            .O(N__33975),
            .I(N__33960));
    LocalMux I__5420 (
            .O(N__33972),
            .I(N__33956));
    InMux I__5419 (
            .O(N__33971),
            .I(N__33949));
    InMux I__5418 (
            .O(N__33970),
            .I(N__33949));
    InMux I__5417 (
            .O(N__33969),
            .I(N__33949));
    InMux I__5416 (
            .O(N__33968),
            .I(N__33939));
    InMux I__5415 (
            .O(N__33967),
            .I(N__33932));
    InMux I__5414 (
            .O(N__33966),
            .I(N__33932));
    InMux I__5413 (
            .O(N__33965),
            .I(N__33927));
    InMux I__5412 (
            .O(N__33964),
            .I(N__33927));
    InMux I__5411 (
            .O(N__33963),
            .I(N__33924));
    InMux I__5410 (
            .O(N__33960),
            .I(N__33919));
    InMux I__5409 (
            .O(N__33959),
            .I(N__33919));
    Span4Mux_v I__5408 (
            .O(N__33956),
            .I(N__33914));
    LocalMux I__5407 (
            .O(N__33949),
            .I(N__33914));
    InMux I__5406 (
            .O(N__33948),
            .I(N__33907));
    InMux I__5405 (
            .O(N__33947),
            .I(N__33907));
    InMux I__5404 (
            .O(N__33946),
            .I(N__33907));
    InMux I__5403 (
            .O(N__33945),
            .I(N__33902));
    InMux I__5402 (
            .O(N__33944),
            .I(N__33902));
    InMux I__5401 (
            .O(N__33943),
            .I(N__33899));
    InMux I__5400 (
            .O(N__33942),
            .I(N__33896));
    LocalMux I__5399 (
            .O(N__33939),
            .I(N__33893));
    InMux I__5398 (
            .O(N__33938),
            .I(N__33890));
    InMux I__5397 (
            .O(N__33937),
            .I(N__33883));
    LocalMux I__5396 (
            .O(N__33932),
            .I(N__33870));
    LocalMux I__5395 (
            .O(N__33927),
            .I(N__33870));
    LocalMux I__5394 (
            .O(N__33924),
            .I(N__33870));
    LocalMux I__5393 (
            .O(N__33919),
            .I(N__33870));
    Span4Mux_v I__5392 (
            .O(N__33914),
            .I(N__33870));
    LocalMux I__5391 (
            .O(N__33907),
            .I(N__33870));
    LocalMux I__5390 (
            .O(N__33902),
            .I(N__33865));
    LocalMux I__5389 (
            .O(N__33899),
            .I(N__33865));
    LocalMux I__5388 (
            .O(N__33896),
            .I(N__33858));
    Span4Mux_h I__5387 (
            .O(N__33893),
            .I(N__33858));
    LocalMux I__5386 (
            .O(N__33890),
            .I(N__33855));
    InMux I__5385 (
            .O(N__33889),
            .I(N__33845));
    InMux I__5384 (
            .O(N__33888),
            .I(N__33845));
    InMux I__5383 (
            .O(N__33887),
            .I(N__33845));
    InMux I__5382 (
            .O(N__33886),
            .I(N__33845));
    LocalMux I__5381 (
            .O(N__33883),
            .I(N__33838));
    Span4Mux_v I__5380 (
            .O(N__33870),
            .I(N__33838));
    Span4Mux_v I__5379 (
            .O(N__33865),
            .I(N__33838));
    InMux I__5378 (
            .O(N__33864),
            .I(N__33835));
    InMux I__5377 (
            .O(N__33863),
            .I(N__33832));
    Span4Mux_h I__5376 (
            .O(N__33858),
            .I(N__33829));
    Span4Mux_h I__5375 (
            .O(N__33855),
            .I(N__33826));
    InMux I__5374 (
            .O(N__33854),
            .I(N__33823));
    LocalMux I__5373 (
            .O(N__33845),
            .I(N__33816));
    Sp12to4 I__5372 (
            .O(N__33838),
            .I(N__33816));
    LocalMux I__5371 (
            .O(N__33835),
            .I(N__33816));
    LocalMux I__5370 (
            .O(N__33832),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__5369 (
            .O(N__33829),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__5368 (
            .O(N__33826),
            .I(\c0.byte_transmit_counter_2 ));
    LocalMux I__5367 (
            .O(N__33823),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv12 I__5366 (
            .O(N__33816),
            .I(\c0.byte_transmit_counter_2 ));
    InMux I__5365 (
            .O(N__33805),
            .I(N__33801));
    InMux I__5364 (
            .O(N__33804),
            .I(N__33798));
    LocalMux I__5363 (
            .O(N__33801),
            .I(N__33795));
    LocalMux I__5362 (
            .O(N__33798),
            .I(data_out_frame_5_7));
    Odrv4 I__5361 (
            .O(N__33795),
            .I(data_out_frame_5_7));
    CascadeMux I__5360 (
            .O(N__33790),
            .I(N__33787));
    InMux I__5359 (
            .O(N__33787),
            .I(N__33784));
    LocalMux I__5358 (
            .O(N__33784),
            .I(N__33781));
    Span4Mux_h I__5357 (
            .O(N__33781),
            .I(N__33778));
    Span4Mux_h I__5356 (
            .O(N__33778),
            .I(N__33775));
    Odrv4 I__5355 (
            .O(N__33775),
            .I(\c0.n24054 ));
    CascadeMux I__5354 (
            .O(N__33772),
            .I(N__33764));
    CascadeMux I__5353 (
            .O(N__33771),
            .I(N__33760));
    InMux I__5352 (
            .O(N__33770),
            .I(N__33757));
    InMux I__5351 (
            .O(N__33769),
            .I(N__33749));
    InMux I__5350 (
            .O(N__33768),
            .I(N__33749));
    InMux I__5349 (
            .O(N__33767),
            .I(N__33749));
    InMux I__5348 (
            .O(N__33764),
            .I(N__33744));
    InMux I__5347 (
            .O(N__33763),
            .I(N__33744));
    InMux I__5346 (
            .O(N__33760),
            .I(N__33741));
    LocalMux I__5345 (
            .O(N__33757),
            .I(N__33738));
    InMux I__5344 (
            .O(N__33756),
            .I(N__33735));
    LocalMux I__5343 (
            .O(N__33749),
            .I(N__33731));
    LocalMux I__5342 (
            .O(N__33744),
            .I(N__33722));
    LocalMux I__5341 (
            .O(N__33741),
            .I(N__33722));
    Span4Mux_v I__5340 (
            .O(N__33738),
            .I(N__33722));
    LocalMux I__5339 (
            .O(N__33735),
            .I(N__33722));
    InMux I__5338 (
            .O(N__33734),
            .I(N__33719));
    Span4Mux_h I__5337 (
            .O(N__33731),
            .I(N__33716));
    Span4Mux_h I__5336 (
            .O(N__33722),
            .I(N__33713));
    LocalMux I__5335 (
            .O(N__33719),
            .I(\c0.tx.r_SM_Main_0 ));
    Odrv4 I__5334 (
            .O(N__33716),
            .I(\c0.tx.r_SM_Main_0 ));
    Odrv4 I__5333 (
            .O(N__33713),
            .I(\c0.tx.r_SM_Main_0 ));
    InMux I__5332 (
            .O(N__33706),
            .I(N__33703));
    LocalMux I__5331 (
            .O(N__33703),
            .I(N__33700));
    Span4Mux_h I__5330 (
            .O(N__33700),
            .I(N__33697));
    Odrv4 I__5329 (
            .O(N__33697),
            .I(\c0.tx.n7086 ));
    CascadeMux I__5328 (
            .O(N__33694),
            .I(N__33673));
    CascadeMux I__5327 (
            .O(N__33693),
            .I(N__33669));
    CascadeMux I__5326 (
            .O(N__33692),
            .I(N__33665));
    CascadeMux I__5325 (
            .O(N__33691),
            .I(N__33660));
    CascadeMux I__5324 (
            .O(N__33690),
            .I(N__33657));
    CascadeMux I__5323 (
            .O(N__33689),
            .I(N__33653));
    CascadeMux I__5322 (
            .O(N__33688),
            .I(N__33649));
    CascadeMux I__5321 (
            .O(N__33687),
            .I(N__33645));
    CascadeMux I__5320 (
            .O(N__33686),
            .I(N__33641));
    CascadeMux I__5319 (
            .O(N__33685),
            .I(N__33637));
    CascadeMux I__5318 (
            .O(N__33684),
            .I(N__33633));
    CascadeMux I__5317 (
            .O(N__33683),
            .I(N__33629));
    CascadeMux I__5316 (
            .O(N__33682),
            .I(N__33625));
    CascadeMux I__5315 (
            .O(N__33681),
            .I(N__33622));
    CascadeMux I__5314 (
            .O(N__33680),
            .I(N__33619));
    CascadeMux I__5313 (
            .O(N__33679),
            .I(N__33616));
    CascadeMux I__5312 (
            .O(N__33678),
            .I(N__33613));
    CascadeMux I__5311 (
            .O(N__33677),
            .I(N__33610));
    CascadeMux I__5310 (
            .O(N__33676),
            .I(N__33607));
    InMux I__5309 (
            .O(N__33673),
            .I(N__33592));
    InMux I__5308 (
            .O(N__33672),
            .I(N__33592));
    InMux I__5307 (
            .O(N__33669),
            .I(N__33592));
    InMux I__5306 (
            .O(N__33668),
            .I(N__33592));
    InMux I__5305 (
            .O(N__33665),
            .I(N__33592));
    InMux I__5304 (
            .O(N__33664),
            .I(N__33592));
    InMux I__5303 (
            .O(N__33663),
            .I(N__33587));
    InMux I__5302 (
            .O(N__33660),
            .I(N__33587));
    InMux I__5301 (
            .O(N__33657),
            .I(N__33570));
    InMux I__5300 (
            .O(N__33656),
            .I(N__33570));
    InMux I__5299 (
            .O(N__33653),
            .I(N__33570));
    InMux I__5298 (
            .O(N__33652),
            .I(N__33570));
    InMux I__5297 (
            .O(N__33649),
            .I(N__33570));
    InMux I__5296 (
            .O(N__33648),
            .I(N__33570));
    InMux I__5295 (
            .O(N__33645),
            .I(N__33570));
    InMux I__5294 (
            .O(N__33644),
            .I(N__33570));
    InMux I__5293 (
            .O(N__33641),
            .I(N__33553));
    InMux I__5292 (
            .O(N__33640),
            .I(N__33553));
    InMux I__5291 (
            .O(N__33637),
            .I(N__33553));
    InMux I__5290 (
            .O(N__33636),
            .I(N__33553));
    InMux I__5289 (
            .O(N__33633),
            .I(N__33553));
    InMux I__5288 (
            .O(N__33632),
            .I(N__33553));
    InMux I__5287 (
            .O(N__33629),
            .I(N__33553));
    InMux I__5286 (
            .O(N__33628),
            .I(N__33553));
    InMux I__5285 (
            .O(N__33625),
            .I(N__33544));
    InMux I__5284 (
            .O(N__33622),
            .I(N__33544));
    InMux I__5283 (
            .O(N__33619),
            .I(N__33544));
    InMux I__5282 (
            .O(N__33616),
            .I(N__33544));
    InMux I__5281 (
            .O(N__33613),
            .I(N__33535));
    InMux I__5280 (
            .O(N__33610),
            .I(N__33535));
    InMux I__5279 (
            .O(N__33607),
            .I(N__33535));
    InMux I__5278 (
            .O(N__33606),
            .I(N__33535));
    InMux I__5277 (
            .O(N__33605),
            .I(N__33532));
    LocalMux I__5276 (
            .O(N__33592),
            .I(N__33527));
    LocalMux I__5275 (
            .O(N__33587),
            .I(N__33527));
    LocalMux I__5274 (
            .O(N__33570),
            .I(N__33522));
    LocalMux I__5273 (
            .O(N__33553),
            .I(N__33522));
    LocalMux I__5272 (
            .O(N__33544),
            .I(N__33517));
    LocalMux I__5271 (
            .O(N__33535),
            .I(N__33517));
    LocalMux I__5270 (
            .O(N__33532),
            .I(N__33514));
    Span4Mux_v I__5269 (
            .O(N__33527),
            .I(N__33509));
    Span4Mux_v I__5268 (
            .O(N__33522),
            .I(N__33509));
    Span4Mux_h I__5267 (
            .O(N__33517),
            .I(N__33506));
    Span4Mux_h I__5266 (
            .O(N__33514),
            .I(N__33499));
    Span4Mux_h I__5265 (
            .O(N__33509),
            .I(N__33499));
    Span4Mux_v I__5264 (
            .O(N__33506),
            .I(N__33499));
    Odrv4 I__5263 (
            .O(N__33499),
            .I(\quad_counter0.n2227 ));
    InMux I__5262 (
            .O(N__33496),
            .I(bfn_14_18_0_));
    CascadeMux I__5261 (
            .O(N__33493),
            .I(\c0.n14474_cascade_ ));
    InMux I__5260 (
            .O(N__33490),
            .I(N__33484));
    InMux I__5259 (
            .O(N__33489),
            .I(N__33484));
    LocalMux I__5258 (
            .O(N__33484),
            .I(data_out_frame_9_1));
    CascadeMux I__5257 (
            .O(N__33481),
            .I(N__33478));
    InMux I__5256 (
            .O(N__33478),
            .I(N__33475));
    LocalMux I__5255 (
            .O(N__33475),
            .I(N__33471));
    InMux I__5254 (
            .O(N__33474),
            .I(N__33468));
    Span4Mux_v I__5253 (
            .O(N__33471),
            .I(N__33465));
    LocalMux I__5252 (
            .O(N__33468),
            .I(data_out_frame_8_1));
    Odrv4 I__5251 (
            .O(N__33465),
            .I(data_out_frame_8_1));
    InMux I__5250 (
            .O(N__33460),
            .I(N__33457));
    LocalMux I__5249 (
            .O(N__33457),
            .I(N__33454));
    Span4Mux_h I__5248 (
            .O(N__33454),
            .I(N__33451));
    Odrv4 I__5247 (
            .O(N__33451),
            .I(\c0.n24186 ));
    InMux I__5246 (
            .O(N__33448),
            .I(N__33445));
    LocalMux I__5245 (
            .O(N__33445),
            .I(n2248));
    InMux I__5244 (
            .O(N__33442),
            .I(N__33439));
    LocalMux I__5243 (
            .O(N__33439),
            .I(n2240));
    InMux I__5242 (
            .O(N__33436),
            .I(N__33433));
    LocalMux I__5241 (
            .O(N__33433),
            .I(N__33429));
    InMux I__5240 (
            .O(N__33432),
            .I(N__33426));
    Span4Mux_h I__5239 (
            .O(N__33429),
            .I(N__33423));
    LocalMux I__5238 (
            .O(N__33426),
            .I(data_out_frame_7_7));
    Odrv4 I__5237 (
            .O(N__33423),
            .I(data_out_frame_7_7));
    CascadeMux I__5236 (
            .O(N__33418),
            .I(N__33415));
    InMux I__5235 (
            .O(N__33415),
            .I(N__33409));
    InMux I__5234 (
            .O(N__33414),
            .I(N__33409));
    LocalMux I__5233 (
            .O(N__33409),
            .I(data_out_frame_5_1));
    InMux I__5232 (
            .O(N__33406),
            .I(bfn_14_17_0_));
    InMux I__5231 (
            .O(N__33403),
            .I(\quad_counter0.n19604 ));
    InMux I__5230 (
            .O(N__33400),
            .I(\quad_counter0.n19605 ));
    InMux I__5229 (
            .O(N__33397),
            .I(\quad_counter0.n19606 ));
    CascadeMux I__5228 (
            .O(N__33394),
            .I(N__33391));
    InMux I__5227 (
            .O(N__33391),
            .I(N__33388));
    LocalMux I__5226 (
            .O(N__33388),
            .I(N__33383));
    CascadeMux I__5225 (
            .O(N__33387),
            .I(N__33380));
    InMux I__5224 (
            .O(N__33386),
            .I(N__33377));
    Span4Mux_h I__5223 (
            .O(N__33383),
            .I(N__33373));
    InMux I__5222 (
            .O(N__33380),
            .I(N__33370));
    LocalMux I__5221 (
            .O(N__33377),
            .I(N__33367));
    CascadeMux I__5220 (
            .O(N__33376),
            .I(N__33363));
    Sp12to4 I__5219 (
            .O(N__33373),
            .I(N__33358));
    LocalMux I__5218 (
            .O(N__33370),
            .I(N__33358));
    Span4Mux_h I__5217 (
            .O(N__33367),
            .I(N__33355));
    InMux I__5216 (
            .O(N__33366),
            .I(N__33350));
    InMux I__5215 (
            .O(N__33363),
            .I(N__33350));
    Odrv12 I__5214 (
            .O(N__33358),
            .I(encoder0_position_27));
    Odrv4 I__5213 (
            .O(N__33355),
            .I(encoder0_position_27));
    LocalMux I__5212 (
            .O(N__33350),
            .I(encoder0_position_27));
    InMux I__5211 (
            .O(N__33343),
            .I(N__33340));
    LocalMux I__5210 (
            .O(N__33340),
            .I(N__33337));
    Odrv12 I__5209 (
            .O(N__33337),
            .I(n2244));
    InMux I__5208 (
            .O(N__33334),
            .I(\quad_counter0.n19607 ));
    InMux I__5207 (
            .O(N__33331),
            .I(\quad_counter0.n19608 ));
    InMux I__5206 (
            .O(N__33328),
            .I(\quad_counter0.n19609 ));
    InMux I__5205 (
            .O(N__33325),
            .I(N__33322));
    LocalMux I__5204 (
            .O(N__33322),
            .I(N__33319));
    Span4Mux_v I__5203 (
            .O(N__33319),
            .I(N__33316));
    Odrv4 I__5202 (
            .O(N__33316),
            .I(n2241));
    InMux I__5201 (
            .O(N__33313),
            .I(\quad_counter0.n19610 ));
    InMux I__5200 (
            .O(N__33310),
            .I(N__33307));
    LocalMux I__5199 (
            .O(N__33307),
            .I(N__33304));
    Odrv4 I__5198 (
            .O(N__33304),
            .I(n2257));
    InMux I__5197 (
            .O(N__33301),
            .I(\quad_counter0.n19594 ));
    InMux I__5196 (
            .O(N__33298),
            .I(bfn_14_16_0_));
    InMux I__5195 (
            .O(N__33295),
            .I(\quad_counter0.n19596 ));
    InMux I__5194 (
            .O(N__33292),
            .I(\quad_counter0.n19597 ));
    InMux I__5193 (
            .O(N__33289),
            .I(\quad_counter0.n19598 ));
    InMux I__5192 (
            .O(N__33286),
            .I(N__33283));
    LocalMux I__5191 (
            .O(N__33283),
            .I(n2252));
    InMux I__5190 (
            .O(N__33280),
            .I(\quad_counter0.n19599 ));
    InMux I__5189 (
            .O(N__33277),
            .I(N__33274));
    LocalMux I__5188 (
            .O(N__33274),
            .I(N__33271));
    Odrv4 I__5187 (
            .O(N__33271),
            .I(n2251));
    InMux I__5186 (
            .O(N__33268),
            .I(\quad_counter0.n19600 ));
    InMux I__5185 (
            .O(N__33265),
            .I(\quad_counter0.n19601 ));
    InMux I__5184 (
            .O(N__33262),
            .I(\quad_counter0.n19602 ));
    InMux I__5183 (
            .O(N__33259),
            .I(\quad_counter0.n19585 ));
    InMux I__5182 (
            .O(N__33256),
            .I(\quad_counter0.n19586 ));
    CascadeMux I__5181 (
            .O(N__33253),
            .I(N__33250));
    InMux I__5180 (
            .O(N__33250),
            .I(N__33246));
    InMux I__5179 (
            .O(N__33249),
            .I(N__33240));
    LocalMux I__5178 (
            .O(N__33246),
            .I(N__33237));
    CascadeMux I__5177 (
            .O(N__33245),
            .I(N__33234));
    InMux I__5176 (
            .O(N__33244),
            .I(N__33231));
    CascadeMux I__5175 (
            .O(N__33243),
            .I(N__33227));
    LocalMux I__5174 (
            .O(N__33240),
            .I(N__33222));
    Span4Mux_v I__5173 (
            .O(N__33237),
            .I(N__33222));
    InMux I__5172 (
            .O(N__33234),
            .I(N__33219));
    LocalMux I__5171 (
            .O(N__33231),
            .I(N__33216));
    InMux I__5170 (
            .O(N__33230),
            .I(N__33213));
    InMux I__5169 (
            .O(N__33227),
            .I(N__33210));
    Odrv4 I__5168 (
            .O(N__33222),
            .I(encoder0_position_7));
    LocalMux I__5167 (
            .O(N__33219),
            .I(encoder0_position_7));
    Odrv4 I__5166 (
            .O(N__33216),
            .I(encoder0_position_7));
    LocalMux I__5165 (
            .O(N__33213),
            .I(encoder0_position_7));
    LocalMux I__5164 (
            .O(N__33210),
            .I(encoder0_position_7));
    InMux I__5163 (
            .O(N__33199),
            .I(N__33196));
    LocalMux I__5162 (
            .O(N__33196),
            .I(n2264));
    InMux I__5161 (
            .O(N__33193),
            .I(bfn_14_15_0_));
    InMux I__5160 (
            .O(N__33190),
            .I(\quad_counter0.n19588 ));
    InMux I__5159 (
            .O(N__33187),
            .I(\quad_counter0.n19589 ));
    InMux I__5158 (
            .O(N__33184),
            .I(\quad_counter0.n19590 ));
    InMux I__5157 (
            .O(N__33181),
            .I(\quad_counter0.n19591 ));
    InMux I__5156 (
            .O(N__33178),
            .I(\quad_counter0.n19592 ));
    InMux I__5155 (
            .O(N__33175),
            .I(N__33172));
    LocalMux I__5154 (
            .O(N__33172),
            .I(N__33169));
    Odrv4 I__5153 (
            .O(N__33169),
            .I(n2258));
    InMux I__5152 (
            .O(N__33166),
            .I(\quad_counter0.n19593 ));
    InMux I__5151 (
            .O(N__33163),
            .I(N__33151));
    InMux I__5150 (
            .O(N__33162),
            .I(N__33151));
    InMux I__5149 (
            .O(N__33161),
            .I(N__33151));
    InMux I__5148 (
            .O(N__33160),
            .I(N__33151));
    LocalMux I__5147 (
            .O(N__33151),
            .I(N__33148));
    Odrv4 I__5146 (
            .O(N__33148),
            .I(\c0.n20160 ));
    CascadeMux I__5145 (
            .O(N__33145),
            .I(N__33142));
    InMux I__5144 (
            .O(N__33142),
            .I(N__33139));
    LocalMux I__5143 (
            .O(N__33139),
            .I(N__33136));
    Span4Mux_v I__5142 (
            .O(N__33136),
            .I(N__33133));
    Span4Mux_v I__5141 (
            .O(N__33133),
            .I(N__33130));
    Span4Mux_h I__5140 (
            .O(N__33130),
            .I(N__33127));
    Odrv4 I__5139 (
            .O(N__33127),
            .I(\quad_counter0.count_direction ));
    InMux I__5138 (
            .O(N__33124),
            .I(\quad_counter0.n19580 ));
    InMux I__5137 (
            .O(N__33121),
            .I(N__33118));
    LocalMux I__5136 (
            .O(N__33118),
            .I(n2270));
    InMux I__5135 (
            .O(N__33115),
            .I(\quad_counter0.n19581 ));
    InMux I__5134 (
            .O(N__33112),
            .I(N__33109));
    LocalMux I__5133 (
            .O(N__33109),
            .I(n2269));
    InMux I__5132 (
            .O(N__33106),
            .I(\quad_counter0.n19582 ));
    InMux I__5131 (
            .O(N__33103),
            .I(N__33100));
    LocalMux I__5130 (
            .O(N__33100),
            .I(N__33097));
    Span4Mux_h I__5129 (
            .O(N__33097),
            .I(N__33094));
    Odrv4 I__5128 (
            .O(N__33094),
            .I(n2268));
    InMux I__5127 (
            .O(N__33091),
            .I(\quad_counter0.n19583 ));
    InMux I__5126 (
            .O(N__33088),
            .I(\quad_counter0.n19584 ));
    InMux I__5125 (
            .O(N__33085),
            .I(N__33081));
    CascadeMux I__5124 (
            .O(N__33084),
            .I(N__33078));
    LocalMux I__5123 (
            .O(N__33081),
            .I(N__33075));
    InMux I__5122 (
            .O(N__33078),
            .I(N__33072));
    Span4Mux_h I__5121 (
            .O(N__33075),
            .I(N__33069));
    LocalMux I__5120 (
            .O(N__33072),
            .I(\c0.n21943 ));
    Odrv4 I__5119 (
            .O(N__33069),
            .I(\c0.n21943 ));
    CascadeMux I__5118 (
            .O(N__33064),
            .I(N__33061));
    InMux I__5117 (
            .O(N__33061),
            .I(N__33051));
    InMux I__5116 (
            .O(N__33060),
            .I(N__33051));
    InMux I__5115 (
            .O(N__33059),
            .I(N__33043));
    InMux I__5114 (
            .O(N__33058),
            .I(N__33043));
    InMux I__5113 (
            .O(N__33057),
            .I(N__33043));
    InMux I__5112 (
            .O(N__33056),
            .I(N__33040));
    LocalMux I__5111 (
            .O(N__33051),
            .I(N__33037));
    InMux I__5110 (
            .O(N__33050),
            .I(N__33034));
    LocalMux I__5109 (
            .O(N__33043),
            .I(N__33031));
    LocalMux I__5108 (
            .O(N__33040),
            .I(\c0.n21196 ));
    Odrv12 I__5107 (
            .O(N__33037),
            .I(\c0.n21196 ));
    LocalMux I__5106 (
            .O(N__33034),
            .I(\c0.n21196 ));
    Odrv4 I__5105 (
            .O(N__33031),
            .I(\c0.n21196 ));
    CascadeMux I__5104 (
            .O(N__33022),
            .I(N__33019));
    InMux I__5103 (
            .O(N__33019),
            .I(N__33014));
    CascadeMux I__5102 (
            .O(N__33018),
            .I(N__33011));
    CascadeMux I__5101 (
            .O(N__33017),
            .I(N__33007));
    LocalMux I__5100 (
            .O(N__33014),
            .I(N__33004));
    InMux I__5099 (
            .O(N__33011),
            .I(N__33001));
    InMux I__5098 (
            .O(N__33010),
            .I(N__32998));
    InMux I__5097 (
            .O(N__33007),
            .I(N__32995));
    Span4Mux_h I__5096 (
            .O(N__33004),
            .I(N__32992));
    LocalMux I__5095 (
            .O(N__33001),
            .I(N__32989));
    LocalMux I__5094 (
            .O(N__32998),
            .I(encoder1_position_25));
    LocalMux I__5093 (
            .O(N__32995),
            .I(encoder1_position_25));
    Odrv4 I__5092 (
            .O(N__32992),
            .I(encoder1_position_25));
    Odrv4 I__5091 (
            .O(N__32989),
            .I(encoder1_position_25));
    CascadeMux I__5090 (
            .O(N__32980),
            .I(N__32976));
    InMux I__5089 (
            .O(N__32979),
            .I(N__32972));
    InMux I__5088 (
            .O(N__32976),
            .I(N__32969));
    CascadeMux I__5087 (
            .O(N__32975),
            .I(N__32966));
    LocalMux I__5086 (
            .O(N__32972),
            .I(N__32962));
    LocalMux I__5085 (
            .O(N__32969),
            .I(N__32959));
    InMux I__5084 (
            .O(N__32966),
            .I(N__32956));
    InMux I__5083 (
            .O(N__32965),
            .I(N__32952));
    Span4Mux_v I__5082 (
            .O(N__32962),
            .I(N__32945));
    Span4Mux_h I__5081 (
            .O(N__32959),
            .I(N__32945));
    LocalMux I__5080 (
            .O(N__32956),
            .I(N__32945));
    InMux I__5079 (
            .O(N__32955),
            .I(N__32942));
    LocalMux I__5078 (
            .O(N__32952),
            .I(encoder1_position_11));
    Odrv4 I__5077 (
            .O(N__32945),
            .I(encoder1_position_11));
    LocalMux I__5076 (
            .O(N__32942),
            .I(encoder1_position_11));
    CascadeMux I__5075 (
            .O(N__32935),
            .I(\c0.n20232_cascade_ ));
    InMux I__5074 (
            .O(N__32932),
            .I(N__32928));
    InMux I__5073 (
            .O(N__32931),
            .I(N__32925));
    LocalMux I__5072 (
            .O(N__32928),
            .I(N__32920));
    LocalMux I__5071 (
            .O(N__32925),
            .I(N__32920));
    Span4Mux_h I__5070 (
            .O(N__32920),
            .I(N__32915));
    InMux I__5069 (
            .O(N__32919),
            .I(N__32910));
    InMux I__5068 (
            .O(N__32918),
            .I(N__32910));
    Odrv4 I__5067 (
            .O(N__32915),
            .I(\c0.n21146 ));
    LocalMux I__5066 (
            .O(N__32910),
            .I(\c0.n21146 ));
    CascadeMux I__5065 (
            .O(N__32905),
            .I(\c0.n21146_cascade_ ));
    InMux I__5064 (
            .O(N__32902),
            .I(N__32897));
    CascadeMux I__5063 (
            .O(N__32901),
            .I(N__32894));
    CascadeMux I__5062 (
            .O(N__32900),
            .I(N__32889));
    LocalMux I__5061 (
            .O(N__32897),
            .I(N__32886));
    InMux I__5060 (
            .O(N__32894),
            .I(N__32883));
    InMux I__5059 (
            .O(N__32893),
            .I(N__32880));
    InMux I__5058 (
            .O(N__32892),
            .I(N__32877));
    InMux I__5057 (
            .O(N__32889),
            .I(N__32874));
    Span4Mux_h I__5056 (
            .O(N__32886),
            .I(N__32871));
    LocalMux I__5055 (
            .O(N__32883),
            .I(N__32868));
    LocalMux I__5054 (
            .O(N__32880),
            .I(encoder1_position_23));
    LocalMux I__5053 (
            .O(N__32877),
            .I(encoder1_position_23));
    LocalMux I__5052 (
            .O(N__32874),
            .I(encoder1_position_23));
    Odrv4 I__5051 (
            .O(N__32871),
            .I(encoder1_position_23));
    Odrv4 I__5050 (
            .O(N__32868),
            .I(encoder1_position_23));
    InMux I__5049 (
            .O(N__32857),
            .I(N__32853));
    InMux I__5048 (
            .O(N__32856),
            .I(N__32849));
    LocalMux I__5047 (
            .O(N__32853),
            .I(N__32846));
    InMux I__5046 (
            .O(N__32852),
            .I(N__32842));
    LocalMux I__5045 (
            .O(N__32849),
            .I(N__32839));
    Span4Mux_h I__5044 (
            .O(N__32846),
            .I(N__32836));
    InMux I__5043 (
            .O(N__32845),
            .I(N__32833));
    LocalMux I__5042 (
            .O(N__32842),
            .I(\c0.n20232 ));
    Odrv4 I__5041 (
            .O(N__32839),
            .I(\c0.n20232 ));
    Odrv4 I__5040 (
            .O(N__32836),
            .I(\c0.n20232 ));
    LocalMux I__5039 (
            .O(N__32833),
            .I(\c0.n20232 ));
    InMux I__5038 (
            .O(N__32824),
            .I(N__32820));
    InMux I__5037 (
            .O(N__32823),
            .I(N__32817));
    LocalMux I__5036 (
            .O(N__32820),
            .I(N__32811));
    LocalMux I__5035 (
            .O(N__32817),
            .I(N__32811));
    InMux I__5034 (
            .O(N__32816),
            .I(N__32808));
    Span4Mux_h I__5033 (
            .O(N__32811),
            .I(N__32805));
    LocalMux I__5032 (
            .O(N__32808),
            .I(\c0.n20744 ));
    Odrv4 I__5031 (
            .O(N__32805),
            .I(\c0.n20744 ));
    CascadeMux I__5030 (
            .O(N__32800),
            .I(N__32796));
    CascadeMux I__5029 (
            .O(N__32799),
            .I(N__32793));
    InMux I__5028 (
            .O(N__32796),
            .I(N__32786));
    InMux I__5027 (
            .O(N__32793),
            .I(N__32781));
    InMux I__5026 (
            .O(N__32792),
            .I(N__32778));
    InMux I__5025 (
            .O(N__32791),
            .I(N__32773));
    InMux I__5024 (
            .O(N__32790),
            .I(N__32773));
    InMux I__5023 (
            .O(N__32789),
            .I(N__32770));
    LocalMux I__5022 (
            .O(N__32786),
            .I(N__32767));
    InMux I__5021 (
            .O(N__32785),
            .I(N__32764));
    InMux I__5020 (
            .O(N__32784),
            .I(N__32761));
    LocalMux I__5019 (
            .O(N__32781),
            .I(N__32758));
    LocalMux I__5018 (
            .O(N__32778),
            .I(N__32753));
    LocalMux I__5017 (
            .O(N__32773),
            .I(N__32753));
    LocalMux I__5016 (
            .O(N__32770),
            .I(encoder1_position_1));
    Odrv12 I__5015 (
            .O(N__32767),
            .I(encoder1_position_1));
    LocalMux I__5014 (
            .O(N__32764),
            .I(encoder1_position_1));
    LocalMux I__5013 (
            .O(N__32761),
            .I(encoder1_position_1));
    Odrv4 I__5012 (
            .O(N__32758),
            .I(encoder1_position_1));
    Odrv12 I__5011 (
            .O(N__32753),
            .I(encoder1_position_1));
    CascadeMux I__5010 (
            .O(N__32740),
            .I(N__32735));
    CascadeMux I__5009 (
            .O(N__32739),
            .I(N__32730));
    CascadeMux I__5008 (
            .O(N__32738),
            .I(N__32727));
    InMux I__5007 (
            .O(N__32735),
            .I(N__32721));
    CascadeMux I__5006 (
            .O(N__32734),
            .I(N__32718));
    InMux I__5005 (
            .O(N__32733),
            .I(N__32715));
    InMux I__5004 (
            .O(N__32730),
            .I(N__32712));
    InMux I__5003 (
            .O(N__32727),
            .I(N__32705));
    InMux I__5002 (
            .O(N__32726),
            .I(N__32705));
    InMux I__5001 (
            .O(N__32725),
            .I(N__32705));
    CascadeMux I__5000 (
            .O(N__32724),
            .I(N__32701));
    LocalMux I__4999 (
            .O(N__32721),
            .I(N__32697));
    InMux I__4998 (
            .O(N__32718),
            .I(N__32694));
    LocalMux I__4997 (
            .O(N__32715),
            .I(N__32691));
    LocalMux I__4996 (
            .O(N__32712),
            .I(N__32688));
    LocalMux I__4995 (
            .O(N__32705),
            .I(N__32685));
    InMux I__4994 (
            .O(N__32704),
            .I(N__32680));
    InMux I__4993 (
            .O(N__32701),
            .I(N__32680));
    InMux I__4992 (
            .O(N__32700),
            .I(N__32677));
    Span4Mux_v I__4991 (
            .O(N__32697),
            .I(N__32670));
    LocalMux I__4990 (
            .O(N__32694),
            .I(N__32670));
    Span4Mux_h I__4989 (
            .O(N__32691),
            .I(N__32670));
    Span4Mux_h I__4988 (
            .O(N__32688),
            .I(N__32667));
    Sp12to4 I__4987 (
            .O(N__32685),
            .I(N__32662));
    LocalMux I__4986 (
            .O(N__32680),
            .I(N__32662));
    LocalMux I__4985 (
            .O(N__32677),
            .I(encoder1_position_5));
    Odrv4 I__4984 (
            .O(N__32670),
            .I(encoder1_position_5));
    Odrv4 I__4983 (
            .O(N__32667),
            .I(encoder1_position_5));
    Odrv12 I__4982 (
            .O(N__32662),
            .I(encoder1_position_5));
    CascadeMux I__4981 (
            .O(N__32653),
            .I(\c0.n22163_cascade_ ));
    InMux I__4980 (
            .O(N__32650),
            .I(N__32647));
    LocalMux I__4979 (
            .O(N__32647),
            .I(\c0.n20_adj_4505 ));
    CascadeMux I__4978 (
            .O(N__32644),
            .I(\c0.n19_adj_4506_cascade_ ));
    InMux I__4977 (
            .O(N__32641),
            .I(N__32638));
    LocalMux I__4976 (
            .O(N__32638),
            .I(N__32634));
    InMux I__4975 (
            .O(N__32637),
            .I(N__32631));
    Odrv4 I__4974 (
            .O(N__32634),
            .I(\c0.n21283 ));
    LocalMux I__4973 (
            .O(N__32631),
            .I(\c0.n21283 ));
    InMux I__4972 (
            .O(N__32626),
            .I(N__32623));
    LocalMux I__4971 (
            .O(N__32623),
            .I(N__32620));
    Odrv4 I__4970 (
            .O(N__32620),
            .I(\c0.n6_adj_4508 ));
    InMux I__4969 (
            .O(N__32617),
            .I(N__32613));
    InMux I__4968 (
            .O(N__32616),
            .I(N__32610));
    LocalMux I__4967 (
            .O(N__32613),
            .I(N__32607));
    LocalMux I__4966 (
            .O(N__32610),
            .I(N__32604));
    Span4Mux_h I__4965 (
            .O(N__32607),
            .I(N__32601));
    Span4Mux_v I__4964 (
            .O(N__32604),
            .I(N__32598));
    Odrv4 I__4963 (
            .O(N__32601),
            .I(\c0.n21116 ));
    Odrv4 I__4962 (
            .O(N__32598),
            .I(\c0.n21116 ));
    InMux I__4961 (
            .O(N__32593),
            .I(N__32589));
    InMux I__4960 (
            .O(N__32592),
            .I(N__32586));
    LocalMux I__4959 (
            .O(N__32589),
            .I(N__32583));
    LocalMux I__4958 (
            .O(N__32586),
            .I(N__32580));
    Span4Mux_h I__4957 (
            .O(N__32583),
            .I(N__32577));
    Odrv12 I__4956 (
            .O(N__32580),
            .I(\c0.n20819 ));
    Odrv4 I__4955 (
            .O(N__32577),
            .I(\c0.n20819 ));
    InMux I__4954 (
            .O(N__32572),
            .I(N__32569));
    LocalMux I__4953 (
            .O(N__32569),
            .I(\c0.n21_adj_4507 ));
    CascadeMux I__4952 (
            .O(N__32566),
            .I(N__32562));
    InMux I__4951 (
            .O(N__32565),
            .I(N__32558));
    InMux I__4950 (
            .O(N__32562),
            .I(N__32555));
    InMux I__4949 (
            .O(N__32561),
            .I(N__32549));
    LocalMux I__4948 (
            .O(N__32558),
            .I(N__32544));
    LocalMux I__4947 (
            .O(N__32555),
            .I(N__32544));
    InMux I__4946 (
            .O(N__32554),
            .I(N__32541));
    InMux I__4945 (
            .O(N__32553),
            .I(N__32538));
    InMux I__4944 (
            .O(N__32552),
            .I(N__32535));
    LocalMux I__4943 (
            .O(N__32549),
            .I(N__32526));
    Span4Mux_h I__4942 (
            .O(N__32544),
            .I(N__32526));
    LocalMux I__4941 (
            .O(N__32541),
            .I(N__32526));
    LocalMux I__4940 (
            .O(N__32538),
            .I(N__32526));
    LocalMux I__4939 (
            .O(N__32535),
            .I(N__32521));
    Span4Mux_v I__4938 (
            .O(N__32526),
            .I(N__32521));
    Odrv4 I__4937 (
            .O(N__32521),
            .I(\c0.n20276 ));
    InMux I__4936 (
            .O(N__32518),
            .I(N__32513));
    InMux I__4935 (
            .O(N__32517),
            .I(N__32509));
    InMux I__4934 (
            .O(N__32516),
            .I(N__32506));
    LocalMux I__4933 (
            .O(N__32513),
            .I(N__32502));
    InMux I__4932 (
            .O(N__32512),
            .I(N__32499));
    LocalMux I__4931 (
            .O(N__32509),
            .I(N__32495));
    LocalMux I__4930 (
            .O(N__32506),
            .I(N__32490));
    InMux I__4929 (
            .O(N__32505),
            .I(N__32487));
    Span4Mux_v I__4928 (
            .O(N__32502),
            .I(N__32482));
    LocalMux I__4927 (
            .O(N__32499),
            .I(N__32482));
    InMux I__4926 (
            .O(N__32498),
            .I(N__32479));
    Span4Mux_h I__4925 (
            .O(N__32495),
            .I(N__32476));
    InMux I__4924 (
            .O(N__32494),
            .I(N__32473));
    InMux I__4923 (
            .O(N__32493),
            .I(N__32470));
    Span4Mux_h I__4922 (
            .O(N__32490),
            .I(N__32465));
    LocalMux I__4921 (
            .O(N__32487),
            .I(N__32465));
    Span4Mux_v I__4920 (
            .O(N__32482),
            .I(N__32460));
    LocalMux I__4919 (
            .O(N__32479),
            .I(N__32460));
    Odrv4 I__4918 (
            .O(N__32476),
            .I(\c0.n21122 ));
    LocalMux I__4917 (
            .O(N__32473),
            .I(\c0.n21122 ));
    LocalMux I__4916 (
            .O(N__32470),
            .I(\c0.n21122 ));
    Odrv4 I__4915 (
            .O(N__32465),
            .I(\c0.n21122 ));
    Odrv4 I__4914 (
            .O(N__32460),
            .I(\c0.n21122 ));
    CascadeMux I__4913 (
            .O(N__32449),
            .I(N__32443));
    CascadeMux I__4912 (
            .O(N__32448),
            .I(N__32439));
    InMux I__4911 (
            .O(N__32447),
            .I(N__32434));
    InMux I__4910 (
            .O(N__32446),
            .I(N__32434));
    InMux I__4909 (
            .O(N__32443),
            .I(N__32431));
    InMux I__4908 (
            .O(N__32442),
            .I(N__32428));
    InMux I__4907 (
            .O(N__32439),
            .I(N__32425));
    LocalMux I__4906 (
            .O(N__32434),
            .I(N__32422));
    LocalMux I__4905 (
            .O(N__32431),
            .I(N__32417));
    LocalMux I__4904 (
            .O(N__32428),
            .I(N__32414));
    LocalMux I__4903 (
            .O(N__32425),
            .I(N__32411));
    Span4Mux_h I__4902 (
            .O(N__32422),
            .I(N__32408));
    InMux I__4901 (
            .O(N__32421),
            .I(N__32403));
    InMux I__4900 (
            .O(N__32420),
            .I(N__32403));
    Span4Mux_v I__4899 (
            .O(N__32417),
            .I(N__32398));
    Span4Mux_h I__4898 (
            .O(N__32414),
            .I(N__32398));
    Odrv4 I__4897 (
            .O(N__32411),
            .I(\c0.n21166 ));
    Odrv4 I__4896 (
            .O(N__32408),
            .I(\c0.n21166 ));
    LocalMux I__4895 (
            .O(N__32403),
            .I(\c0.n21166 ));
    Odrv4 I__4894 (
            .O(N__32398),
            .I(\c0.n21166 ));
    CascadeMux I__4893 (
            .O(N__32389),
            .I(N__32386));
    InMux I__4892 (
            .O(N__32386),
            .I(N__32381));
    CascadeMux I__4891 (
            .O(N__32385),
            .I(N__32377));
    CascadeMux I__4890 (
            .O(N__32384),
            .I(N__32374));
    LocalMux I__4889 (
            .O(N__32381),
            .I(N__32368));
    InMux I__4888 (
            .O(N__32380),
            .I(N__32364));
    InMux I__4887 (
            .O(N__32377),
            .I(N__32361));
    InMux I__4886 (
            .O(N__32374),
            .I(N__32358));
    InMux I__4885 (
            .O(N__32373),
            .I(N__32355));
    InMux I__4884 (
            .O(N__32372),
            .I(N__32352));
    InMux I__4883 (
            .O(N__32371),
            .I(N__32349));
    Span4Mux_v I__4882 (
            .O(N__32368),
            .I(N__32346));
    InMux I__4881 (
            .O(N__32367),
            .I(N__32343));
    LocalMux I__4880 (
            .O(N__32364),
            .I(N__32334));
    LocalMux I__4879 (
            .O(N__32361),
            .I(N__32334));
    LocalMux I__4878 (
            .O(N__32358),
            .I(N__32334));
    LocalMux I__4877 (
            .O(N__32355),
            .I(N__32334));
    LocalMux I__4876 (
            .O(N__32352),
            .I(\c0.n13480 ));
    LocalMux I__4875 (
            .O(N__32349),
            .I(\c0.n13480 ));
    Odrv4 I__4874 (
            .O(N__32346),
            .I(\c0.n13480 ));
    LocalMux I__4873 (
            .O(N__32343),
            .I(\c0.n13480 ));
    Odrv4 I__4872 (
            .O(N__32334),
            .I(\c0.n13480 ));
    InMux I__4871 (
            .O(N__32323),
            .I(N__32320));
    LocalMux I__4870 (
            .O(N__32320),
            .I(N__32317));
    Span4Mux_h I__4869 (
            .O(N__32317),
            .I(N__32314));
    Odrv4 I__4868 (
            .O(N__32314),
            .I(\c0.n22078 ));
    CascadeMux I__4867 (
            .O(N__32311),
            .I(N__32306));
    CascadeMux I__4866 (
            .O(N__32310),
            .I(N__32303));
    CascadeMux I__4865 (
            .O(N__32309),
            .I(N__32299));
    InMux I__4864 (
            .O(N__32306),
            .I(N__32296));
    InMux I__4863 (
            .O(N__32303),
            .I(N__32293));
    CascadeMux I__4862 (
            .O(N__32302),
            .I(N__32290));
    InMux I__4861 (
            .O(N__32299),
            .I(N__32287));
    LocalMux I__4860 (
            .O(N__32296),
            .I(N__32283));
    LocalMux I__4859 (
            .O(N__32293),
            .I(N__32280));
    InMux I__4858 (
            .O(N__32290),
            .I(N__32277));
    LocalMux I__4857 (
            .O(N__32287),
            .I(N__32274));
    InMux I__4856 (
            .O(N__32286),
            .I(N__32270));
    Span4Mux_v I__4855 (
            .O(N__32283),
            .I(N__32263));
    Span4Mux_v I__4854 (
            .O(N__32280),
            .I(N__32263));
    LocalMux I__4853 (
            .O(N__32277),
            .I(N__32263));
    Span4Mux_h I__4852 (
            .O(N__32274),
            .I(N__32260));
    InMux I__4851 (
            .O(N__32273),
            .I(N__32257));
    LocalMux I__4850 (
            .O(N__32270),
            .I(encoder1_position_9));
    Odrv4 I__4849 (
            .O(N__32263),
            .I(encoder1_position_9));
    Odrv4 I__4848 (
            .O(N__32260),
            .I(encoder1_position_9));
    LocalMux I__4847 (
            .O(N__32257),
            .I(encoder1_position_9));
    InMux I__4846 (
            .O(N__32248),
            .I(N__32242));
    InMux I__4845 (
            .O(N__32247),
            .I(N__32237));
    InMux I__4844 (
            .O(N__32246),
            .I(N__32237));
    InMux I__4843 (
            .O(N__32245),
            .I(N__32234));
    LocalMux I__4842 (
            .O(N__32242),
            .I(N__32228));
    LocalMux I__4841 (
            .O(N__32237),
            .I(N__32228));
    LocalMux I__4840 (
            .O(N__32234),
            .I(N__32225));
    InMux I__4839 (
            .O(N__32233),
            .I(N__32222));
    Span4Mux_h I__4838 (
            .O(N__32228),
            .I(N__32219));
    Odrv12 I__4837 (
            .O(N__32225),
            .I(\c0.n21112 ));
    LocalMux I__4836 (
            .O(N__32222),
            .I(\c0.n21112 ));
    Odrv4 I__4835 (
            .O(N__32219),
            .I(\c0.n21112 ));
    InMux I__4834 (
            .O(N__32212),
            .I(N__32207));
    InMux I__4833 (
            .O(N__32211),
            .I(N__32201));
    InMux I__4832 (
            .O(N__32210),
            .I(N__32198));
    LocalMux I__4831 (
            .O(N__32207),
            .I(N__32195));
    InMux I__4830 (
            .O(N__32206),
            .I(N__32190));
    InMux I__4829 (
            .O(N__32205),
            .I(N__32190));
    InMux I__4828 (
            .O(N__32204),
            .I(N__32187));
    LocalMux I__4827 (
            .O(N__32201),
            .I(N__32179));
    LocalMux I__4826 (
            .O(N__32198),
            .I(N__32179));
    Span4Mux_h I__4825 (
            .O(N__32195),
            .I(N__32179));
    LocalMux I__4824 (
            .O(N__32190),
            .I(N__32176));
    LocalMux I__4823 (
            .O(N__32187),
            .I(N__32173));
    InMux I__4822 (
            .O(N__32186),
            .I(N__32170));
    Span4Mux_v I__4821 (
            .O(N__32179),
            .I(N__32167));
    Span4Mux_h I__4820 (
            .O(N__32176),
            .I(N__32162));
    Span4Mux_v I__4819 (
            .O(N__32173),
            .I(N__32162));
    LocalMux I__4818 (
            .O(N__32170),
            .I(N__32159));
    Odrv4 I__4817 (
            .O(N__32167),
            .I(\c0.n21253 ));
    Odrv4 I__4816 (
            .O(N__32162),
            .I(\c0.n21253 ));
    Odrv4 I__4815 (
            .O(N__32159),
            .I(\c0.n21253 ));
    CascadeMux I__4814 (
            .O(N__32152),
            .I(\c0.n20180_cascade_ ));
    InMux I__4813 (
            .O(N__32149),
            .I(N__32145));
    InMux I__4812 (
            .O(N__32148),
            .I(N__32142));
    LocalMux I__4811 (
            .O(N__32145),
            .I(N__32136));
    LocalMux I__4810 (
            .O(N__32142),
            .I(N__32136));
    InMux I__4809 (
            .O(N__32141),
            .I(N__32132));
    Span4Mux_v I__4808 (
            .O(N__32136),
            .I(N__32129));
    InMux I__4807 (
            .O(N__32135),
            .I(N__32126));
    LocalMux I__4806 (
            .O(N__32132),
            .I(N__32123));
    Odrv4 I__4805 (
            .O(N__32129),
            .I(\c0.data_out_frame_29__7__N_1144 ));
    LocalMux I__4804 (
            .O(N__32126),
            .I(\c0.data_out_frame_29__7__N_1144 ));
    Odrv4 I__4803 (
            .O(N__32123),
            .I(\c0.data_out_frame_29__7__N_1144 ));
    InMux I__4802 (
            .O(N__32116),
            .I(N__32110));
    InMux I__4801 (
            .O(N__32115),
            .I(N__32106));
    InMux I__4800 (
            .O(N__32114),
            .I(N__32101));
    InMux I__4799 (
            .O(N__32113),
            .I(N__32101));
    LocalMux I__4798 (
            .O(N__32110),
            .I(N__32097));
    InMux I__4797 (
            .O(N__32109),
            .I(N__32094));
    LocalMux I__4796 (
            .O(N__32106),
            .I(N__32089));
    LocalMux I__4795 (
            .O(N__32101),
            .I(N__32089));
    InMux I__4794 (
            .O(N__32100),
            .I(N__32086));
    Span4Mux_v I__4793 (
            .O(N__32097),
            .I(N__32083));
    LocalMux I__4792 (
            .O(N__32094),
            .I(N__32080));
    Span4Mux_h I__4791 (
            .O(N__32089),
            .I(N__32075));
    LocalMux I__4790 (
            .O(N__32086),
            .I(N__32075));
    Odrv4 I__4789 (
            .O(N__32083),
            .I(\c0.n20465 ));
    Odrv12 I__4788 (
            .O(N__32080),
            .I(\c0.n20465 ));
    Odrv4 I__4787 (
            .O(N__32075),
            .I(\c0.n20465 ));
    InMux I__4786 (
            .O(N__32068),
            .I(N__32065));
    LocalMux I__4785 (
            .O(N__32065),
            .I(N__32061));
    InMux I__4784 (
            .O(N__32064),
            .I(N__32058));
    Span4Mux_v I__4783 (
            .O(N__32061),
            .I(N__32055));
    LocalMux I__4782 (
            .O(N__32058),
            .I(data_out_frame_13_7));
    Odrv4 I__4781 (
            .O(N__32055),
            .I(data_out_frame_13_7));
    CascadeMux I__4780 (
            .O(N__32050),
            .I(N__32047));
    InMux I__4779 (
            .O(N__32047),
            .I(N__32043));
    CascadeMux I__4778 (
            .O(N__32046),
            .I(N__32040));
    LocalMux I__4777 (
            .O(N__32043),
            .I(N__32036));
    InMux I__4776 (
            .O(N__32040),
            .I(N__32030));
    InMux I__4775 (
            .O(N__32039),
            .I(N__32030));
    Span4Mux_h I__4774 (
            .O(N__32036),
            .I(N__32027));
    InMux I__4773 (
            .O(N__32035),
            .I(N__32024));
    LocalMux I__4772 (
            .O(N__32030),
            .I(N__32021));
    Odrv4 I__4771 (
            .O(N__32027),
            .I(\c0.n21056 ));
    LocalMux I__4770 (
            .O(N__32024),
            .I(\c0.n21056 ));
    Odrv4 I__4769 (
            .O(N__32021),
            .I(\c0.n21056 ));
    InMux I__4768 (
            .O(N__32014),
            .I(N__32010));
    InMux I__4767 (
            .O(N__32013),
            .I(N__32007));
    LocalMux I__4766 (
            .O(N__32010),
            .I(\c0.n22177 ));
    LocalMux I__4765 (
            .O(N__32007),
            .I(\c0.n22177 ));
    InMux I__4764 (
            .O(N__32002),
            .I(N__31999));
    LocalMux I__4763 (
            .O(N__31999),
            .I(\c0.n22072 ));
    CascadeMux I__4762 (
            .O(N__31996),
            .I(\c0.n22072_cascade_ ));
    InMux I__4761 (
            .O(N__31993),
            .I(N__31990));
    LocalMux I__4760 (
            .O(N__31990),
            .I(N__31985));
    InMux I__4759 (
            .O(N__31989),
            .I(N__31982));
    InMux I__4758 (
            .O(N__31988),
            .I(N__31979));
    Span4Mux_h I__4757 (
            .O(N__31985),
            .I(N__31974));
    LocalMux I__4756 (
            .O(N__31982),
            .I(N__31974));
    LocalMux I__4755 (
            .O(N__31979),
            .I(\c0.n22073 ));
    Odrv4 I__4754 (
            .O(N__31974),
            .I(\c0.n22073 ));
    InMux I__4753 (
            .O(N__31969),
            .I(N__31965));
    InMux I__4752 (
            .O(N__31968),
            .I(N__31961));
    LocalMux I__4751 (
            .O(N__31965),
            .I(N__31958));
    InMux I__4750 (
            .O(N__31964),
            .I(N__31953));
    LocalMux I__4749 (
            .O(N__31961),
            .I(N__31948));
    Span4Mux_v I__4748 (
            .O(N__31958),
            .I(N__31948));
    InMux I__4747 (
            .O(N__31957),
            .I(N__31943));
    InMux I__4746 (
            .O(N__31956),
            .I(N__31943));
    LocalMux I__4745 (
            .O(N__31953),
            .I(N__31940));
    Span4Mux_v I__4744 (
            .O(N__31948),
            .I(N__31935));
    LocalMux I__4743 (
            .O(N__31943),
            .I(N__31935));
    Odrv4 I__4742 (
            .O(N__31940),
            .I(\c0.n20175 ));
    Odrv4 I__4741 (
            .O(N__31935),
            .I(\c0.n20175 ));
    CascadeMux I__4740 (
            .O(N__31930),
            .I(\c0.n20249_cascade_ ));
    InMux I__4739 (
            .O(N__31927),
            .I(N__31923));
    InMux I__4738 (
            .O(N__31926),
            .I(N__31919));
    LocalMux I__4737 (
            .O(N__31923),
            .I(N__31916));
    InMux I__4736 (
            .O(N__31922),
            .I(N__31913));
    LocalMux I__4735 (
            .O(N__31919),
            .I(N__31909));
    Span4Mux_v I__4734 (
            .O(N__31916),
            .I(N__31904));
    LocalMux I__4733 (
            .O(N__31913),
            .I(N__31904));
    InMux I__4732 (
            .O(N__31912),
            .I(N__31901));
    Odrv4 I__4731 (
            .O(N__31909),
            .I(\c0.n12528 ));
    Odrv4 I__4730 (
            .O(N__31904),
            .I(\c0.n12528 ));
    LocalMux I__4729 (
            .O(N__31901),
            .I(\c0.n12528 ));
    InMux I__4728 (
            .O(N__31894),
            .I(N__31887));
    InMux I__4727 (
            .O(N__31893),
            .I(N__31887));
    CascadeMux I__4726 (
            .O(N__31892),
            .I(N__31883));
    LocalMux I__4725 (
            .O(N__31887),
            .I(N__31878));
    InMux I__4724 (
            .O(N__31886),
            .I(N__31872));
    InMux I__4723 (
            .O(N__31883),
            .I(N__31872));
    InMux I__4722 (
            .O(N__31882),
            .I(N__31867));
    InMux I__4721 (
            .O(N__31881),
            .I(N__31867));
    Span4Mux_h I__4720 (
            .O(N__31878),
            .I(N__31864));
    InMux I__4719 (
            .O(N__31877),
            .I(N__31861));
    LocalMux I__4718 (
            .O(N__31872),
            .I(\c0.n21065 ));
    LocalMux I__4717 (
            .O(N__31867),
            .I(\c0.n21065 ));
    Odrv4 I__4716 (
            .O(N__31864),
            .I(\c0.n21065 ));
    LocalMux I__4715 (
            .O(N__31861),
            .I(\c0.n21065 ));
    InMux I__4714 (
            .O(N__31852),
            .I(N__31849));
    LocalMux I__4713 (
            .O(N__31849),
            .I(N__31846));
    Span4Mux_h I__4712 (
            .O(N__31846),
            .I(N__31843));
    Odrv4 I__4711 (
            .O(N__31843),
            .I(\c0.n21842 ));
    InMux I__4710 (
            .O(N__31840),
            .I(N__31835));
    InMux I__4709 (
            .O(N__31839),
            .I(N__31832));
    CascadeMux I__4708 (
            .O(N__31838),
            .I(N__31829));
    LocalMux I__4707 (
            .O(N__31835),
            .I(N__31824));
    LocalMux I__4706 (
            .O(N__31832),
            .I(N__31824));
    InMux I__4705 (
            .O(N__31829),
            .I(N__31821));
    Span4Mux_h I__4704 (
            .O(N__31824),
            .I(N__31818));
    LocalMux I__4703 (
            .O(N__31821),
            .I(\c0.n20230 ));
    Odrv4 I__4702 (
            .O(N__31818),
            .I(\c0.n20230 ));
    InMux I__4701 (
            .O(N__31813),
            .I(N__31810));
    LocalMux I__4700 (
            .O(N__31810),
            .I(N__31807));
    Span12Mux_v I__4699 (
            .O(N__31807),
            .I(N__31804));
    Odrv12 I__4698 (
            .O(N__31804),
            .I(\c0.n6_adj_4394 ));
    CascadeMux I__4697 (
            .O(N__31801),
            .I(\c0.n6_adj_4497_cascade_ ));
    InMux I__4696 (
            .O(N__31798),
            .I(N__31794));
    InMux I__4695 (
            .O(N__31797),
            .I(N__31791));
    LocalMux I__4694 (
            .O(N__31794),
            .I(N__31788));
    LocalMux I__4693 (
            .O(N__31791),
            .I(N__31785));
    Span4Mux_h I__4692 (
            .O(N__31788),
            .I(N__31782));
    Odrv4 I__4691 (
            .O(N__31785),
            .I(\c0.n20151 ));
    Odrv4 I__4690 (
            .O(N__31782),
            .I(\c0.n20151 ));
    InMux I__4689 (
            .O(N__31777),
            .I(N__31774));
    LocalMux I__4688 (
            .O(N__31774),
            .I(\c0.data_out_frame_29_6 ));
    InMux I__4687 (
            .O(N__31771),
            .I(N__31767));
    InMux I__4686 (
            .O(N__31770),
            .I(N__31764));
    LocalMux I__4685 (
            .O(N__31767),
            .I(N__31761));
    LocalMux I__4684 (
            .O(N__31764),
            .I(N__31758));
    Span4Mux_h I__4683 (
            .O(N__31761),
            .I(N__31754));
    Span4Mux_v I__4682 (
            .O(N__31758),
            .I(N__31751));
    InMux I__4681 (
            .O(N__31757),
            .I(N__31748));
    Odrv4 I__4680 (
            .O(N__31754),
            .I(\c0.n21848 ));
    Odrv4 I__4679 (
            .O(N__31751),
            .I(\c0.n21848 ));
    LocalMux I__4678 (
            .O(N__31748),
            .I(\c0.n21848 ));
    InMux I__4677 (
            .O(N__31741),
            .I(N__31738));
    LocalMux I__4676 (
            .O(N__31738),
            .I(N__31735));
    Odrv4 I__4675 (
            .O(N__31735),
            .I(\c0.n20253 ));
    CascadeMux I__4674 (
            .O(N__31732),
            .I(\c0.n21852_cascade_ ));
    InMux I__4673 (
            .O(N__31729),
            .I(N__31723));
    InMux I__4672 (
            .O(N__31728),
            .I(N__31723));
    LocalMux I__4671 (
            .O(N__31723),
            .I(\c0.n22346 ));
    InMux I__4670 (
            .O(N__31720),
            .I(N__31714));
    InMux I__4669 (
            .O(N__31719),
            .I(N__31714));
    LocalMux I__4668 (
            .O(N__31714),
            .I(N__31711));
    Odrv12 I__4667 (
            .O(N__31711),
            .I(\c0.n22126 ));
    InMux I__4666 (
            .O(N__31708),
            .I(N__31704));
    InMux I__4665 (
            .O(N__31707),
            .I(N__31701));
    LocalMux I__4664 (
            .O(N__31704),
            .I(\c0.n20298 ));
    LocalMux I__4663 (
            .O(N__31701),
            .I(\c0.n20298 ));
    CascadeMux I__4662 (
            .O(N__31696),
            .I(\c0.n10_adj_4512_cascade_ ));
    CascadeMux I__4661 (
            .O(N__31693),
            .I(N__31689));
    InMux I__4660 (
            .O(N__31692),
            .I(N__31684));
    InMux I__4659 (
            .O(N__31689),
            .I(N__31679));
    InMux I__4658 (
            .O(N__31688),
            .I(N__31676));
    InMux I__4657 (
            .O(N__31687),
            .I(N__31673));
    LocalMux I__4656 (
            .O(N__31684),
            .I(N__31670));
    InMux I__4655 (
            .O(N__31683),
            .I(N__31667));
    InMux I__4654 (
            .O(N__31682),
            .I(N__31664));
    LocalMux I__4653 (
            .O(N__31679),
            .I(N__31657));
    LocalMux I__4652 (
            .O(N__31676),
            .I(N__31657));
    LocalMux I__4651 (
            .O(N__31673),
            .I(N__31657));
    Span4Mux_v I__4650 (
            .O(N__31670),
            .I(N__31653));
    LocalMux I__4649 (
            .O(N__31667),
            .I(N__31646));
    LocalMux I__4648 (
            .O(N__31664),
            .I(N__31646));
    Span4Mux_h I__4647 (
            .O(N__31657),
            .I(N__31646));
    InMux I__4646 (
            .O(N__31656),
            .I(N__31643));
    Odrv4 I__4645 (
            .O(N__31653),
            .I(\c0.n10496 ));
    Odrv4 I__4644 (
            .O(N__31646),
            .I(\c0.n10496 ));
    LocalMux I__4643 (
            .O(N__31643),
            .I(\c0.n10496 ));
    InMux I__4642 (
            .O(N__31636),
            .I(N__31627));
    InMux I__4641 (
            .O(N__31635),
            .I(N__31624));
    InMux I__4640 (
            .O(N__31634),
            .I(N__31618));
    InMux I__4639 (
            .O(N__31633),
            .I(N__31618));
    InMux I__4638 (
            .O(N__31632),
            .I(N__31613));
    InMux I__4637 (
            .O(N__31631),
            .I(N__31613));
    InMux I__4636 (
            .O(N__31630),
            .I(N__31610));
    LocalMux I__4635 (
            .O(N__31627),
            .I(N__31607));
    LocalMux I__4634 (
            .O(N__31624),
            .I(N__31604));
    InMux I__4633 (
            .O(N__31623),
            .I(N__31601));
    LocalMux I__4632 (
            .O(N__31618),
            .I(N__31594));
    LocalMux I__4631 (
            .O(N__31613),
            .I(N__31594));
    LocalMux I__4630 (
            .O(N__31610),
            .I(N__31594));
    Span4Mux_h I__4629 (
            .O(N__31607),
            .I(N__31587));
    Span4Mux_v I__4628 (
            .O(N__31604),
            .I(N__31587));
    LocalMux I__4627 (
            .O(N__31601),
            .I(N__31587));
    Odrv4 I__4626 (
            .O(N__31594),
            .I(\c0.n20274 ));
    Odrv4 I__4625 (
            .O(N__31587),
            .I(\c0.n20274 ));
    InMux I__4624 (
            .O(N__31582),
            .I(N__31579));
    LocalMux I__4623 (
            .O(N__31579),
            .I(N__31576));
    Span4Mux_v I__4622 (
            .O(N__31576),
            .I(N__31573));
    Odrv4 I__4621 (
            .O(N__31573),
            .I(\c0.n21231 ));
    InMux I__4620 (
            .O(N__31570),
            .I(N__31566));
    InMux I__4619 (
            .O(N__31569),
            .I(N__31562));
    LocalMux I__4618 (
            .O(N__31566),
            .I(N__31558));
    InMux I__4617 (
            .O(N__31565),
            .I(N__31555));
    LocalMux I__4616 (
            .O(N__31562),
            .I(N__31552));
    InMux I__4615 (
            .O(N__31561),
            .I(N__31549));
    Odrv4 I__4614 (
            .O(N__31558),
            .I(\c0.n22736 ));
    LocalMux I__4613 (
            .O(N__31555),
            .I(\c0.n22736 ));
    Odrv4 I__4612 (
            .O(N__31552),
            .I(\c0.n22736 ));
    LocalMux I__4611 (
            .O(N__31549),
            .I(\c0.n22736 ));
    CascadeMux I__4610 (
            .O(N__31540),
            .I(\c0.n21162_cascade_ ));
    InMux I__4609 (
            .O(N__31537),
            .I(N__31531));
    InMux I__4608 (
            .O(N__31536),
            .I(N__31531));
    LocalMux I__4607 (
            .O(N__31531),
            .I(\c0.n12526 ));
    InMux I__4606 (
            .O(N__31528),
            .I(N__31522));
    InMux I__4605 (
            .O(N__31527),
            .I(N__31522));
    LocalMux I__4604 (
            .O(N__31522),
            .I(\c0.n20201 ));
    CascadeMux I__4603 (
            .O(N__31519),
            .I(N__31516));
    InMux I__4602 (
            .O(N__31516),
            .I(N__31510));
    InMux I__4601 (
            .O(N__31515),
            .I(N__31510));
    LocalMux I__4600 (
            .O(N__31510),
            .I(N__31507));
    Odrv4 I__4599 (
            .O(N__31507),
            .I(\c0.n21876 ));
    CascadeMux I__4598 (
            .O(N__31504),
            .I(N__31501));
    InMux I__4597 (
            .O(N__31501),
            .I(N__31498));
    LocalMux I__4596 (
            .O(N__31498),
            .I(N__31495));
    Span4Mux_v I__4595 (
            .O(N__31495),
            .I(N__31492));
    Odrv4 I__4594 (
            .O(N__31492),
            .I(\c0.n24119 ));
    InMux I__4593 (
            .O(N__31489),
            .I(N__31486));
    LocalMux I__4592 (
            .O(N__31486),
            .I(N__31482));
    InMux I__4591 (
            .O(N__31485),
            .I(N__31479));
    Span4Mux_h I__4590 (
            .O(N__31482),
            .I(N__31476));
    LocalMux I__4589 (
            .O(N__31479),
            .I(N__31473));
    Odrv4 I__4588 (
            .O(N__31476),
            .I(\c0.n21050 ));
    Odrv12 I__4587 (
            .O(N__31473),
            .I(\c0.n21050 ));
    InMux I__4586 (
            .O(N__31468),
            .I(N__31465));
    LocalMux I__4585 (
            .O(N__31465),
            .I(\c0.n6_adj_4402 ));
    InMux I__4584 (
            .O(N__31462),
            .I(N__31459));
    LocalMux I__4583 (
            .O(N__31459),
            .I(N__31454));
    InMux I__4582 (
            .O(N__31458),
            .I(N__31451));
    InMux I__4581 (
            .O(N__31457),
            .I(N__31448));
    Odrv4 I__4580 (
            .O(N__31454),
            .I(\c0.n22188 ));
    LocalMux I__4579 (
            .O(N__31451),
            .I(\c0.n22188 ));
    LocalMux I__4578 (
            .O(N__31448),
            .I(\c0.n22188 ));
    CascadeMux I__4577 (
            .O(N__31441),
            .I(\c0.n20658_cascade_ ));
    InMux I__4576 (
            .O(N__31438),
            .I(N__31435));
    LocalMux I__4575 (
            .O(N__31435),
            .I(N__31431));
    InMux I__4574 (
            .O(N__31434),
            .I(N__31428));
    Span4Mux_h I__4573 (
            .O(N__31431),
            .I(N__31425));
    LocalMux I__4572 (
            .O(N__31428),
            .I(\c0.n22166 ));
    Odrv4 I__4571 (
            .O(N__31425),
            .I(\c0.n22166 ));
    CascadeMux I__4570 (
            .O(N__31420),
            .I(N__31412));
    CascadeMux I__4569 (
            .O(N__31419),
            .I(N__31409));
    CascadeMux I__4568 (
            .O(N__31418),
            .I(N__31406));
    CascadeMux I__4567 (
            .O(N__31417),
            .I(N__31401));
    CascadeMux I__4566 (
            .O(N__31416),
            .I(N__31398));
    InMux I__4565 (
            .O(N__31415),
            .I(N__31391));
    InMux I__4564 (
            .O(N__31412),
            .I(N__31391));
    InMux I__4563 (
            .O(N__31409),
            .I(N__31391));
    InMux I__4562 (
            .O(N__31406),
            .I(N__31386));
    InMux I__4561 (
            .O(N__31405),
            .I(N__31386));
    InMux I__4560 (
            .O(N__31404),
            .I(N__31383));
    InMux I__4559 (
            .O(N__31401),
            .I(N__31378));
    InMux I__4558 (
            .O(N__31398),
            .I(N__31378));
    LocalMux I__4557 (
            .O(N__31391),
            .I(N__31374));
    LocalMux I__4556 (
            .O(N__31386),
            .I(N__31367));
    LocalMux I__4555 (
            .O(N__31383),
            .I(N__31367));
    LocalMux I__4554 (
            .O(N__31378),
            .I(N__31367));
    InMux I__4553 (
            .O(N__31377),
            .I(N__31364));
    Span12Mux_h I__4552 (
            .O(N__31374),
            .I(N__31361));
    Span4Mux_v I__4551 (
            .O(N__31367),
            .I(N__31358));
    LocalMux I__4550 (
            .O(N__31364),
            .I(\c0.n10467 ));
    Odrv12 I__4549 (
            .O(N__31361),
            .I(\c0.n10467 ));
    Odrv4 I__4548 (
            .O(N__31358),
            .I(\c0.n10467 ));
    CascadeMux I__4547 (
            .O(N__31351),
            .I(N__31345));
    InMux I__4546 (
            .O(N__31350),
            .I(N__31342));
    CascadeMux I__4545 (
            .O(N__31349),
            .I(N__31338));
    CascadeMux I__4544 (
            .O(N__31348),
            .I(N__31334));
    InMux I__4543 (
            .O(N__31345),
            .I(N__31331));
    LocalMux I__4542 (
            .O(N__31342),
            .I(N__31328));
    InMux I__4541 (
            .O(N__31341),
            .I(N__31325));
    InMux I__4540 (
            .O(N__31338),
            .I(N__31322));
    InMux I__4539 (
            .O(N__31337),
            .I(N__31319));
    InMux I__4538 (
            .O(N__31334),
            .I(N__31316));
    LocalMux I__4537 (
            .O(N__31331),
            .I(N__31313));
    Span4Mux_v I__4536 (
            .O(N__31328),
            .I(N__31310));
    LocalMux I__4535 (
            .O(N__31325),
            .I(\c0.n22180 ));
    LocalMux I__4534 (
            .O(N__31322),
            .I(\c0.n22180 ));
    LocalMux I__4533 (
            .O(N__31319),
            .I(\c0.n22180 ));
    LocalMux I__4532 (
            .O(N__31316),
            .I(\c0.n22180 ));
    Odrv4 I__4531 (
            .O(N__31313),
            .I(\c0.n22180 ));
    Odrv4 I__4530 (
            .O(N__31310),
            .I(\c0.n22180 ));
    InMux I__4529 (
            .O(N__31297),
            .I(N__31289));
    InMux I__4528 (
            .O(N__31296),
            .I(N__31289));
    InMux I__4527 (
            .O(N__31295),
            .I(N__31286));
    InMux I__4526 (
            .O(N__31294),
            .I(N__31282));
    LocalMux I__4525 (
            .O(N__31289),
            .I(N__31277));
    LocalMux I__4524 (
            .O(N__31286),
            .I(N__31277));
    InMux I__4523 (
            .O(N__31285),
            .I(N__31274));
    LocalMux I__4522 (
            .O(N__31282),
            .I(N__31269));
    Span4Mux_v I__4521 (
            .O(N__31277),
            .I(N__31266));
    LocalMux I__4520 (
            .O(N__31274),
            .I(N__31263));
    InMux I__4519 (
            .O(N__31273),
            .I(N__31258));
    InMux I__4518 (
            .O(N__31272),
            .I(N__31258));
    Span4Mux_h I__4517 (
            .O(N__31269),
            .I(N__31253));
    Span4Mux_v I__4516 (
            .O(N__31266),
            .I(N__31249));
    Span4Mux_h I__4515 (
            .O(N__31263),
            .I(N__31244));
    LocalMux I__4514 (
            .O(N__31258),
            .I(N__31244));
    InMux I__4513 (
            .O(N__31257),
            .I(N__31241));
    InMux I__4512 (
            .O(N__31256),
            .I(N__31238));
    Span4Mux_v I__4511 (
            .O(N__31253),
            .I(N__31235));
    InMux I__4510 (
            .O(N__31252),
            .I(N__31232));
    Odrv4 I__4509 (
            .O(N__31249),
            .I(\c0.n20330 ));
    Odrv4 I__4508 (
            .O(N__31244),
            .I(\c0.n20330 ));
    LocalMux I__4507 (
            .O(N__31241),
            .I(\c0.n20330 ));
    LocalMux I__4506 (
            .O(N__31238),
            .I(\c0.n20330 ));
    Odrv4 I__4505 (
            .O(N__31235),
            .I(\c0.n20330 ));
    LocalMux I__4504 (
            .O(N__31232),
            .I(\c0.n20330 ));
    CascadeMux I__4503 (
            .O(N__31219),
            .I(N__31214));
    InMux I__4502 (
            .O(N__31218),
            .I(N__31210));
    InMux I__4501 (
            .O(N__31217),
            .I(N__31203));
    InMux I__4500 (
            .O(N__31214),
            .I(N__31203));
    InMux I__4499 (
            .O(N__31213),
            .I(N__31200));
    LocalMux I__4498 (
            .O(N__31210),
            .I(N__31197));
    InMux I__4497 (
            .O(N__31209),
            .I(N__31194));
    InMux I__4496 (
            .O(N__31208),
            .I(N__31191));
    LocalMux I__4495 (
            .O(N__31203),
            .I(N__31185));
    LocalMux I__4494 (
            .O(N__31200),
            .I(N__31185));
    Span4Mux_v I__4493 (
            .O(N__31197),
            .I(N__31182));
    LocalMux I__4492 (
            .O(N__31194),
            .I(N__31177));
    LocalMux I__4491 (
            .O(N__31191),
            .I(N__31177));
    InMux I__4490 (
            .O(N__31190),
            .I(N__31174));
    Span4Mux_h I__4489 (
            .O(N__31185),
            .I(N__31171));
    Span4Mux_h I__4488 (
            .O(N__31182),
            .I(N__31166));
    Span4Mux_v I__4487 (
            .O(N__31177),
            .I(N__31166));
    LocalMux I__4486 (
            .O(N__31174),
            .I(\c0.n10434 ));
    Odrv4 I__4485 (
            .O(N__31171),
            .I(\c0.n10434 ));
    Odrv4 I__4484 (
            .O(N__31166),
            .I(\c0.n10434 ));
    InMux I__4483 (
            .O(N__31159),
            .I(N__31153));
    InMux I__4482 (
            .O(N__31158),
            .I(N__31153));
    LocalMux I__4481 (
            .O(N__31153),
            .I(N__31148));
    InMux I__4480 (
            .O(N__31152),
            .I(N__31145));
    InMux I__4479 (
            .O(N__31151),
            .I(N__31142));
    Span4Mux_h I__4478 (
            .O(N__31148),
            .I(N__31139));
    LocalMux I__4477 (
            .O(N__31145),
            .I(\c0.n10513 ));
    LocalMux I__4476 (
            .O(N__31142),
            .I(\c0.n10513 ));
    Odrv4 I__4475 (
            .O(N__31139),
            .I(\c0.n10513 ));
    InMux I__4474 (
            .O(N__31132),
            .I(N__31123));
    InMux I__4473 (
            .O(N__31131),
            .I(N__31123));
    InMux I__4472 (
            .O(N__31130),
            .I(N__31120));
    InMux I__4471 (
            .O(N__31129),
            .I(N__31115));
    InMux I__4470 (
            .O(N__31128),
            .I(N__31115));
    LocalMux I__4469 (
            .O(N__31123),
            .I(N__31110));
    LocalMux I__4468 (
            .O(N__31120),
            .I(N__31110));
    LocalMux I__4467 (
            .O(N__31115),
            .I(N__31107));
    Odrv4 I__4466 (
            .O(N__31110),
            .I(\c0.n21189 ));
    Odrv4 I__4465 (
            .O(N__31107),
            .I(\c0.n21189 ));
    CascadeMux I__4464 (
            .O(N__31102),
            .I(N__31099));
    InMux I__4463 (
            .O(N__31099),
            .I(N__31096));
    LocalMux I__4462 (
            .O(N__31096),
            .I(\c0.n21135 ));
    InMux I__4461 (
            .O(N__31093),
            .I(N__31090));
    LocalMux I__4460 (
            .O(N__31090),
            .I(N__31085));
    InMux I__4459 (
            .O(N__31089),
            .I(N__31082));
    InMux I__4458 (
            .O(N__31088),
            .I(N__31079));
    Odrv12 I__4457 (
            .O(N__31085),
            .I(\c0.n21219 ));
    LocalMux I__4456 (
            .O(N__31082),
            .I(\c0.n21219 ));
    LocalMux I__4455 (
            .O(N__31079),
            .I(\c0.n21219 ));
    InMux I__4454 (
            .O(N__31072),
            .I(N__31067));
    InMux I__4453 (
            .O(N__31071),
            .I(N__31064));
    InMux I__4452 (
            .O(N__31070),
            .I(N__31061));
    LocalMux I__4451 (
            .O(N__31067),
            .I(\c0.n21811 ));
    LocalMux I__4450 (
            .O(N__31064),
            .I(\c0.n21811 ));
    LocalMux I__4449 (
            .O(N__31061),
            .I(\c0.n21811 ));
    CascadeMux I__4448 (
            .O(N__31054),
            .I(\c0.n21135_cascade_ ));
    InMux I__4447 (
            .O(N__31051),
            .I(\c0.tx.n19545 ));
    InMux I__4446 (
            .O(N__31048),
            .I(N__31044));
    InMux I__4445 (
            .O(N__31047),
            .I(N__31039));
    LocalMux I__4444 (
            .O(N__31044),
            .I(N__31036));
    InMux I__4443 (
            .O(N__31043),
            .I(N__31031));
    InMux I__4442 (
            .O(N__31042),
            .I(N__31031));
    LocalMux I__4441 (
            .O(N__31039),
            .I(r_Clock_Count_7));
    Odrv4 I__4440 (
            .O(N__31036),
            .I(r_Clock_Count_7));
    LocalMux I__4439 (
            .O(N__31031),
            .I(r_Clock_Count_7));
    InMux I__4438 (
            .O(N__31024),
            .I(N__31021));
    LocalMux I__4437 (
            .O(N__31021),
            .I(N__31018));
    Odrv4 I__4436 (
            .O(N__31018),
            .I(n314));
    InMux I__4435 (
            .O(N__31015),
            .I(\c0.tx.n19546 ));
    InMux I__4434 (
            .O(N__31012),
            .I(bfn_13_22_0_));
    InMux I__4433 (
            .O(N__31009),
            .I(N__31006));
    LocalMux I__4432 (
            .O(N__31006),
            .I(\c0.n12878 ));
    SRMux I__4431 (
            .O(N__31003),
            .I(N__31000));
    LocalMux I__4430 (
            .O(N__31000),
            .I(N__30997));
    Span4Mux_h I__4429 (
            .O(N__30997),
            .I(N__30994));
    Span4Mux_h I__4428 (
            .O(N__30994),
            .I(N__30991));
    Odrv4 I__4427 (
            .O(N__30991),
            .I(\c0.n21360 ));
    SRMux I__4426 (
            .O(N__30988),
            .I(N__30985));
    LocalMux I__4425 (
            .O(N__30985),
            .I(\c0.n21356 ));
    InMux I__4424 (
            .O(N__30982),
            .I(N__30978));
    InMux I__4423 (
            .O(N__30981),
            .I(N__30975));
    LocalMux I__4422 (
            .O(N__30978),
            .I(N__30972));
    LocalMux I__4421 (
            .O(N__30975),
            .I(\c0.n22317 ));
    Odrv4 I__4420 (
            .O(N__30972),
            .I(\c0.n22317 ));
    InMux I__4419 (
            .O(N__30967),
            .I(N__30964));
    LocalMux I__4418 (
            .O(N__30964),
            .I(\c0.n6_adj_4305 ));
    CascadeMux I__4417 (
            .O(N__30961),
            .I(\c0.tx.n6_cascade_ ));
    InMux I__4416 (
            .O(N__30958),
            .I(N__30955));
    LocalMux I__4415 (
            .O(N__30955),
            .I(\c0.tx.n31 ));
    CascadeMux I__4414 (
            .O(N__30952),
            .I(\c0.tx.n31_cascade_ ));
    InMux I__4413 (
            .O(N__30949),
            .I(N__30946));
    LocalMux I__4412 (
            .O(N__30946),
            .I(\c0.tx.n47 ));
    CascadeMux I__4411 (
            .O(N__30943),
            .I(N__30940));
    InMux I__4410 (
            .O(N__30940),
            .I(N__30937));
    LocalMux I__4409 (
            .O(N__30937),
            .I(\c0.tx.n10 ));
    InMux I__4408 (
            .O(N__30934),
            .I(N__30930));
    InMux I__4407 (
            .O(N__30933),
            .I(N__30926));
    LocalMux I__4406 (
            .O(N__30930),
            .I(N__30923));
    InMux I__4405 (
            .O(N__30929),
            .I(N__30920));
    LocalMux I__4404 (
            .O(N__30926),
            .I(N__30915));
    Span4Mux_v I__4403 (
            .O(N__30923),
            .I(N__30915));
    LocalMux I__4402 (
            .O(N__30920),
            .I(\c0.tx.r_Clock_Count_0 ));
    Odrv4 I__4401 (
            .O(N__30915),
            .I(\c0.tx.r_Clock_Count_0 ));
    InMux I__4400 (
            .O(N__30910),
            .I(N__30907));
    LocalMux I__4399 (
            .O(N__30907),
            .I(N__30904));
    Odrv12 I__4398 (
            .O(N__30904),
            .I(\c0.tx.n23960 ));
    InMux I__4397 (
            .O(N__30901),
            .I(bfn_13_21_0_));
    InMux I__4396 (
            .O(N__30898),
            .I(N__30893));
    InMux I__4395 (
            .O(N__30897),
            .I(N__30890));
    InMux I__4394 (
            .O(N__30896),
            .I(N__30887));
    LocalMux I__4393 (
            .O(N__30893),
            .I(\c0.tx.r_Clock_Count_1 ));
    LocalMux I__4392 (
            .O(N__30890),
            .I(\c0.tx.r_Clock_Count_1 ));
    LocalMux I__4391 (
            .O(N__30887),
            .I(\c0.tx.r_Clock_Count_1 ));
    InMux I__4390 (
            .O(N__30880),
            .I(N__30877));
    LocalMux I__4389 (
            .O(N__30877),
            .I(\c0.tx.n23961 ));
    InMux I__4388 (
            .O(N__30874),
            .I(\c0.tx.n19540 ));
    InMux I__4387 (
            .O(N__30871),
            .I(N__30866));
    InMux I__4386 (
            .O(N__30870),
            .I(N__30863));
    InMux I__4385 (
            .O(N__30869),
            .I(N__30860));
    LocalMux I__4384 (
            .O(N__30866),
            .I(\c0.tx.r_Clock_Count_2 ));
    LocalMux I__4383 (
            .O(N__30863),
            .I(\c0.tx.r_Clock_Count_2 ));
    LocalMux I__4382 (
            .O(N__30860),
            .I(\c0.tx.r_Clock_Count_2 ));
    InMux I__4381 (
            .O(N__30853),
            .I(N__30850));
    LocalMux I__4380 (
            .O(N__30850),
            .I(\c0.tx.n23958 ));
    InMux I__4379 (
            .O(N__30847),
            .I(\c0.tx.n19541 ));
    InMux I__4378 (
            .O(N__30844),
            .I(N__30839));
    InMux I__4377 (
            .O(N__30843),
            .I(N__30836));
    InMux I__4376 (
            .O(N__30842),
            .I(N__30833));
    LocalMux I__4375 (
            .O(N__30839),
            .I(\c0.tx.r_Clock_Count_3 ));
    LocalMux I__4374 (
            .O(N__30836),
            .I(\c0.tx.r_Clock_Count_3 ));
    LocalMux I__4373 (
            .O(N__30833),
            .I(\c0.tx.r_Clock_Count_3 ));
    InMux I__4372 (
            .O(N__30826),
            .I(N__30823));
    LocalMux I__4371 (
            .O(N__30823),
            .I(\c0.tx.n23963 ));
    InMux I__4370 (
            .O(N__30820),
            .I(\c0.tx.n19542 ));
    InMux I__4369 (
            .O(N__30817),
            .I(N__30813));
    InMux I__4368 (
            .O(N__30816),
            .I(N__30810));
    LocalMux I__4367 (
            .O(N__30813),
            .I(N__30804));
    LocalMux I__4366 (
            .O(N__30810),
            .I(N__30804));
    InMux I__4365 (
            .O(N__30809),
            .I(N__30801));
    Span4Mux_v I__4364 (
            .O(N__30804),
            .I(N__30798));
    LocalMux I__4363 (
            .O(N__30801),
            .I(\c0.tx.r_Clock_Count_4 ));
    Odrv4 I__4362 (
            .O(N__30798),
            .I(\c0.tx.r_Clock_Count_4 ));
    InMux I__4361 (
            .O(N__30793),
            .I(N__30790));
    LocalMux I__4360 (
            .O(N__30790),
            .I(N__30787));
    Odrv12 I__4359 (
            .O(N__30787),
            .I(\c0.tx.n23953 ));
    InMux I__4358 (
            .O(N__30784),
            .I(\c0.tx.n19543 ));
    InMux I__4357 (
            .O(N__30781),
            .I(N__30775));
    InMux I__4356 (
            .O(N__30780),
            .I(N__30772));
    InMux I__4355 (
            .O(N__30779),
            .I(N__30767));
    InMux I__4354 (
            .O(N__30778),
            .I(N__30767));
    LocalMux I__4353 (
            .O(N__30775),
            .I(r_Clock_Count_5));
    LocalMux I__4352 (
            .O(N__30772),
            .I(r_Clock_Count_5));
    LocalMux I__4351 (
            .O(N__30767),
            .I(r_Clock_Count_5));
    InMux I__4350 (
            .O(N__30760),
            .I(N__30757));
    LocalMux I__4349 (
            .O(N__30757),
            .I(n316));
    InMux I__4348 (
            .O(N__30754),
            .I(\c0.tx.n19544 ));
    CascadeMux I__4347 (
            .O(N__30751),
            .I(o_Tx_Serial_N_3783_cascade_));
    InMux I__4346 (
            .O(N__30748),
            .I(N__30745));
    LocalMux I__4345 (
            .O(N__30745),
            .I(N__30742));
    Span4Mux_v I__4344 (
            .O(N__30742),
            .I(N__30739));
    Odrv4 I__4343 (
            .O(N__30739),
            .I(\c0.tx.n12 ));
    CascadeMux I__4342 (
            .O(N__30736),
            .I(N__30732));
    InMux I__4341 (
            .O(N__30735),
            .I(N__30722));
    InMux I__4340 (
            .O(N__30732),
            .I(N__30722));
    InMux I__4339 (
            .O(N__30731),
            .I(N__30722));
    InMux I__4338 (
            .O(N__30730),
            .I(N__30715));
    InMux I__4337 (
            .O(N__30729),
            .I(N__30715));
    LocalMux I__4336 (
            .O(N__30722),
            .I(N__30712));
    CascadeMux I__4335 (
            .O(N__30721),
            .I(N__30708));
    InMux I__4334 (
            .O(N__30720),
            .I(N__30700));
    LocalMux I__4333 (
            .O(N__30715),
            .I(N__30697));
    Span4Mux_h I__4332 (
            .O(N__30712),
            .I(N__30694));
    InMux I__4331 (
            .O(N__30711),
            .I(N__30691));
    InMux I__4330 (
            .O(N__30708),
            .I(N__30684));
    InMux I__4329 (
            .O(N__30707),
            .I(N__30684));
    InMux I__4328 (
            .O(N__30706),
            .I(N__30684));
    InMux I__4327 (
            .O(N__30705),
            .I(N__30677));
    InMux I__4326 (
            .O(N__30704),
            .I(N__30677));
    InMux I__4325 (
            .O(N__30703),
            .I(N__30677));
    LocalMux I__4324 (
            .O(N__30700),
            .I(r_SM_Main_1_adj_4550));
    Odrv12 I__4323 (
            .O(N__30697),
            .I(r_SM_Main_1_adj_4550));
    Odrv4 I__4322 (
            .O(N__30694),
            .I(r_SM_Main_1_adj_4550));
    LocalMux I__4321 (
            .O(N__30691),
            .I(r_SM_Main_1_adj_4550));
    LocalMux I__4320 (
            .O(N__30684),
            .I(r_SM_Main_1_adj_4550));
    LocalMux I__4319 (
            .O(N__30677),
            .I(r_SM_Main_1_adj_4550));
    CascadeMux I__4318 (
            .O(N__30664),
            .I(\c0.tx.n6_adj_4214_cascade_ ));
    CascadeMux I__4317 (
            .O(N__30661),
            .I(N__30657));
    InMux I__4316 (
            .O(N__30660),
            .I(N__30654));
    InMux I__4315 (
            .O(N__30657),
            .I(N__30651));
    LocalMux I__4314 (
            .O(N__30654),
            .I(N__30645));
    LocalMux I__4313 (
            .O(N__30651),
            .I(N__30645));
    InMux I__4312 (
            .O(N__30650),
            .I(N__30639));
    Span4Mux_h I__4311 (
            .O(N__30645),
            .I(N__30636));
    InMux I__4310 (
            .O(N__30644),
            .I(N__30629));
    InMux I__4309 (
            .O(N__30643),
            .I(N__30629));
    InMux I__4308 (
            .O(N__30642),
            .I(N__30629));
    LocalMux I__4307 (
            .O(N__30639),
            .I(\c0.tx.n16630 ));
    Odrv4 I__4306 (
            .O(N__30636),
            .I(\c0.tx.n16630 ));
    LocalMux I__4305 (
            .O(N__30629),
            .I(\c0.tx.n16630 ));
    CascadeMux I__4304 (
            .O(N__30622),
            .I(n8_cascade_));
    InMux I__4303 (
            .O(N__30619),
            .I(N__30615));
    InMux I__4302 (
            .O(N__30618),
            .I(N__30612));
    LocalMux I__4301 (
            .O(N__30615),
            .I(N__30608));
    LocalMux I__4300 (
            .O(N__30612),
            .I(N__30605));
    InMux I__4299 (
            .O(N__30611),
            .I(N__30602));
    Span12Mux_h I__4298 (
            .O(N__30608),
            .I(N__30597));
    Sp12to4 I__4297 (
            .O(N__30605),
            .I(N__30597));
    LocalMux I__4296 (
            .O(N__30602),
            .I(data_in_0_2));
    Odrv12 I__4295 (
            .O(N__30597),
            .I(data_in_0_2));
    InMux I__4294 (
            .O(N__30592),
            .I(N__30588));
    InMux I__4293 (
            .O(N__30591),
            .I(N__30585));
    LocalMux I__4292 (
            .O(N__30588),
            .I(\c0.n13006 ));
    LocalMux I__4291 (
            .O(N__30585),
            .I(\c0.n13006 ));
    InMux I__4290 (
            .O(N__30580),
            .I(N__30576));
    InMux I__4289 (
            .O(N__30579),
            .I(N__30573));
    LocalMux I__4288 (
            .O(N__30576),
            .I(\c0.n21767 ));
    LocalMux I__4287 (
            .O(N__30573),
            .I(\c0.n21767 ));
    InMux I__4286 (
            .O(N__30568),
            .I(N__30565));
    LocalMux I__4285 (
            .O(N__30565),
            .I(N__30562));
    Odrv4 I__4284 (
            .O(N__30562),
            .I(\c0.tx.n14296 ));
    CascadeMux I__4283 (
            .O(N__30559),
            .I(N__30554));
    CascadeMux I__4282 (
            .O(N__30558),
            .I(N__30551));
    InMux I__4281 (
            .O(N__30557),
            .I(N__30547));
    InMux I__4280 (
            .O(N__30554),
            .I(N__30544));
    InMux I__4279 (
            .O(N__30551),
            .I(N__30541));
    InMux I__4278 (
            .O(N__30550),
            .I(N__30538));
    LocalMux I__4277 (
            .O(N__30547),
            .I(N__30535));
    LocalMux I__4276 (
            .O(N__30544),
            .I(data_in_1_0));
    LocalMux I__4275 (
            .O(N__30541),
            .I(data_in_1_0));
    LocalMux I__4274 (
            .O(N__30538),
            .I(data_in_1_0));
    Odrv4 I__4273 (
            .O(N__30535),
            .I(data_in_1_0));
    InMux I__4272 (
            .O(N__30526),
            .I(N__30522));
    InMux I__4271 (
            .O(N__30525),
            .I(N__30519));
    LocalMux I__4270 (
            .O(N__30522),
            .I(data_in_0_0));
    LocalMux I__4269 (
            .O(N__30519),
            .I(data_in_0_0));
    CascadeMux I__4268 (
            .O(N__30514),
            .I(N__30510));
    InMux I__4267 (
            .O(N__30513),
            .I(N__30505));
    InMux I__4266 (
            .O(N__30510),
            .I(N__30505));
    LocalMux I__4265 (
            .O(N__30505),
            .I(data_in_0_4));
    InMux I__4264 (
            .O(N__30502),
            .I(N__30499));
    LocalMux I__4263 (
            .O(N__30499),
            .I(N__30495));
    InMux I__4262 (
            .O(N__30498),
            .I(N__30491));
    Span4Mux_v I__4261 (
            .O(N__30495),
            .I(N__30488));
    InMux I__4260 (
            .O(N__30494),
            .I(N__30485));
    LocalMux I__4259 (
            .O(N__30491),
            .I(data_in_1_7));
    Odrv4 I__4258 (
            .O(N__30488),
            .I(data_in_1_7));
    LocalMux I__4257 (
            .O(N__30485),
            .I(data_in_1_7));
    InMux I__4256 (
            .O(N__30478),
            .I(N__30475));
    LocalMux I__4255 (
            .O(N__30475),
            .I(\c0.n10_adj_4494 ));
    CascadeMux I__4254 (
            .O(N__30472),
            .I(N__30469));
    InMux I__4253 (
            .O(N__30469),
            .I(N__30466));
    LocalMux I__4252 (
            .O(N__30466),
            .I(N__30463));
    Odrv4 I__4251 (
            .O(N__30463),
            .I(\c0.n16_adj_4476 ));
    InMux I__4250 (
            .O(N__30460),
            .I(N__30457));
    LocalMux I__4249 (
            .O(N__30457),
            .I(\c0.n17_adj_4477 ));
    InMux I__4248 (
            .O(N__30454),
            .I(N__30447));
    CascadeMux I__4247 (
            .O(N__30453),
            .I(N__30444));
    InMux I__4246 (
            .O(N__30452),
            .I(N__30436));
    InMux I__4245 (
            .O(N__30451),
            .I(N__30436));
    InMux I__4244 (
            .O(N__30450),
            .I(N__30436));
    LocalMux I__4243 (
            .O(N__30447),
            .I(N__30433));
    InMux I__4242 (
            .O(N__30444),
            .I(N__30427));
    InMux I__4241 (
            .O(N__30443),
            .I(N__30427));
    LocalMux I__4240 (
            .O(N__30436),
            .I(N__30424));
    Span4Mux_h I__4239 (
            .O(N__30433),
            .I(N__30421));
    InMux I__4238 (
            .O(N__30432),
            .I(N__30418));
    LocalMux I__4237 (
            .O(N__30427),
            .I(r_Bit_Index_0_adj_4553));
    Odrv4 I__4236 (
            .O(N__30424),
            .I(r_Bit_Index_0_adj_4553));
    Odrv4 I__4235 (
            .O(N__30421),
            .I(r_Bit_Index_0_adj_4553));
    LocalMux I__4234 (
            .O(N__30418),
            .I(r_Bit_Index_0_adj_4553));
    InMux I__4233 (
            .O(N__30409),
            .I(N__30406));
    LocalMux I__4232 (
            .O(N__30406),
            .I(N__30403));
    Odrv4 I__4231 (
            .O(N__30403),
            .I(n24192));
    InMux I__4230 (
            .O(N__30400),
            .I(N__30397));
    LocalMux I__4229 (
            .O(N__30397),
            .I(N__30394));
    Span4Mux_h I__4228 (
            .O(N__30394),
            .I(N__30391));
    Odrv4 I__4227 (
            .O(N__30391),
            .I(n24198));
    InMux I__4226 (
            .O(N__30388),
            .I(N__30385));
    LocalMux I__4225 (
            .O(N__30385),
            .I(N__30381));
    InMux I__4224 (
            .O(N__30384),
            .I(N__30378));
    Span4Mux_h I__4223 (
            .O(N__30381),
            .I(N__30375));
    LocalMux I__4222 (
            .O(N__30378),
            .I(data_out_frame_6_4));
    Odrv4 I__4221 (
            .O(N__30375),
            .I(data_out_frame_6_4));
    InMux I__4220 (
            .O(N__30370),
            .I(N__30367));
    LocalMux I__4219 (
            .O(N__30367),
            .I(N__30363));
    InMux I__4218 (
            .O(N__30366),
            .I(N__30360));
    Odrv4 I__4217 (
            .O(N__30363),
            .I(\c0.n13003 ));
    LocalMux I__4216 (
            .O(N__30360),
            .I(\c0.n13003 ));
    InMux I__4215 (
            .O(N__30355),
            .I(N__30352));
    LocalMux I__4214 (
            .O(N__30352),
            .I(\c0.n19_adj_4367 ));
    CascadeMux I__4213 (
            .O(N__30349),
            .I(\c0.n20_adj_4362_cascade_ ));
    InMux I__4212 (
            .O(N__30346),
            .I(N__30343));
    LocalMux I__4211 (
            .O(N__30343),
            .I(\c0.n23834 ));
    InMux I__4210 (
            .O(N__30340),
            .I(N__30335));
    InMux I__4209 (
            .O(N__30339),
            .I(N__30332));
    InMux I__4208 (
            .O(N__30338),
            .I(N__30329));
    LocalMux I__4207 (
            .O(N__30335),
            .I(N__30325));
    LocalMux I__4206 (
            .O(N__30332),
            .I(N__30322));
    LocalMux I__4205 (
            .O(N__30329),
            .I(N__30319));
    InMux I__4204 (
            .O(N__30328),
            .I(N__30316));
    Span4Mux_v I__4203 (
            .O(N__30325),
            .I(N__30313));
    Span4Mux_h I__4202 (
            .O(N__30322),
            .I(N__30310));
    Odrv12 I__4201 (
            .O(N__30319),
            .I(data_in_1_2));
    LocalMux I__4200 (
            .O(N__30316),
            .I(data_in_1_2));
    Odrv4 I__4199 (
            .O(N__30313),
            .I(data_in_1_2));
    Odrv4 I__4198 (
            .O(N__30310),
            .I(data_in_1_2));
    CascadeMux I__4197 (
            .O(N__30301),
            .I(N__30296));
    InMux I__4196 (
            .O(N__30300),
            .I(N__30293));
    InMux I__4195 (
            .O(N__30299),
            .I(N__30288));
    InMux I__4194 (
            .O(N__30296),
            .I(N__30288));
    LocalMux I__4193 (
            .O(N__30293),
            .I(data_in_0_5));
    LocalMux I__4192 (
            .O(N__30288),
            .I(data_in_0_5));
    InMux I__4191 (
            .O(N__30283),
            .I(N__30280));
    LocalMux I__4190 (
            .O(N__30280),
            .I(N__30274));
    InMux I__4189 (
            .O(N__30279),
            .I(N__30269));
    InMux I__4188 (
            .O(N__30278),
            .I(N__30269));
    InMux I__4187 (
            .O(N__30277),
            .I(N__30266));
    Odrv12 I__4186 (
            .O(N__30274),
            .I(data_in_1_6));
    LocalMux I__4185 (
            .O(N__30269),
            .I(data_in_1_6));
    LocalMux I__4184 (
            .O(N__30266),
            .I(data_in_1_6));
    CascadeMux I__4183 (
            .O(N__30259),
            .I(\c0.n17_adj_4479_cascade_ ));
    CascadeMux I__4182 (
            .O(N__30256),
            .I(N__30253));
    InMux I__4181 (
            .O(N__30253),
            .I(N__30249));
    InMux I__4180 (
            .O(N__30252),
            .I(N__30246));
    LocalMux I__4179 (
            .O(N__30249),
            .I(\c0.n13023 ));
    LocalMux I__4178 (
            .O(N__30246),
            .I(\c0.n13023 ));
    CascadeMux I__4177 (
            .O(N__30241),
            .I(\c0.n21914_cascade_ ));
    InMux I__4176 (
            .O(N__30238),
            .I(N__30235));
    LocalMux I__4175 (
            .O(N__30235),
            .I(\c0.n21_adj_4320 ));
    CascadeMux I__4174 (
            .O(N__30232),
            .I(N__30228));
    InMux I__4173 (
            .O(N__30231),
            .I(N__30225));
    InMux I__4172 (
            .O(N__30228),
            .I(N__30222));
    LocalMux I__4171 (
            .O(N__30225),
            .I(N__30219));
    LocalMux I__4170 (
            .O(N__30222),
            .I(data_out_frame_8_4));
    Odrv12 I__4169 (
            .O(N__30219),
            .I(data_out_frame_8_4));
    CascadeMux I__4168 (
            .O(N__30214),
            .I(N__30211));
    InMux I__4167 (
            .O(N__30211),
            .I(N__30208));
    LocalMux I__4166 (
            .O(N__30208),
            .I(N__30205));
    Span4Mux_h I__4165 (
            .O(N__30205),
            .I(N__30202));
    Span4Mux_h I__4164 (
            .O(N__30202),
            .I(N__30199));
    Odrv4 I__4163 (
            .O(N__30199),
            .I(\c0.n23880 ));
    CascadeMux I__4162 (
            .O(N__30196),
            .I(N__30193));
    InMux I__4161 (
            .O(N__30193),
            .I(N__30187));
    InMux I__4160 (
            .O(N__30192),
            .I(N__30187));
    LocalMux I__4159 (
            .O(N__30187),
            .I(data_out_frame_9_4));
    InMux I__4158 (
            .O(N__30184),
            .I(N__30181));
    LocalMux I__4157 (
            .O(N__30181),
            .I(N__30178));
    Odrv4 I__4156 (
            .O(N__30178),
            .I(n2178));
    CascadeMux I__4155 (
            .O(N__30175),
            .I(N__30172));
    InMux I__4154 (
            .O(N__30172),
            .I(N__30168));
    CascadeMux I__4153 (
            .O(N__30171),
            .I(N__30165));
    LocalMux I__4152 (
            .O(N__30168),
            .I(N__30160));
    InMux I__4151 (
            .O(N__30165),
            .I(N__30157));
    InMux I__4150 (
            .O(N__30164),
            .I(N__30154));
    InMux I__4149 (
            .O(N__30163),
            .I(N__30151));
    Span4Mux_h I__4148 (
            .O(N__30160),
            .I(N__30148));
    LocalMux I__4147 (
            .O(N__30157),
            .I(N__30145));
    LocalMux I__4146 (
            .O(N__30154),
            .I(N__30142));
    LocalMux I__4145 (
            .O(N__30151),
            .I(encoder1_position_27));
    Odrv4 I__4144 (
            .O(N__30148),
            .I(encoder1_position_27));
    Odrv12 I__4143 (
            .O(N__30145),
            .I(encoder1_position_27));
    Odrv12 I__4142 (
            .O(N__30142),
            .I(encoder1_position_27));
    InMux I__4141 (
            .O(N__30133),
            .I(N__30130));
    LocalMux I__4140 (
            .O(N__30130),
            .I(N__30126));
    InMux I__4139 (
            .O(N__30129),
            .I(N__30123));
    Span4Mux_v I__4138 (
            .O(N__30126),
            .I(N__30120));
    LocalMux I__4137 (
            .O(N__30123),
            .I(data_out_frame_10_2));
    Odrv4 I__4136 (
            .O(N__30120),
            .I(data_out_frame_10_2));
    InMux I__4135 (
            .O(N__30115),
            .I(N__30112));
    LocalMux I__4134 (
            .O(N__30112),
            .I(N__30108));
    InMux I__4133 (
            .O(N__30111),
            .I(N__30105));
    Span4Mux_v I__4132 (
            .O(N__30108),
            .I(N__30102));
    LocalMux I__4131 (
            .O(N__30105),
            .I(data_out_frame_5_4));
    Odrv4 I__4130 (
            .O(N__30102),
            .I(data_out_frame_5_4));
    InMux I__4129 (
            .O(N__30097),
            .I(N__30094));
    LocalMux I__4128 (
            .O(N__30094),
            .I(N__30091));
    Sp12to4 I__4127 (
            .O(N__30091),
            .I(N__30088));
    Span12Mux_v I__4126 (
            .O(N__30088),
            .I(N__30085));
    Odrv12 I__4125 (
            .O(N__30085),
            .I(\c0.n11 ));
    InMux I__4124 (
            .O(N__30082),
            .I(N__30079));
    LocalMux I__4123 (
            .O(N__30079),
            .I(N__30076));
    Odrv12 I__4122 (
            .O(N__30076),
            .I(\c0.n14_adj_4329 ));
    InMux I__4121 (
            .O(N__30073),
            .I(N__30070));
    LocalMux I__4120 (
            .O(N__30070),
            .I(N__30067));
    Span4Mux_h I__4119 (
            .O(N__30067),
            .I(N__30064));
    Odrv4 I__4118 (
            .O(N__30064),
            .I(n2198));
    InMux I__4117 (
            .O(N__30061),
            .I(N__30058));
    LocalMux I__4116 (
            .O(N__30058),
            .I(N__30055));
    Span4Mux_h I__4115 (
            .O(N__30055),
            .I(N__30052));
    Odrv4 I__4114 (
            .O(N__30052),
            .I(n2192));
    InMux I__4113 (
            .O(N__30049),
            .I(N__30046));
    LocalMux I__4112 (
            .O(N__30046),
            .I(N__30043));
    Span4Mux_v I__4111 (
            .O(N__30043),
            .I(N__30040));
    Sp12to4 I__4110 (
            .O(N__30040),
            .I(N__30037));
    Odrv12 I__4109 (
            .O(N__30037),
            .I(n2186));
    InMux I__4108 (
            .O(N__30034),
            .I(N__30031));
    LocalMux I__4107 (
            .O(N__30031),
            .I(N__30026));
    CascadeMux I__4106 (
            .O(N__30030),
            .I(N__30022));
    InMux I__4105 (
            .O(N__30029),
            .I(N__30019));
    Span4Mux_v I__4104 (
            .O(N__30026),
            .I(N__30016));
    InMux I__4103 (
            .O(N__30025),
            .I(N__30011));
    InMux I__4102 (
            .O(N__30022),
            .I(N__30011));
    LocalMux I__4101 (
            .O(N__30019),
            .I(encoder1_position_19));
    Odrv4 I__4100 (
            .O(N__30016),
            .I(encoder1_position_19));
    LocalMux I__4099 (
            .O(N__30011),
            .I(encoder1_position_19));
    InMux I__4098 (
            .O(N__30004),
            .I(N__30001));
    LocalMux I__4097 (
            .O(N__30001),
            .I(\c0.n19_adj_4319 ));
    InMux I__4096 (
            .O(N__29998),
            .I(N__29995));
    LocalMux I__4095 (
            .O(N__29995),
            .I(\c0.n23557 ));
    InMux I__4094 (
            .O(N__29992),
            .I(N__29989));
    LocalMux I__4093 (
            .O(N__29989),
            .I(N__29986));
    Span4Mux_h I__4092 (
            .O(N__29986),
            .I(N__29983));
    Odrv4 I__4091 (
            .O(N__29983),
            .I(n2180));
    InMux I__4090 (
            .O(N__29980),
            .I(N__29968));
    InMux I__4089 (
            .O(N__29979),
            .I(N__29968));
    InMux I__4088 (
            .O(N__29978),
            .I(N__29968));
    InMux I__4087 (
            .O(N__29977),
            .I(N__29968));
    LocalMux I__4086 (
            .O(N__29968),
            .I(\c0.n20767 ));
    CascadeMux I__4085 (
            .O(N__29965),
            .I(\c0.n20767_cascade_ ));
    CascadeMux I__4084 (
            .O(N__29962),
            .I(N__29959));
    InMux I__4083 (
            .O(N__29959),
            .I(N__29954));
    InMux I__4082 (
            .O(N__29958),
            .I(N__29951));
    CascadeMux I__4081 (
            .O(N__29957),
            .I(N__29948));
    LocalMux I__4080 (
            .O(N__29954),
            .I(N__29944));
    LocalMux I__4079 (
            .O(N__29951),
            .I(N__29941));
    InMux I__4078 (
            .O(N__29948),
            .I(N__29938));
    InMux I__4077 (
            .O(N__29947),
            .I(N__29934));
    Span4Mux_v I__4076 (
            .O(N__29944),
            .I(N__29929));
    Span4Mux_h I__4075 (
            .O(N__29941),
            .I(N__29929));
    LocalMux I__4074 (
            .O(N__29938),
            .I(N__29926));
    InMux I__4073 (
            .O(N__29937),
            .I(N__29923));
    LocalMux I__4072 (
            .O(N__29934),
            .I(encoder1_position_24));
    Odrv4 I__4071 (
            .O(N__29929),
            .I(encoder1_position_24));
    Odrv4 I__4070 (
            .O(N__29926),
            .I(encoder1_position_24));
    LocalMux I__4069 (
            .O(N__29923),
            .I(encoder1_position_24));
    InMux I__4068 (
            .O(N__29914),
            .I(N__29911));
    LocalMux I__4067 (
            .O(N__29911),
            .I(N__29908));
    Span4Mux_h I__4066 (
            .O(N__29908),
            .I(N__29905));
    Odrv4 I__4065 (
            .O(N__29905),
            .I(n2195));
    CascadeMux I__4064 (
            .O(N__29902),
            .I(N__29899));
    InMux I__4063 (
            .O(N__29899),
            .I(N__29895));
    InMux I__4062 (
            .O(N__29898),
            .I(N__29892));
    LocalMux I__4061 (
            .O(N__29895),
            .I(data_out_frame_9_6));
    LocalMux I__4060 (
            .O(N__29892),
            .I(data_out_frame_9_6));
    InMux I__4059 (
            .O(N__29887),
            .I(N__29884));
    LocalMux I__4058 (
            .O(N__29884),
            .I(N__29880));
    InMux I__4057 (
            .O(N__29883),
            .I(N__29877));
    Span4Mux_h I__4056 (
            .O(N__29880),
            .I(N__29874));
    LocalMux I__4055 (
            .O(N__29877),
            .I(N__29869));
    Span4Mux_h I__4054 (
            .O(N__29874),
            .I(N__29869));
    Odrv4 I__4053 (
            .O(N__29869),
            .I(data_out_frame_13_6));
    InMux I__4052 (
            .O(N__29866),
            .I(N__29863));
    LocalMux I__4051 (
            .O(N__29863),
            .I(N__29860));
    Span4Mux_h I__4050 (
            .O(N__29860),
            .I(N__29857));
    Odrv4 I__4049 (
            .O(N__29857),
            .I(n2194));
    InMux I__4048 (
            .O(N__29854),
            .I(N__29847));
    InMux I__4047 (
            .O(N__29853),
            .I(N__29844));
    InMux I__4046 (
            .O(N__29852),
            .I(N__29837));
    InMux I__4045 (
            .O(N__29851),
            .I(N__29837));
    InMux I__4044 (
            .O(N__29850),
            .I(N__29837));
    LocalMux I__4043 (
            .O(N__29847),
            .I(\c0.n21175 ));
    LocalMux I__4042 (
            .O(N__29844),
            .I(\c0.n21175 ));
    LocalMux I__4041 (
            .O(N__29837),
            .I(\c0.n21175 ));
    CascadeMux I__4040 (
            .O(N__29830),
            .I(N__29826));
    InMux I__4039 (
            .O(N__29829),
            .I(N__29821));
    InMux I__4038 (
            .O(N__29826),
            .I(N__29816));
    InMux I__4037 (
            .O(N__29825),
            .I(N__29816));
    InMux I__4036 (
            .O(N__29824),
            .I(N__29813));
    LocalMux I__4035 (
            .O(N__29821),
            .I(\c0.n21156 ));
    LocalMux I__4034 (
            .O(N__29816),
            .I(\c0.n21156 ));
    LocalMux I__4033 (
            .O(N__29813),
            .I(\c0.n21156 ));
    InMux I__4032 (
            .O(N__29806),
            .I(N__29801));
    InMux I__4031 (
            .O(N__29805),
            .I(N__29796));
    InMux I__4030 (
            .O(N__29804),
            .I(N__29796));
    LocalMux I__4029 (
            .O(N__29801),
            .I(N__29791));
    LocalMux I__4028 (
            .O(N__29796),
            .I(N__29791));
    Odrv4 I__4027 (
            .O(N__29791),
            .I(\c0.n12554 ));
    InMux I__4026 (
            .O(N__29788),
            .I(N__29785));
    LocalMux I__4025 (
            .O(N__29785),
            .I(N__29782));
    Span4Mux_h I__4024 (
            .O(N__29782),
            .I(N__29777));
    InMux I__4023 (
            .O(N__29781),
            .I(N__29772));
    InMux I__4022 (
            .O(N__29780),
            .I(N__29772));
    Odrv4 I__4021 (
            .O(N__29777),
            .I(\c0.n20931 ));
    LocalMux I__4020 (
            .O(N__29772),
            .I(\c0.n20931 ));
    InMux I__4019 (
            .O(N__29767),
            .I(N__29761));
    InMux I__4018 (
            .O(N__29766),
            .I(N__29758));
    InMux I__4017 (
            .O(N__29765),
            .I(N__29753));
    InMux I__4016 (
            .O(N__29764),
            .I(N__29753));
    LocalMux I__4015 (
            .O(N__29761),
            .I(\c0.n22991 ));
    LocalMux I__4014 (
            .O(N__29758),
            .I(\c0.n22991 ));
    LocalMux I__4013 (
            .O(N__29753),
            .I(\c0.n22991 ));
    CascadeMux I__4012 (
            .O(N__29746),
            .I(\c0.n21189_cascade_ ));
    InMux I__4011 (
            .O(N__29743),
            .I(N__29739));
    InMux I__4010 (
            .O(N__29742),
            .I(N__29736));
    LocalMux I__4009 (
            .O(N__29739),
            .I(N__29733));
    LocalMux I__4008 (
            .O(N__29736),
            .I(\c0.n21058 ));
    Odrv4 I__4007 (
            .O(N__29733),
            .I(\c0.n21058 ));
    InMux I__4006 (
            .O(N__29728),
            .I(N__29722));
    InMux I__4005 (
            .O(N__29727),
            .I(N__29722));
    LocalMux I__4004 (
            .O(N__29722),
            .I(N__29718));
    InMux I__4003 (
            .O(N__29721),
            .I(N__29715));
    Odrv4 I__4002 (
            .O(N__29718),
            .I(\c0.n21192 ));
    LocalMux I__4001 (
            .O(N__29715),
            .I(\c0.n21192 ));
    InMux I__4000 (
            .O(N__29710),
            .I(N__29707));
    LocalMux I__3999 (
            .O(N__29707),
            .I(N__29702));
    InMux I__3998 (
            .O(N__29706),
            .I(N__29699));
    CascadeMux I__3997 (
            .O(N__29705),
            .I(N__29696));
    Span4Mux_v I__3996 (
            .O(N__29702),
            .I(N__29692));
    LocalMux I__3995 (
            .O(N__29699),
            .I(N__29689));
    InMux I__3994 (
            .O(N__29696),
            .I(N__29684));
    InMux I__3993 (
            .O(N__29695),
            .I(N__29684));
    Span4Mux_v I__3992 (
            .O(N__29692),
            .I(N__29679));
    Span4Mux_v I__3991 (
            .O(N__29689),
            .I(N__29679));
    LocalMux I__3990 (
            .O(N__29684),
            .I(N__29676));
    Odrv4 I__3989 (
            .O(N__29679),
            .I(\c0.n13349 ));
    Odrv12 I__3988 (
            .O(N__29676),
            .I(\c0.n13349 ));
    CascadeMux I__3987 (
            .O(N__29671),
            .I(\c0.n13480_cascade_ ));
    CascadeMux I__3986 (
            .O(N__29668),
            .I(\c0.n21122_cascade_ ));
    CascadeMux I__3985 (
            .O(N__29665),
            .I(N__29661));
    InMux I__3984 (
            .O(N__29664),
            .I(N__29656));
    InMux I__3983 (
            .O(N__29661),
            .I(N__29652));
    InMux I__3982 (
            .O(N__29660),
            .I(N__29647));
    InMux I__3981 (
            .O(N__29659),
            .I(N__29647));
    LocalMux I__3980 (
            .O(N__29656),
            .I(N__29644));
    InMux I__3979 (
            .O(N__29655),
            .I(N__29641));
    LocalMux I__3978 (
            .O(N__29652),
            .I(N__29636));
    LocalMux I__3977 (
            .O(N__29647),
            .I(N__29631));
    Span4Mux_v I__3976 (
            .O(N__29644),
            .I(N__29631));
    LocalMux I__3975 (
            .O(N__29641),
            .I(N__29628));
    InMux I__3974 (
            .O(N__29640),
            .I(N__29623));
    InMux I__3973 (
            .O(N__29639),
            .I(N__29623));
    Span4Mux_v I__3972 (
            .O(N__29636),
            .I(N__29618));
    Span4Mux_h I__3971 (
            .O(N__29631),
            .I(N__29618));
    Odrv4 I__3970 (
            .O(N__29628),
            .I(encoder1_position_14));
    LocalMux I__3969 (
            .O(N__29623),
            .I(encoder1_position_14));
    Odrv4 I__3968 (
            .O(N__29618),
            .I(encoder1_position_14));
    CascadeMux I__3967 (
            .O(N__29611),
            .I(\c0.n6_adj_4509_cascade_ ));
    InMux I__3966 (
            .O(N__29608),
            .I(N__29605));
    LocalMux I__3965 (
            .O(N__29605),
            .I(\c0.n22393 ));
    InMux I__3964 (
            .O(N__29602),
            .I(N__29597));
    InMux I__3963 (
            .O(N__29601),
            .I(N__29594));
    InMux I__3962 (
            .O(N__29600),
            .I(N__29591));
    LocalMux I__3961 (
            .O(N__29597),
            .I(\c0.n10498 ));
    LocalMux I__3960 (
            .O(N__29594),
            .I(\c0.n10498 ));
    LocalMux I__3959 (
            .O(N__29591),
            .I(\c0.n10498 ));
    CascadeMux I__3958 (
            .O(N__29584),
            .I(\c0.n22393_cascade_ ));
    CascadeMux I__3957 (
            .O(N__29581),
            .I(\c0.n14_adj_4510_cascade_ ));
    InMux I__3956 (
            .O(N__29578),
            .I(N__29570));
    InMux I__3955 (
            .O(N__29577),
            .I(N__29570));
    InMux I__3954 (
            .O(N__29576),
            .I(N__29565));
    InMux I__3953 (
            .O(N__29575),
            .I(N__29565));
    LocalMux I__3952 (
            .O(N__29570),
            .I(N__29559));
    LocalMux I__3951 (
            .O(N__29565),
            .I(N__29556));
    InMux I__3950 (
            .O(N__29564),
            .I(N__29553));
    InMux I__3949 (
            .O(N__29563),
            .I(N__29550));
    InMux I__3948 (
            .O(N__29562),
            .I(N__29547));
    Span4Mux_h I__3947 (
            .O(N__29559),
            .I(N__29544));
    Span4Mux_h I__3946 (
            .O(N__29556),
            .I(N__29537));
    LocalMux I__3945 (
            .O(N__29553),
            .I(N__29537));
    LocalMux I__3944 (
            .O(N__29550),
            .I(N__29537));
    LocalMux I__3943 (
            .O(N__29547),
            .I(\c0.n10462 ));
    Odrv4 I__3942 (
            .O(N__29544),
            .I(\c0.n10462 ));
    Odrv4 I__3941 (
            .O(N__29537),
            .I(\c0.n10462 ));
    InMux I__3940 (
            .O(N__29530),
            .I(N__29524));
    InMux I__3939 (
            .O(N__29529),
            .I(N__29524));
    LocalMux I__3938 (
            .O(N__29524),
            .I(N__29521));
    Span4Mux_h I__3937 (
            .O(N__29521),
            .I(N__29517));
    InMux I__3936 (
            .O(N__29520),
            .I(N__29514));
    Odrv4 I__3935 (
            .O(N__29517),
            .I(\c0.n21150 ));
    LocalMux I__3934 (
            .O(N__29514),
            .I(\c0.n21150 ));
    InMux I__3933 (
            .O(N__29509),
            .I(N__29506));
    LocalMux I__3932 (
            .O(N__29506),
            .I(\c0.n10_adj_4511 ));
    InMux I__3931 (
            .O(N__29503),
            .I(N__29500));
    LocalMux I__3930 (
            .O(N__29500),
            .I(\c0.n10_adj_4330 ));
    CascadeMux I__3929 (
            .O(N__29497),
            .I(\c0.n21192_cascade_ ));
    CascadeMux I__3928 (
            .O(N__29494),
            .I(\c0.n20931_cascade_ ));
    InMux I__3927 (
            .O(N__29491),
            .I(N__29488));
    LocalMux I__3926 (
            .O(N__29488),
            .I(\c0.n22151 ));
    CascadeMux I__3925 (
            .O(N__29485),
            .I(\c0.n22151_cascade_ ));
    CascadeMux I__3924 (
            .O(N__29482),
            .I(\c0.n6_adj_4397_cascade_ ));
    InMux I__3923 (
            .O(N__29479),
            .I(N__29476));
    LocalMux I__3922 (
            .O(N__29476),
            .I(\c0.data_out_frame_28_0 ));
    CascadeMux I__3921 (
            .O(N__29473),
            .I(N__29470));
    InMux I__3920 (
            .O(N__29470),
            .I(N__29467));
    LocalMux I__3919 (
            .O(N__29467),
            .I(N__29463));
    InMux I__3918 (
            .O(N__29466),
            .I(N__29460));
    Odrv4 I__3917 (
            .O(N__29463),
            .I(\c0.n22018 ));
    LocalMux I__3916 (
            .O(N__29460),
            .I(\c0.n22018 ));
    InMux I__3915 (
            .O(N__29455),
            .I(N__29452));
    LocalMux I__3914 (
            .O(N__29452),
            .I(\c0.data_out_frame_29_5 ));
    InMux I__3913 (
            .O(N__29449),
            .I(N__29446));
    LocalMux I__3912 (
            .O(N__29446),
            .I(\c0.data_out_frame_28_5 ));
    InMux I__3911 (
            .O(N__29443),
            .I(N__29440));
    LocalMux I__3910 (
            .O(N__29440),
            .I(N__29437));
    Span4Mux_h I__3909 (
            .O(N__29437),
            .I(N__29434));
    Sp12to4 I__3908 (
            .O(N__29434),
            .I(N__29431));
    Span12Mux_v I__3907 (
            .O(N__29431),
            .I(N__29428));
    Odrv12 I__3906 (
            .O(N__29428),
            .I(\c0.n26_adj_4347 ));
    InMux I__3905 (
            .O(N__29425),
            .I(N__29420));
    InMux I__3904 (
            .O(N__29424),
            .I(N__29417));
    InMux I__3903 (
            .O(N__29423),
            .I(N__29413));
    LocalMux I__3902 (
            .O(N__29420),
            .I(N__29408));
    LocalMux I__3901 (
            .O(N__29417),
            .I(N__29405));
    InMux I__3900 (
            .O(N__29416),
            .I(N__29402));
    LocalMux I__3899 (
            .O(N__29413),
            .I(N__29399));
    InMux I__3898 (
            .O(N__29412),
            .I(N__29394));
    InMux I__3897 (
            .O(N__29411),
            .I(N__29394));
    Span4Mux_v I__3896 (
            .O(N__29408),
            .I(N__29389));
    Span4Mux_v I__3895 (
            .O(N__29405),
            .I(N__29389));
    LocalMux I__3894 (
            .O(N__29402),
            .I(\c0.n20376 ));
    Odrv4 I__3893 (
            .O(N__29399),
            .I(\c0.n20376 ));
    LocalMux I__3892 (
            .O(N__29394),
            .I(\c0.n20376 ));
    Odrv4 I__3891 (
            .O(N__29389),
            .I(\c0.n20376 ));
    CascadeMux I__3890 (
            .O(N__29380),
            .I(\c0.n22018_cascade_ ));
    CascadeMux I__3889 (
            .O(N__29377),
            .I(N__29374));
    InMux I__3888 (
            .O(N__29374),
            .I(N__29371));
    LocalMux I__3887 (
            .O(N__29371),
            .I(N__29368));
    Span4Mux_h I__3886 (
            .O(N__29368),
            .I(N__29365));
    Odrv4 I__3885 (
            .O(N__29365),
            .I(\c0.n21946 ));
    CascadeMux I__3884 (
            .O(N__29362),
            .I(\c0.n21946_cascade_ ));
    InMux I__3883 (
            .O(N__29359),
            .I(N__29355));
    InMux I__3882 (
            .O(N__29358),
            .I(N__29350));
    LocalMux I__3881 (
            .O(N__29355),
            .I(N__29347));
    InMux I__3880 (
            .O(N__29354),
            .I(N__29344));
    InMux I__3879 (
            .O(N__29353),
            .I(N__29341));
    LocalMux I__3878 (
            .O(N__29350),
            .I(N__29338));
    Span4Mux_h I__3877 (
            .O(N__29347),
            .I(N__29335));
    LocalMux I__3876 (
            .O(N__29344),
            .I(N__29332));
    LocalMux I__3875 (
            .O(N__29341),
            .I(N__29327));
    Span4Mux_h I__3874 (
            .O(N__29338),
            .I(N__29327));
    Odrv4 I__3873 (
            .O(N__29335),
            .I(\c0.n12532 ));
    Odrv4 I__3872 (
            .O(N__29332),
            .I(\c0.n12532 ));
    Odrv4 I__3871 (
            .O(N__29327),
            .I(\c0.n12532 ));
    CascadeMux I__3870 (
            .O(N__29320),
            .I(\c0.n12491_cascade_ ));
    InMux I__3869 (
            .O(N__29317),
            .I(N__29314));
    LocalMux I__3868 (
            .O(N__29314),
            .I(\c0.data_out_frame_28_6 ));
    InMux I__3867 (
            .O(N__29311),
            .I(N__29308));
    LocalMux I__3866 (
            .O(N__29308),
            .I(N__29305));
    Span4Mux_v I__3865 (
            .O(N__29305),
            .I(N__29302));
    Span4Mux_v I__3864 (
            .O(N__29302),
            .I(N__29299));
    Odrv4 I__3863 (
            .O(N__29299),
            .I(\c0.n26_adj_4351 ));
    CascadeMux I__3862 (
            .O(N__29296),
            .I(\c0.n7_adj_4307_cascade_ ));
    InMux I__3861 (
            .O(N__29293),
            .I(N__29289));
    InMux I__3860 (
            .O(N__29292),
            .I(N__29286));
    LocalMux I__3859 (
            .O(N__29289),
            .I(N__29283));
    LocalMux I__3858 (
            .O(N__29286),
            .I(N__29280));
    Span4Mux_h I__3857 (
            .O(N__29283),
            .I(N__29277));
    Odrv4 I__3856 (
            .O(N__29280),
            .I(data_out_frame_29__3__N_1662));
    Odrv4 I__3855 (
            .O(N__29277),
            .I(data_out_frame_29__3__N_1662));
    InMux I__3854 (
            .O(N__29272),
            .I(N__29267));
    InMux I__3853 (
            .O(N__29271),
            .I(N__29264));
    InMux I__3852 (
            .O(N__29270),
            .I(N__29261));
    LocalMux I__3851 (
            .O(N__29267),
            .I(\c0.n22024 ));
    LocalMux I__3850 (
            .O(N__29264),
            .I(\c0.n22024 ));
    LocalMux I__3849 (
            .O(N__29261),
            .I(\c0.n22024 ));
    InMux I__3848 (
            .O(N__29254),
            .I(N__29251));
    LocalMux I__3847 (
            .O(N__29251),
            .I(N__29248));
    Odrv12 I__3846 (
            .O(N__29248),
            .I(\c0.data_out_frame_29_4 ));
    SRMux I__3845 (
            .O(N__29245),
            .I(N__29242));
    LocalMux I__3844 (
            .O(N__29242),
            .I(N__29239));
    Span4Mux_h I__3843 (
            .O(N__29239),
            .I(N__29236));
    Odrv4 I__3842 (
            .O(N__29236),
            .I(\c0.n21376 ));
    SRMux I__3841 (
            .O(N__29233),
            .I(N__29230));
    LocalMux I__3840 (
            .O(N__29230),
            .I(\c0.n21362 ));
    CascadeMux I__3839 (
            .O(N__29227),
            .I(N__29224));
    InMux I__3838 (
            .O(N__29224),
            .I(N__29221));
    LocalMux I__3837 (
            .O(N__29221),
            .I(N__29218));
    Odrv4 I__3836 (
            .O(N__29218),
            .I(\c0.n21128 ));
    InMux I__3835 (
            .O(N__29215),
            .I(N__29212));
    LocalMux I__3834 (
            .O(N__29212),
            .I(\c0.n12_adj_4516 ));
    InMux I__3833 (
            .O(N__29209),
            .I(N__29206));
    LocalMux I__3832 (
            .O(N__29206),
            .I(\c0.n9_adj_4339 ));
    CascadeMux I__3831 (
            .O(N__29203),
            .I(\c0.tx.n16631_cascade_ ));
    InMux I__3830 (
            .O(N__29200),
            .I(N__29194));
    InMux I__3829 (
            .O(N__29199),
            .I(N__29194));
    LocalMux I__3828 (
            .O(N__29194),
            .I(N__29189));
    InMux I__3827 (
            .O(N__29193),
            .I(N__29186));
    InMux I__3826 (
            .O(N__29192),
            .I(N__29183));
    Span4Mux_h I__3825 (
            .O(N__29189),
            .I(N__29180));
    LocalMux I__3824 (
            .O(N__29186),
            .I(n14442));
    LocalMux I__3823 (
            .O(N__29183),
            .I(n14442));
    Odrv4 I__3822 (
            .O(N__29180),
            .I(n14442));
    SRMux I__3821 (
            .O(N__29173),
            .I(N__29170));
    LocalMux I__3820 (
            .O(N__29170),
            .I(N__29167));
    Odrv4 I__3819 (
            .O(N__29167),
            .I(\c0.n21370 ));
    CascadeMux I__3818 (
            .O(N__29164),
            .I(\c0.n10_adj_4231_cascade_ ));
    InMux I__3817 (
            .O(N__29161),
            .I(N__29158));
    LocalMux I__3816 (
            .O(N__29158),
            .I(\c0.n14 ));
    InMux I__3815 (
            .O(N__29155),
            .I(N__29149));
    InMux I__3814 (
            .O(N__29154),
            .I(N__29146));
    InMux I__3813 (
            .O(N__29153),
            .I(N__29139));
    InMux I__3812 (
            .O(N__29152),
            .I(N__29139));
    LocalMux I__3811 (
            .O(N__29149),
            .I(N__29136));
    LocalMux I__3810 (
            .O(N__29146),
            .I(N__29132));
    InMux I__3809 (
            .O(N__29145),
            .I(N__29127));
    InMux I__3808 (
            .O(N__29144),
            .I(N__29127));
    LocalMux I__3807 (
            .O(N__29139),
            .I(N__29124));
    Span4Mux_v I__3806 (
            .O(N__29136),
            .I(N__29121));
    InMux I__3805 (
            .O(N__29135),
            .I(N__29118));
    Span12Mux_s11_h I__3804 (
            .O(N__29132),
            .I(N__29114));
    LocalMux I__3803 (
            .O(N__29127),
            .I(N__29111));
    Span4Mux_h I__3802 (
            .O(N__29124),
            .I(N__29108));
    Span4Mux_v I__3801 (
            .O(N__29121),
            .I(N__29103));
    LocalMux I__3800 (
            .O(N__29118),
            .I(N__29103));
    InMux I__3799 (
            .O(N__29117),
            .I(N__29100));
    Odrv12 I__3798 (
            .O(N__29114),
            .I(n9539));
    Odrv12 I__3797 (
            .O(N__29111),
            .I(n9539));
    Odrv4 I__3796 (
            .O(N__29108),
            .I(n9539));
    Odrv4 I__3795 (
            .O(N__29103),
            .I(n9539));
    LocalMux I__3794 (
            .O(N__29100),
            .I(n9539));
    CascadeMux I__3793 (
            .O(N__29089),
            .I(N__29085));
    InMux I__3792 (
            .O(N__29088),
            .I(N__29082));
    InMux I__3791 (
            .O(N__29085),
            .I(N__29079));
    LocalMux I__3790 (
            .O(N__29082),
            .I(data_out_frame_10_0));
    LocalMux I__3789 (
            .O(N__29079),
            .I(data_out_frame_10_0));
    InMux I__3788 (
            .O(N__29074),
            .I(N__29071));
    LocalMux I__3787 (
            .O(N__29071),
            .I(N__29065));
    InMux I__3786 (
            .O(N__29070),
            .I(N__29062));
    InMux I__3785 (
            .O(N__29069),
            .I(N__29057));
    InMux I__3784 (
            .O(N__29068),
            .I(N__29057));
    Odrv4 I__3783 (
            .O(N__29065),
            .I(data_in_3_3));
    LocalMux I__3782 (
            .O(N__29062),
            .I(data_in_3_3));
    LocalMux I__3781 (
            .O(N__29057),
            .I(data_in_3_3));
    CascadeMux I__3780 (
            .O(N__29050),
            .I(N__29046));
    CascadeMux I__3779 (
            .O(N__29049),
            .I(N__29043));
    InMux I__3778 (
            .O(N__29046),
            .I(N__29039));
    InMux I__3777 (
            .O(N__29043),
            .I(N__29036));
    InMux I__3776 (
            .O(N__29042),
            .I(N__29033));
    LocalMux I__3775 (
            .O(N__29039),
            .I(N__29029));
    LocalMux I__3774 (
            .O(N__29036),
            .I(N__29024));
    LocalMux I__3773 (
            .O(N__29033),
            .I(N__29024));
    InMux I__3772 (
            .O(N__29032),
            .I(N__29021));
    Span4Mux_h I__3771 (
            .O(N__29029),
            .I(N__29016));
    Span4Mux_h I__3770 (
            .O(N__29024),
            .I(N__29016));
    LocalMux I__3769 (
            .O(N__29021),
            .I(encoder1_position_18));
    Odrv4 I__3768 (
            .O(N__29016),
            .I(encoder1_position_18));
    CascadeMux I__3767 (
            .O(N__29011),
            .I(N__29007));
    InMux I__3766 (
            .O(N__29010),
            .I(N__29004));
    InMux I__3765 (
            .O(N__29007),
            .I(N__29001));
    LocalMux I__3764 (
            .O(N__29004),
            .I(data_out_frame_11_2));
    LocalMux I__3763 (
            .O(N__29001),
            .I(data_out_frame_11_2));
    InMux I__3762 (
            .O(N__28996),
            .I(N__28993));
    LocalMux I__3761 (
            .O(N__28993),
            .I(N__28990));
    Span4Mux_v I__3760 (
            .O(N__28990),
            .I(N__28987));
    Odrv4 I__3759 (
            .O(N__28987),
            .I(\c0.n24177 ));
    InMux I__3758 (
            .O(N__28984),
            .I(N__28980));
    InMux I__3757 (
            .O(N__28983),
            .I(N__28977));
    LocalMux I__3756 (
            .O(N__28980),
            .I(N__28974));
    LocalMux I__3755 (
            .O(N__28977),
            .I(N__28969));
    Span4Mux_h I__3754 (
            .O(N__28974),
            .I(N__28969));
    Odrv4 I__3753 (
            .O(N__28969),
            .I(data_out_frame_5_0));
    InMux I__3752 (
            .O(N__28966),
            .I(N__28962));
    CascadeMux I__3751 (
            .O(N__28965),
            .I(N__28959));
    LocalMux I__3750 (
            .O(N__28962),
            .I(N__28955));
    InMux I__3749 (
            .O(N__28959),
            .I(N__28951));
    InMux I__3748 (
            .O(N__28958),
            .I(N__28948));
    Span4Mux_v I__3747 (
            .O(N__28955),
            .I(N__28945));
    InMux I__3746 (
            .O(N__28954),
            .I(N__28942));
    LocalMux I__3745 (
            .O(N__28951),
            .I(N__28939));
    LocalMux I__3744 (
            .O(N__28948),
            .I(encoder1_position_29));
    Odrv4 I__3743 (
            .O(N__28945),
            .I(encoder1_position_29));
    LocalMux I__3742 (
            .O(N__28942),
            .I(encoder1_position_29));
    Odrv12 I__3741 (
            .O(N__28939),
            .I(encoder1_position_29));
    CascadeMux I__3740 (
            .O(N__28930),
            .I(N__28926));
    InMux I__3739 (
            .O(N__28929),
            .I(N__28923));
    InMux I__3738 (
            .O(N__28926),
            .I(N__28920));
    LocalMux I__3737 (
            .O(N__28923),
            .I(N__28917));
    LocalMux I__3736 (
            .O(N__28920),
            .I(data_out_frame_10_5));
    Odrv4 I__3735 (
            .O(N__28917),
            .I(data_out_frame_10_5));
    InMux I__3734 (
            .O(N__28912),
            .I(N__28908));
    InMux I__3733 (
            .O(N__28911),
            .I(N__28905));
    LocalMux I__3732 (
            .O(N__28908),
            .I(data_out_frame_12_3));
    LocalMux I__3731 (
            .O(N__28905),
            .I(data_out_frame_12_3));
    CascadeMux I__3730 (
            .O(N__28900),
            .I(\c0.n7_adj_4492_cascade_ ));
    CascadeMux I__3729 (
            .O(N__28897),
            .I(N__28893));
    InMux I__3728 (
            .O(N__28896),
            .I(N__28890));
    InMux I__3727 (
            .O(N__28893),
            .I(N__28885));
    LocalMux I__3726 (
            .O(N__28890),
            .I(N__28882));
    InMux I__3725 (
            .O(N__28889),
            .I(N__28877));
    InMux I__3724 (
            .O(N__28888),
            .I(N__28877));
    LocalMux I__3723 (
            .O(N__28885),
            .I(data_in_1_5));
    Odrv4 I__3722 (
            .O(N__28882),
            .I(data_in_1_5));
    LocalMux I__3721 (
            .O(N__28877),
            .I(data_in_1_5));
    InMux I__3720 (
            .O(N__28870),
            .I(N__28867));
    LocalMux I__3719 (
            .O(N__28867),
            .I(\c0.n9_adj_4493 ));
    InMux I__3718 (
            .O(N__28864),
            .I(N__28861));
    LocalMux I__3717 (
            .O(N__28861),
            .I(\c0.n23600 ));
    InMux I__3716 (
            .O(N__28858),
            .I(N__28849));
    InMux I__3715 (
            .O(N__28857),
            .I(N__28849));
    InMux I__3714 (
            .O(N__28856),
            .I(N__28849));
    LocalMux I__3713 (
            .O(N__28849),
            .I(data_in_0_6));
    InMux I__3712 (
            .O(N__28846),
            .I(N__28840));
    InMux I__3711 (
            .O(N__28845),
            .I(N__28837));
    InMux I__3710 (
            .O(N__28844),
            .I(N__28832));
    InMux I__3709 (
            .O(N__28843),
            .I(N__28832));
    LocalMux I__3708 (
            .O(N__28840),
            .I(N__28825));
    LocalMux I__3707 (
            .O(N__28837),
            .I(N__28825));
    LocalMux I__3706 (
            .O(N__28832),
            .I(N__28825));
    Odrv4 I__3705 (
            .O(N__28825),
            .I(data_in_2_2));
    CascadeMux I__3704 (
            .O(N__28822),
            .I(N__28819));
    InMux I__3703 (
            .O(N__28819),
            .I(N__28815));
    InMux I__3702 (
            .O(N__28818),
            .I(N__28812));
    LocalMux I__3701 (
            .O(N__28815),
            .I(N__28806));
    LocalMux I__3700 (
            .O(N__28812),
            .I(N__28806));
    InMux I__3699 (
            .O(N__28811),
            .I(N__28803));
    Span4Mux_v I__3698 (
            .O(N__28806),
            .I(N__28800));
    LocalMux I__3697 (
            .O(N__28803),
            .I(data_in_0_3));
    Odrv4 I__3696 (
            .O(N__28800),
            .I(data_in_0_3));
    CascadeMux I__3695 (
            .O(N__28795),
            .I(\c0.n14_adj_4495_cascade_ ));
    InMux I__3694 (
            .O(N__28792),
            .I(N__28789));
    LocalMux I__3693 (
            .O(N__28789),
            .I(\c0.n15_adj_4496 ));
    CascadeMux I__3692 (
            .O(N__28786),
            .I(N__28783));
    InMux I__3691 (
            .O(N__28783),
            .I(N__28778));
    InMux I__3690 (
            .O(N__28782),
            .I(N__28775));
    InMux I__3689 (
            .O(N__28781),
            .I(N__28772));
    LocalMux I__3688 (
            .O(N__28778),
            .I(N__28767));
    LocalMux I__3687 (
            .O(N__28775),
            .I(N__28762));
    LocalMux I__3686 (
            .O(N__28772),
            .I(N__28762));
    InMux I__3685 (
            .O(N__28771),
            .I(N__28759));
    InMux I__3684 (
            .O(N__28770),
            .I(N__28756));
    Span4Mux_h I__3683 (
            .O(N__28767),
            .I(N__28753));
    Span4Mux_v I__3682 (
            .O(N__28762),
            .I(N__28750));
    LocalMux I__3681 (
            .O(N__28759),
            .I(encoder1_position_31));
    LocalMux I__3680 (
            .O(N__28756),
            .I(encoder1_position_31));
    Odrv4 I__3679 (
            .O(N__28753),
            .I(encoder1_position_31));
    Odrv4 I__3678 (
            .O(N__28750),
            .I(encoder1_position_31));
    CascadeMux I__3677 (
            .O(N__28741),
            .I(N__28737));
    InMux I__3676 (
            .O(N__28740),
            .I(N__28734));
    InMux I__3675 (
            .O(N__28737),
            .I(N__28731));
    LocalMux I__3674 (
            .O(N__28734),
            .I(N__28728));
    LocalMux I__3673 (
            .O(N__28731),
            .I(data_out_frame_10_7));
    Odrv4 I__3672 (
            .O(N__28728),
            .I(data_out_frame_10_7));
    InMux I__3671 (
            .O(N__28723),
            .I(N__28719));
    InMux I__3670 (
            .O(N__28722),
            .I(N__28716));
    LocalMux I__3669 (
            .O(N__28719),
            .I(N__28713));
    LocalMux I__3668 (
            .O(N__28716),
            .I(data_out_frame_8_7));
    Odrv4 I__3667 (
            .O(N__28713),
            .I(data_out_frame_8_7));
    InMux I__3666 (
            .O(N__28708),
            .I(N__28705));
    LocalMux I__3665 (
            .O(N__28705),
            .I(N__28701));
    InMux I__3664 (
            .O(N__28704),
            .I(N__28698));
    Span4Mux_v I__3663 (
            .O(N__28701),
            .I(N__28695));
    LocalMux I__3662 (
            .O(N__28698),
            .I(data_out_frame_11_7));
    Odrv4 I__3661 (
            .O(N__28695),
            .I(data_out_frame_11_7));
    InMux I__3660 (
            .O(N__28690),
            .I(N__28687));
    LocalMux I__3659 (
            .O(N__28687),
            .I(N__28684));
    Span4Mux_v I__3658 (
            .O(N__28684),
            .I(N__28681));
    Odrv4 I__3657 (
            .O(N__28681),
            .I(n2181));
    InMux I__3656 (
            .O(N__28678),
            .I(N__28675));
    LocalMux I__3655 (
            .O(N__28675),
            .I(N__28672));
    Span4Mux_h I__3654 (
            .O(N__28672),
            .I(N__28669));
    Odrv4 I__3653 (
            .O(N__28669),
            .I(\c0.n22224 ));
    CascadeMux I__3652 (
            .O(N__28666),
            .I(\c0.n22224_cascade_ ));
    CascadeMux I__3651 (
            .O(N__28663),
            .I(\c0.n13349_cascade_ ));
    InMux I__3650 (
            .O(N__28660),
            .I(N__28657));
    LocalMux I__3649 (
            .O(N__28657),
            .I(N__28654));
    Odrv4 I__3648 (
            .O(N__28654),
            .I(\c0.n6_adj_4334 ));
    InMux I__3647 (
            .O(N__28651),
            .I(N__28648));
    LocalMux I__3646 (
            .O(N__28648),
            .I(N__28645));
    Span4Mux_h I__3645 (
            .O(N__28645),
            .I(N__28642));
    Odrv4 I__3644 (
            .O(N__28642),
            .I(n24104));
    InMux I__3643 (
            .O(N__28639),
            .I(N__28636));
    LocalMux I__3642 (
            .O(N__28636),
            .I(\c0.n22405 ));
    InMux I__3641 (
            .O(N__28633),
            .I(N__28630));
    LocalMux I__3640 (
            .O(N__28630),
            .I(\c0.n22102 ));
    CascadeMux I__3639 (
            .O(N__28627),
            .I(\c0.n22361_cascade_ ));
    InMux I__3638 (
            .O(N__28624),
            .I(N__28621));
    LocalMux I__3637 (
            .O(N__28621),
            .I(N__28618));
    Odrv4 I__3636 (
            .O(N__28618),
            .I(\c0.n10_adj_4314 ));
    CascadeMux I__3635 (
            .O(N__28615),
            .I(N__28612));
    InMux I__3634 (
            .O(N__28612),
            .I(N__28607));
    InMux I__3633 (
            .O(N__28611),
            .I(N__28603));
    InMux I__3632 (
            .O(N__28610),
            .I(N__28600));
    LocalMux I__3631 (
            .O(N__28607),
            .I(N__28597));
    InMux I__3630 (
            .O(N__28606),
            .I(N__28594));
    LocalMux I__3629 (
            .O(N__28603),
            .I(N__28591));
    LocalMux I__3628 (
            .O(N__28600),
            .I(encoder1_position_21));
    Odrv12 I__3627 (
            .O(N__28597),
            .I(encoder1_position_21));
    LocalMux I__3626 (
            .O(N__28594),
            .I(encoder1_position_21));
    Odrv4 I__3625 (
            .O(N__28591),
            .I(encoder1_position_21));
    InMux I__3624 (
            .O(N__28582),
            .I(N__28579));
    LocalMux I__3623 (
            .O(N__28579),
            .I(N__28576));
    Span4Mux_v I__3622 (
            .O(N__28576),
            .I(N__28573));
    Span4Mux_h I__3621 (
            .O(N__28573),
            .I(N__28570));
    Odrv4 I__3620 (
            .O(N__28570),
            .I(\c0.n24153 ));
    CascadeMux I__3619 (
            .O(N__28567),
            .I(N__28563));
    InMux I__3618 (
            .O(N__28566),
            .I(N__28558));
    InMux I__3617 (
            .O(N__28563),
            .I(N__28558));
    LocalMux I__3616 (
            .O(N__28558),
            .I(data_out_frame_8_6));
    InMux I__3615 (
            .O(N__28555),
            .I(N__28552));
    LocalMux I__3614 (
            .O(N__28552),
            .I(N__28549));
    Span4Mux_h I__3613 (
            .O(N__28549),
            .I(N__28546));
    Odrv4 I__3612 (
            .O(N__28546),
            .I(\c0.n24156 ));
    InMux I__3611 (
            .O(N__28543),
            .I(N__28540));
    LocalMux I__3610 (
            .O(N__28540),
            .I(N__28536));
    InMux I__3609 (
            .O(N__28539),
            .I(N__28533));
    Span4Mux_h I__3608 (
            .O(N__28536),
            .I(N__28530));
    LocalMux I__3607 (
            .O(N__28533),
            .I(data_out_frame_12_6));
    Odrv4 I__3606 (
            .O(N__28530),
            .I(data_out_frame_12_6));
    CascadeMux I__3605 (
            .O(N__28525),
            .I(N__28522));
    InMux I__3604 (
            .O(N__28522),
            .I(N__28518));
    CascadeMux I__3603 (
            .O(N__28521),
            .I(N__28515));
    LocalMux I__3602 (
            .O(N__28518),
            .I(N__28512));
    InMux I__3601 (
            .O(N__28515),
            .I(N__28509));
    Span4Mux_v I__3600 (
            .O(N__28512),
            .I(N__28506));
    LocalMux I__3599 (
            .O(N__28509),
            .I(data_out_frame_11_3));
    Odrv4 I__3598 (
            .O(N__28506),
            .I(data_out_frame_11_3));
    CascadeMux I__3597 (
            .O(N__28501),
            .I(\c0.n21110_cascade_ ));
    InMux I__3596 (
            .O(N__28498),
            .I(N__28495));
    LocalMux I__3595 (
            .O(N__28495),
            .I(N__28492));
    Odrv12 I__3594 (
            .O(N__28492),
            .I(\c0.n14_adj_4514 ));
    InMux I__3593 (
            .O(N__28489),
            .I(N__28482));
    InMux I__3592 (
            .O(N__28488),
            .I(N__28482));
    CascadeMux I__3591 (
            .O(N__28487),
            .I(N__28478));
    LocalMux I__3590 (
            .O(N__28482),
            .I(N__28475));
    InMux I__3589 (
            .O(N__28481),
            .I(N__28471));
    InMux I__3588 (
            .O(N__28478),
            .I(N__28467));
    Span4Mux_v I__3587 (
            .O(N__28475),
            .I(N__28464));
    InMux I__3586 (
            .O(N__28474),
            .I(N__28461));
    LocalMux I__3585 (
            .O(N__28471),
            .I(N__28458));
    InMux I__3584 (
            .O(N__28470),
            .I(N__28455));
    LocalMux I__3583 (
            .O(N__28467),
            .I(N__28452));
    Span4Mux_h I__3582 (
            .O(N__28464),
            .I(N__28447));
    LocalMux I__3581 (
            .O(N__28461),
            .I(N__28447));
    Odrv4 I__3580 (
            .O(N__28458),
            .I(encoder1_position_22));
    LocalMux I__3579 (
            .O(N__28455),
            .I(encoder1_position_22));
    Odrv4 I__3578 (
            .O(N__28452),
            .I(encoder1_position_22));
    Odrv4 I__3577 (
            .O(N__28447),
            .I(encoder1_position_22));
    InMux I__3576 (
            .O(N__28438),
            .I(N__28435));
    LocalMux I__3575 (
            .O(N__28435),
            .I(N__28432));
    Span4Mux_h I__3574 (
            .O(N__28432),
            .I(N__28429));
    Odrv4 I__3573 (
            .O(N__28429),
            .I(n2201));
    InMux I__3572 (
            .O(N__28426),
            .I(N__28423));
    LocalMux I__3571 (
            .O(N__28423),
            .I(N__28419));
    InMux I__3570 (
            .O(N__28422),
            .I(N__28416));
    Span4Mux_h I__3569 (
            .O(N__28419),
            .I(N__28413));
    LocalMux I__3568 (
            .O(N__28416),
            .I(N__28410));
    Odrv4 I__3567 (
            .O(N__28413),
            .I(\c0.n22277 ));
    Odrv12 I__3566 (
            .O(N__28410),
            .I(\c0.n22277 ));
    CascadeMux I__3565 (
            .O(N__28405),
            .I(\c0.n22102_cascade_ ));
    InMux I__3564 (
            .O(N__28402),
            .I(N__28399));
    LocalMux I__3563 (
            .O(N__28399),
            .I(\c0.n22293 ));
    CascadeMux I__3562 (
            .O(N__28396),
            .I(\c0.n15_adj_4325_cascade_ ));
    InMux I__3561 (
            .O(N__28393),
            .I(N__28384));
    InMux I__3560 (
            .O(N__28392),
            .I(N__28384));
    InMux I__3559 (
            .O(N__28391),
            .I(N__28384));
    LocalMux I__3558 (
            .O(N__28384),
            .I(N__28381));
    Odrv4 I__3557 (
            .O(N__28381),
            .I(\c0.n21041 ));
    CascadeMux I__3556 (
            .O(N__28378),
            .I(\c0.n21041_cascade_ ));
    CascadeMux I__3555 (
            .O(N__28375),
            .I(\c0.n6_adj_4313_cascade_ ));
    CascadeMux I__3554 (
            .O(N__28372),
            .I(\c0.n21156_cascade_ ));
    CascadeMux I__3553 (
            .O(N__28369),
            .I(\c0.n21175_cascade_ ));
    CascadeMux I__3552 (
            .O(N__28366),
            .I(\c0.n20276_cascade_ ));
    InMux I__3551 (
            .O(N__28363),
            .I(N__28360));
    LocalMux I__3550 (
            .O(N__28360),
            .I(\c0.n22066 ));
    CascadeMux I__3549 (
            .O(N__28357),
            .I(N__28353));
    CascadeMux I__3548 (
            .O(N__28356),
            .I(N__28349));
    InMux I__3547 (
            .O(N__28353),
            .I(N__28346));
    InMux I__3546 (
            .O(N__28352),
            .I(N__28339));
    InMux I__3545 (
            .O(N__28349),
            .I(N__28339));
    LocalMux I__3544 (
            .O(N__28346),
            .I(N__28335));
    InMux I__3543 (
            .O(N__28345),
            .I(N__28329));
    InMux I__3542 (
            .O(N__28344),
            .I(N__28329));
    LocalMux I__3541 (
            .O(N__28339),
            .I(N__28326));
    InMux I__3540 (
            .O(N__28338),
            .I(N__28322));
    Span4Mux_h I__3539 (
            .O(N__28335),
            .I(N__28318));
    InMux I__3538 (
            .O(N__28334),
            .I(N__28315));
    LocalMux I__3537 (
            .O(N__28329),
            .I(N__28312));
    Span4Mux_v I__3536 (
            .O(N__28326),
            .I(N__28308));
    InMux I__3535 (
            .O(N__28325),
            .I(N__28305));
    LocalMux I__3534 (
            .O(N__28322),
            .I(N__28302));
    InMux I__3533 (
            .O(N__28321),
            .I(N__28299));
    Span4Mux_v I__3532 (
            .O(N__28318),
            .I(N__28292));
    LocalMux I__3531 (
            .O(N__28315),
            .I(N__28292));
    Span4Mux_h I__3530 (
            .O(N__28312),
            .I(N__28292));
    InMux I__3529 (
            .O(N__28311),
            .I(N__28289));
    Span4Mux_h I__3528 (
            .O(N__28308),
            .I(N__28286));
    LocalMux I__3527 (
            .O(N__28305),
            .I(encoder1_position_3));
    Odrv4 I__3526 (
            .O(N__28302),
            .I(encoder1_position_3));
    LocalMux I__3525 (
            .O(N__28299),
            .I(encoder1_position_3));
    Odrv4 I__3524 (
            .O(N__28292),
            .I(encoder1_position_3));
    LocalMux I__3523 (
            .O(N__28289),
            .I(encoder1_position_3));
    Odrv4 I__3522 (
            .O(N__28286),
            .I(encoder1_position_3));
    CascadeMux I__3521 (
            .O(N__28273),
            .I(\c0.n21071_cascade_ ));
    InMux I__3520 (
            .O(N__28270),
            .I(N__28266));
    InMux I__3519 (
            .O(N__28269),
            .I(N__28263));
    LocalMux I__3518 (
            .O(N__28266),
            .I(N__28258));
    LocalMux I__3517 (
            .O(N__28263),
            .I(N__28258));
    Odrv4 I__3516 (
            .O(N__28258),
            .I(data_out_frame_29__2__N_1749));
    InMux I__3515 (
            .O(N__28255),
            .I(N__28252));
    LocalMux I__3514 (
            .O(N__28252),
            .I(\c0.n17_adj_4501 ));
    InMux I__3513 (
            .O(N__28249),
            .I(N__28246));
    LocalMux I__3512 (
            .O(N__28246),
            .I(\c0.data_out_frame_29_0 ));
    InMux I__3511 (
            .O(N__28243),
            .I(N__28240));
    LocalMux I__3510 (
            .O(N__28240),
            .I(N__28237));
    Span4Mux_v I__3509 (
            .O(N__28237),
            .I(N__28234));
    Span4Mux_v I__3508 (
            .O(N__28234),
            .I(N__28231));
    Span4Mux_v I__3507 (
            .O(N__28231),
            .I(N__28228));
    Odrv4 I__3506 (
            .O(N__28228),
            .I(\c0.n26_adj_4423 ));
    InMux I__3505 (
            .O(N__28225),
            .I(N__28222));
    LocalMux I__3504 (
            .O(N__28222),
            .I(\c0.n16_adj_4500 ));
    CascadeMux I__3503 (
            .O(N__28219),
            .I(N__28215));
    CascadeMux I__3502 (
            .O(N__28218),
            .I(N__28212));
    InMux I__3501 (
            .O(N__28215),
            .I(N__28209));
    InMux I__3500 (
            .O(N__28212),
            .I(N__28206));
    LocalMux I__3499 (
            .O(N__28209),
            .I(N__28203));
    LocalMux I__3498 (
            .O(N__28206),
            .I(N__28200));
    Span4Mux_h I__3497 (
            .O(N__28203),
            .I(N__28195));
    Span4Mux_h I__3496 (
            .O(N__28200),
            .I(N__28195));
    Odrv4 I__3495 (
            .O(N__28195),
            .I(\c0.n10422 ));
    CascadeMux I__3494 (
            .O(N__28192),
            .I(\c0.n14_adj_4340_cascade_ ));
    InMux I__3493 (
            .O(N__28189),
            .I(N__28186));
    LocalMux I__3492 (
            .O(N__28186),
            .I(\c0.n20320 ));
    CascadeMux I__3491 (
            .O(N__28183),
            .I(\c0.n20320_cascade_ ));
    CascadeMux I__3490 (
            .O(N__28180),
            .I(\c0.n22180_cascade_ ));
    CascadeMux I__3489 (
            .O(N__28177),
            .I(\c0.n10498_cascade_ ));
    CascadeMux I__3488 (
            .O(N__28174),
            .I(\c0.n20253_cascade_ ));
    InMux I__3487 (
            .O(N__28171),
            .I(N__28166));
    InMux I__3486 (
            .O(N__28170),
            .I(N__28161));
    InMux I__3485 (
            .O(N__28169),
            .I(N__28161));
    LocalMux I__3484 (
            .O(N__28166),
            .I(N__28156));
    LocalMux I__3483 (
            .O(N__28161),
            .I(N__28156));
    Odrv4 I__3482 (
            .O(N__28156),
            .I(\c0.n21229 ));
    InMux I__3481 (
            .O(N__28153),
            .I(N__28150));
    LocalMux I__3480 (
            .O(N__28150),
            .I(\c0.n15_adj_4513 ));
    InMux I__3479 (
            .O(N__28147),
            .I(N__28144));
    LocalMux I__3478 (
            .O(N__28144),
            .I(\quad_counter0.n28_adj_4202 ));
    CascadeMux I__3477 (
            .O(N__28141),
            .I(\quad_counter0.n27_adj_4204_cascade_ ));
    InMux I__3476 (
            .O(N__28138),
            .I(N__28135));
    LocalMux I__3475 (
            .O(N__28135),
            .I(\quad_counter0.n25_adj_4205 ));
    InMux I__3474 (
            .O(N__28132),
            .I(N__28126));
    InMux I__3473 (
            .O(N__28131),
            .I(N__28126));
    LocalMux I__3472 (
            .O(N__28126),
            .I(n9821));
    InMux I__3471 (
            .O(N__28123),
            .I(N__28119));
    InMux I__3470 (
            .O(N__28122),
            .I(N__28116));
    LocalMux I__3469 (
            .O(N__28119),
            .I(\quad_counter0.a_delay_counter_12 ));
    LocalMux I__3468 (
            .O(N__28116),
            .I(\quad_counter0.a_delay_counter_12 ));
    InMux I__3467 (
            .O(N__28111),
            .I(N__28107));
    InMux I__3466 (
            .O(N__28110),
            .I(N__28104));
    LocalMux I__3465 (
            .O(N__28107),
            .I(\quad_counter0.a_delay_counter_13 ));
    LocalMux I__3464 (
            .O(N__28104),
            .I(\quad_counter0.a_delay_counter_13 ));
    CascadeMux I__3463 (
            .O(N__28099),
            .I(N__28095));
    InMux I__3462 (
            .O(N__28098),
            .I(N__28092));
    InMux I__3461 (
            .O(N__28095),
            .I(N__28089));
    LocalMux I__3460 (
            .O(N__28092),
            .I(\quad_counter0.a_delay_counter_6 ));
    LocalMux I__3459 (
            .O(N__28089),
            .I(\quad_counter0.a_delay_counter_6 ));
    InMux I__3458 (
            .O(N__28084),
            .I(N__28080));
    InMux I__3457 (
            .O(N__28083),
            .I(N__28077));
    LocalMux I__3456 (
            .O(N__28080),
            .I(\quad_counter0.a_delay_counter_9 ));
    LocalMux I__3455 (
            .O(N__28077),
            .I(\quad_counter0.a_delay_counter_9 ));
    InMux I__3454 (
            .O(N__28072),
            .I(N__28069));
    LocalMux I__3453 (
            .O(N__28069),
            .I(\quad_counter0.n26_adj_4203 ));
    InMux I__3452 (
            .O(N__28066),
            .I(N__28062));
    InMux I__3451 (
            .O(N__28065),
            .I(N__28059));
    LocalMux I__3450 (
            .O(N__28062),
            .I(N__28056));
    LocalMux I__3449 (
            .O(N__28059),
            .I(N__28053));
    Span4Mux_v I__3448 (
            .O(N__28056),
            .I(N__28050));
    Span4Mux_v I__3447 (
            .O(N__28053),
            .I(N__28047));
    Odrv4 I__3446 (
            .O(N__28050),
            .I(data_out_frame_28__3__N_1881));
    Odrv4 I__3445 (
            .O(N__28047),
            .I(data_out_frame_28__3__N_1881));
    CascadeMux I__3444 (
            .O(N__28042),
            .I(N__28039));
    InMux I__3443 (
            .O(N__28039),
            .I(N__28036));
    LocalMux I__3442 (
            .O(N__28036),
            .I(N__28032));
    InMux I__3441 (
            .O(N__28035),
            .I(N__28029));
    Span4Mux_h I__3440 (
            .O(N__28032),
            .I(N__28026));
    LocalMux I__3439 (
            .O(N__28029),
            .I(N__28023));
    Span4Mux_v I__3438 (
            .O(N__28026),
            .I(N__28020));
    Span4Mux_h I__3437 (
            .O(N__28023),
            .I(N__28017));
    Odrv4 I__3436 (
            .O(N__28020),
            .I(\c0.n20257 ));
    Odrv4 I__3435 (
            .O(N__28017),
            .I(\c0.n20257 ));
    InMux I__3434 (
            .O(N__28012),
            .I(N__28009));
    LocalMux I__3433 (
            .O(N__28009),
            .I(\c0.n21062 ));
    InMux I__3432 (
            .O(N__28006),
            .I(N__28003));
    LocalMux I__3431 (
            .O(N__28003),
            .I(N__28000));
    Odrv4 I__3430 (
            .O(N__28000),
            .I(\c0.data_out_frame_28_1 ));
    InMux I__3429 (
            .O(N__27997),
            .I(N__27994));
    LocalMux I__3428 (
            .O(N__27994),
            .I(\c0.data_out_frame_29_1 ));
    InMux I__3427 (
            .O(N__27991),
            .I(N__27988));
    LocalMux I__3426 (
            .O(N__27988),
            .I(N__27985));
    Span4Mux_v I__3425 (
            .O(N__27985),
            .I(N__27982));
    Span4Mux_v I__3424 (
            .O(N__27982),
            .I(N__27979));
    Odrv4 I__3423 (
            .O(N__27979),
            .I(\c0.n26_adj_4519 ));
    CascadeMux I__3422 (
            .O(N__27976),
            .I(\c0.n12542_cascade_ ));
    InMux I__3421 (
            .O(N__27973),
            .I(N__27966));
    InMux I__3420 (
            .O(N__27972),
            .I(N__27966));
    InMux I__3419 (
            .O(N__27971),
            .I(N__27963));
    LocalMux I__3418 (
            .O(N__27966),
            .I(\quad_counter0.B_delayed ));
    LocalMux I__3417 (
            .O(N__27963),
            .I(\quad_counter0.B_delayed ));
    InMux I__3416 (
            .O(N__27958),
            .I(N__27954));
    InMux I__3415 (
            .O(N__27957),
            .I(N__27951));
    LocalMux I__3414 (
            .O(N__27954),
            .I(\quad_counter0.a_delay_counter_3 ));
    LocalMux I__3413 (
            .O(N__27951),
            .I(\quad_counter0.a_delay_counter_3 ));
    InMux I__3412 (
            .O(N__27946),
            .I(N__27942));
    InMux I__3411 (
            .O(N__27945),
            .I(N__27939));
    LocalMux I__3410 (
            .O(N__27942),
            .I(\quad_counter0.a_delay_counter_8 ));
    LocalMux I__3409 (
            .O(N__27939),
            .I(\quad_counter0.a_delay_counter_8 ));
    CascadeMux I__3408 (
            .O(N__27934),
            .I(N__27930));
    InMux I__3407 (
            .O(N__27933),
            .I(N__27927));
    InMux I__3406 (
            .O(N__27930),
            .I(N__27924));
    LocalMux I__3405 (
            .O(N__27927),
            .I(\quad_counter0.a_delay_counter_2 ));
    LocalMux I__3404 (
            .O(N__27924),
            .I(\quad_counter0.a_delay_counter_2 ));
    InMux I__3403 (
            .O(N__27919),
            .I(N__27915));
    InMux I__3402 (
            .O(N__27918),
            .I(N__27912));
    LocalMux I__3401 (
            .O(N__27915),
            .I(\quad_counter0.a_delay_counter_1 ));
    LocalMux I__3400 (
            .O(N__27912),
            .I(\quad_counter0.a_delay_counter_1 ));
    InMux I__3399 (
            .O(N__27907),
            .I(N__27903));
    InMux I__3398 (
            .O(N__27906),
            .I(N__27900));
    LocalMux I__3397 (
            .O(N__27903),
            .I(\quad_counter0.a_delay_counter_5 ));
    LocalMux I__3396 (
            .O(N__27900),
            .I(\quad_counter0.a_delay_counter_5 ));
    InMux I__3395 (
            .O(N__27895),
            .I(N__27891));
    InMux I__3394 (
            .O(N__27894),
            .I(N__27888));
    LocalMux I__3393 (
            .O(N__27891),
            .I(\quad_counter0.a_delay_counter_11 ));
    LocalMux I__3392 (
            .O(N__27888),
            .I(\quad_counter0.a_delay_counter_11 ));
    CascadeMux I__3391 (
            .O(N__27883),
            .I(N__27879));
    InMux I__3390 (
            .O(N__27882),
            .I(N__27876));
    InMux I__3389 (
            .O(N__27879),
            .I(N__27873));
    LocalMux I__3388 (
            .O(N__27876),
            .I(\quad_counter0.a_delay_counter_4 ));
    LocalMux I__3387 (
            .O(N__27873),
            .I(\quad_counter0.a_delay_counter_4 ));
    CascadeMux I__3386 (
            .O(N__27868),
            .I(N__27865));
    InMux I__3385 (
            .O(N__27865),
            .I(N__27860));
    InMux I__3384 (
            .O(N__27864),
            .I(N__27855));
    InMux I__3383 (
            .O(N__27863),
            .I(N__27852));
    LocalMux I__3382 (
            .O(N__27860),
            .I(N__27849));
    InMux I__3381 (
            .O(N__27859),
            .I(N__27844));
    InMux I__3380 (
            .O(N__27858),
            .I(N__27844));
    LocalMux I__3379 (
            .O(N__27855),
            .I(N__27841));
    LocalMux I__3378 (
            .O(N__27852),
            .I(A_filtered));
    Odrv4 I__3377 (
            .O(N__27849),
            .I(A_filtered));
    LocalMux I__3376 (
            .O(N__27844),
            .I(A_filtered));
    Odrv4 I__3375 (
            .O(N__27841),
            .I(A_filtered));
    InMux I__3374 (
            .O(N__27832),
            .I(N__27826));
    InMux I__3373 (
            .O(N__27831),
            .I(N__27826));
    LocalMux I__3372 (
            .O(N__27826),
            .I(N__27821));
    InMux I__3371 (
            .O(N__27825),
            .I(N__27818));
    InMux I__3370 (
            .O(N__27824),
            .I(N__27815));
    Span4Mux_h I__3369 (
            .O(N__27821),
            .I(N__27808));
    LocalMux I__3368 (
            .O(N__27818),
            .I(N__27808));
    LocalMux I__3367 (
            .O(N__27815),
            .I(N__27808));
    Span4Mux_v I__3366 (
            .O(N__27808),
            .I(N__27805));
    Sp12to4 I__3365 (
            .O(N__27805),
            .I(N__27802));
    Odrv12 I__3364 (
            .O(N__27802),
            .I(PIN_7_c));
    CascadeMux I__3363 (
            .O(N__27799),
            .I(N__27796));
    InMux I__3362 (
            .O(N__27796),
            .I(N__27790));
    InMux I__3361 (
            .O(N__27795),
            .I(N__27790));
    LocalMux I__3360 (
            .O(N__27790),
            .I(N__27786));
    InMux I__3359 (
            .O(N__27789),
            .I(N__27783));
    Span4Mux_h I__3358 (
            .O(N__27786),
            .I(N__27780));
    LocalMux I__3357 (
            .O(N__27783),
            .I(N__27777));
    Odrv4 I__3356 (
            .O(N__27780),
            .I(quadA_delayed));
    Odrv4 I__3355 (
            .O(N__27777),
            .I(quadA_delayed));
    CEMux I__3354 (
            .O(N__27772),
            .I(N__27769));
    LocalMux I__3353 (
            .O(N__27769),
            .I(N__27765));
    CEMux I__3352 (
            .O(N__27768),
            .I(N__27762));
    Span4Mux_h I__3351 (
            .O(N__27765),
            .I(N__27759));
    LocalMux I__3350 (
            .O(N__27762),
            .I(N__27756));
    Span4Mux_h I__3349 (
            .O(N__27759),
            .I(N__27753));
    Odrv4 I__3348 (
            .O(N__27756),
            .I(n14421));
    Odrv4 I__3347 (
            .O(N__27753),
            .I(n14421));
    SRMux I__3346 (
            .O(N__27748),
            .I(N__27743));
    SRMux I__3345 (
            .O(N__27747),
            .I(N__27740));
    InMux I__3344 (
            .O(N__27746),
            .I(N__27737));
    LocalMux I__3343 (
            .O(N__27743),
            .I(N__27734));
    LocalMux I__3342 (
            .O(N__27740),
            .I(N__27729));
    LocalMux I__3341 (
            .O(N__27737),
            .I(N__27729));
    Odrv4 I__3340 (
            .O(N__27734),
            .I(a_delay_counter_15__N_4124));
    Odrv4 I__3339 (
            .O(N__27729),
            .I(a_delay_counter_15__N_4124));
    InMux I__3338 (
            .O(N__27724),
            .I(N__27721));
    LocalMux I__3337 (
            .O(N__27721),
            .I(n39));
    CascadeMux I__3336 (
            .O(N__27718),
            .I(n14421_cascade_));
    InMux I__3335 (
            .O(N__27715),
            .I(N__27710));
    InMux I__3334 (
            .O(N__27714),
            .I(N__27707));
    InMux I__3333 (
            .O(N__27713),
            .I(N__27704));
    LocalMux I__3332 (
            .O(N__27710),
            .I(a_delay_counter_0));
    LocalMux I__3331 (
            .O(N__27707),
            .I(a_delay_counter_0));
    LocalMux I__3330 (
            .O(N__27704),
            .I(a_delay_counter_0));
    InMux I__3329 (
            .O(N__27697),
            .I(N__27693));
    InMux I__3328 (
            .O(N__27696),
            .I(N__27690));
    LocalMux I__3327 (
            .O(N__27693),
            .I(\quad_counter0.a_delay_counter_14 ));
    LocalMux I__3326 (
            .O(N__27690),
            .I(\quad_counter0.a_delay_counter_14 ));
    InMux I__3325 (
            .O(N__27685),
            .I(N__27681));
    InMux I__3324 (
            .O(N__27684),
            .I(N__27678));
    LocalMux I__3323 (
            .O(N__27681),
            .I(\quad_counter0.a_delay_counter_15 ));
    LocalMux I__3322 (
            .O(N__27678),
            .I(\quad_counter0.a_delay_counter_15 ));
    CascadeMux I__3321 (
            .O(N__27673),
            .I(N__27669));
    InMux I__3320 (
            .O(N__27672),
            .I(N__27666));
    InMux I__3319 (
            .O(N__27669),
            .I(N__27663));
    LocalMux I__3318 (
            .O(N__27666),
            .I(\quad_counter0.a_delay_counter_7 ));
    LocalMux I__3317 (
            .O(N__27663),
            .I(\quad_counter0.a_delay_counter_7 ));
    InMux I__3316 (
            .O(N__27658),
            .I(N__27654));
    InMux I__3315 (
            .O(N__27657),
            .I(N__27651));
    LocalMux I__3314 (
            .O(N__27654),
            .I(\quad_counter0.a_delay_counter_10 ));
    LocalMux I__3313 (
            .O(N__27651),
            .I(\quad_counter0.a_delay_counter_10 ));
    InMux I__3312 (
            .O(N__27646),
            .I(N__27642));
    InMux I__3311 (
            .O(N__27645),
            .I(N__27639));
    LocalMux I__3310 (
            .O(N__27642),
            .I(\quad_counter0.b_delay_counter_3 ));
    LocalMux I__3309 (
            .O(N__27639),
            .I(\quad_counter0.b_delay_counter_3 ));
    InMux I__3308 (
            .O(N__27634),
            .I(N__27630));
    InMux I__3307 (
            .O(N__27633),
            .I(N__27627));
    LocalMux I__3306 (
            .O(N__27630),
            .I(\quad_counter0.b_delay_counter_9 ));
    LocalMux I__3305 (
            .O(N__27627),
            .I(\quad_counter0.b_delay_counter_9 ));
    CascadeMux I__3304 (
            .O(N__27622),
            .I(N__27618));
    InMux I__3303 (
            .O(N__27621),
            .I(N__27615));
    InMux I__3302 (
            .O(N__27618),
            .I(N__27612));
    LocalMux I__3301 (
            .O(N__27615),
            .I(\quad_counter0.b_delay_counter_4 ));
    LocalMux I__3300 (
            .O(N__27612),
            .I(\quad_counter0.b_delay_counter_4 ));
    CascadeMux I__3299 (
            .O(N__27607),
            .I(N__27603));
    InMux I__3298 (
            .O(N__27606),
            .I(N__27599));
    InMux I__3297 (
            .O(N__27603),
            .I(N__27596));
    InMux I__3296 (
            .O(N__27602),
            .I(N__27593));
    LocalMux I__3295 (
            .O(N__27599),
            .I(N__27590));
    LocalMux I__3294 (
            .O(N__27596),
            .I(b_delay_counter_0));
    LocalMux I__3293 (
            .O(N__27593),
            .I(b_delay_counter_0));
    Odrv4 I__3292 (
            .O(N__27590),
            .I(b_delay_counter_0));
    InMux I__3291 (
            .O(N__27583),
            .I(N__27580));
    LocalMux I__3290 (
            .O(N__27580),
            .I(N__27575));
    InMux I__3289 (
            .O(N__27579),
            .I(N__27569));
    InMux I__3288 (
            .O(N__27578),
            .I(N__27569));
    Span4Mux_v I__3287 (
            .O(N__27575),
            .I(N__27566));
    InMux I__3286 (
            .O(N__27574),
            .I(N__27563));
    LocalMux I__3285 (
            .O(N__27569),
            .I(N__27560));
    Span4Mux_h I__3284 (
            .O(N__27566),
            .I(N__27555));
    LocalMux I__3283 (
            .O(N__27563),
            .I(N__27555));
    Sp12to4 I__3282 (
            .O(N__27560),
            .I(N__27552));
    Span4Mux_h I__3281 (
            .O(N__27555),
            .I(N__27549));
    Span12Mux_v I__3280 (
            .O(N__27552),
            .I(N__27546));
    Span4Mux_v I__3279 (
            .O(N__27549),
            .I(N__27543));
    Odrv12 I__3278 (
            .O(N__27546),
            .I(PIN_8_c));
    Odrv4 I__3277 (
            .O(N__27543),
            .I(PIN_8_c));
    CascadeMux I__3276 (
            .O(N__27538),
            .I(N__27535));
    InMux I__3275 (
            .O(N__27535),
            .I(N__27532));
    LocalMux I__3274 (
            .O(N__27532),
            .I(N__27527));
    InMux I__3273 (
            .O(N__27531),
            .I(N__27522));
    InMux I__3272 (
            .O(N__27530),
            .I(N__27522));
    Span4Mux_v I__3271 (
            .O(N__27527),
            .I(N__27519));
    LocalMux I__3270 (
            .O(N__27522),
            .I(N__27516));
    Span4Mux_h I__3269 (
            .O(N__27519),
            .I(N__27513));
    Span4Mux_v I__3268 (
            .O(N__27516),
            .I(N__27510));
    Odrv4 I__3267 (
            .O(N__27513),
            .I(quadB_delayed));
    Odrv4 I__3266 (
            .O(N__27510),
            .I(quadB_delayed));
    InMux I__3265 (
            .O(N__27505),
            .I(N__27496));
    InMux I__3264 (
            .O(N__27504),
            .I(N__27496));
    InMux I__3263 (
            .O(N__27503),
            .I(N__27496));
    LocalMux I__3262 (
            .O(N__27496),
            .I(B_filtered));
    InMux I__3261 (
            .O(N__27493),
            .I(N__27489));
    InMux I__3260 (
            .O(N__27492),
            .I(N__27486));
    LocalMux I__3259 (
            .O(N__27489),
            .I(\quad_counter0.b_delay_counter_13 ));
    LocalMux I__3258 (
            .O(N__27486),
            .I(\quad_counter0.b_delay_counter_13 ));
    InMux I__3257 (
            .O(N__27481),
            .I(N__27477));
    InMux I__3256 (
            .O(N__27480),
            .I(N__27474));
    LocalMux I__3255 (
            .O(N__27477),
            .I(\quad_counter0.b_delay_counter_1 ));
    LocalMux I__3254 (
            .O(N__27474),
            .I(\quad_counter0.b_delay_counter_1 ));
    CascadeMux I__3253 (
            .O(N__27469),
            .I(N__27465));
    InMux I__3252 (
            .O(N__27468),
            .I(N__27462));
    InMux I__3251 (
            .O(N__27465),
            .I(N__27459));
    LocalMux I__3250 (
            .O(N__27462),
            .I(\quad_counter0.b_delay_counter_2 ));
    LocalMux I__3249 (
            .O(N__27459),
            .I(\quad_counter0.b_delay_counter_2 ));
    InMux I__3248 (
            .O(N__27454),
            .I(N__27450));
    InMux I__3247 (
            .O(N__27453),
            .I(N__27447));
    LocalMux I__3246 (
            .O(N__27450),
            .I(\quad_counter0.b_delay_counter_5 ));
    LocalMux I__3245 (
            .O(N__27447),
            .I(\quad_counter0.b_delay_counter_5 ));
    InMux I__3244 (
            .O(N__27442),
            .I(N__27438));
    InMux I__3243 (
            .O(N__27441),
            .I(N__27435));
    LocalMux I__3242 (
            .O(N__27438),
            .I(\quad_counter0.b_delay_counter_11 ));
    LocalMux I__3241 (
            .O(N__27435),
            .I(\quad_counter0.b_delay_counter_11 ));
    InMux I__3240 (
            .O(N__27430),
            .I(N__27426));
    InMux I__3239 (
            .O(N__27429),
            .I(N__27423));
    LocalMux I__3238 (
            .O(N__27426),
            .I(\quad_counter0.b_delay_counter_10 ));
    LocalMux I__3237 (
            .O(N__27423),
            .I(\quad_counter0.b_delay_counter_10 ));
    CascadeMux I__3236 (
            .O(N__27418),
            .I(N__27414));
    InMux I__3235 (
            .O(N__27417),
            .I(N__27411));
    InMux I__3234 (
            .O(N__27414),
            .I(N__27408));
    LocalMux I__3233 (
            .O(N__27411),
            .I(\quad_counter0.b_delay_counter_8 ));
    LocalMux I__3232 (
            .O(N__27408),
            .I(\quad_counter0.b_delay_counter_8 ));
    InMux I__3231 (
            .O(N__27403),
            .I(N__27399));
    InMux I__3230 (
            .O(N__27402),
            .I(N__27396));
    LocalMux I__3229 (
            .O(N__27399),
            .I(\quad_counter0.b_delay_counter_6 ));
    LocalMux I__3228 (
            .O(N__27396),
            .I(\quad_counter0.b_delay_counter_6 ));
    InMux I__3227 (
            .O(N__27391),
            .I(N__27388));
    LocalMux I__3226 (
            .O(N__27388),
            .I(\quad_counter0.n28_adj_4198 ));
    CascadeMux I__3225 (
            .O(N__27385),
            .I(\quad_counter0.n26_adj_4199_cascade_ ));
    InMux I__3224 (
            .O(N__27382),
            .I(N__27379));
    LocalMux I__3223 (
            .O(N__27379),
            .I(\quad_counter0.n25_adj_4201 ));
    InMux I__3222 (
            .O(N__27376),
            .I(N__27373));
    LocalMux I__3221 (
            .O(N__27373),
            .I(N__27369));
    InMux I__3220 (
            .O(N__27372),
            .I(N__27366));
    Span4Mux_h I__3219 (
            .O(N__27369),
            .I(N__27363));
    LocalMux I__3218 (
            .O(N__27366),
            .I(n12909));
    Odrv4 I__3217 (
            .O(N__27363),
            .I(n12909));
    InMux I__3216 (
            .O(N__27358),
            .I(N__27355));
    LocalMux I__3215 (
            .O(N__27355),
            .I(\quad_counter0.A_delayed ));
    InMux I__3214 (
            .O(N__27352),
            .I(N__27349));
    LocalMux I__3213 (
            .O(N__27349),
            .I(N__27346));
    Odrv4 I__3212 (
            .O(N__27346),
            .I(n10_adj_4535));
    CascadeMux I__3211 (
            .O(N__27343),
            .I(N__27339));
    CascadeMux I__3210 (
            .O(N__27342),
            .I(N__27335));
    InMux I__3209 (
            .O(N__27339),
            .I(N__27331));
    InMux I__3208 (
            .O(N__27338),
            .I(N__27326));
    InMux I__3207 (
            .O(N__27335),
            .I(N__27323));
    CascadeMux I__3206 (
            .O(N__27334),
            .I(N__27319));
    LocalMux I__3205 (
            .O(N__27331),
            .I(N__27316));
    InMux I__3204 (
            .O(N__27330),
            .I(N__27311));
    InMux I__3203 (
            .O(N__27329),
            .I(N__27311));
    LocalMux I__3202 (
            .O(N__27326),
            .I(N__27305));
    LocalMux I__3201 (
            .O(N__27323),
            .I(N__27302));
    InMux I__3200 (
            .O(N__27322),
            .I(N__27297));
    InMux I__3199 (
            .O(N__27319),
            .I(N__27297));
    Span4Mux_v I__3198 (
            .O(N__27316),
            .I(N__27292));
    LocalMux I__3197 (
            .O(N__27311),
            .I(N__27292));
    InMux I__3196 (
            .O(N__27310),
            .I(N__27289));
    InMux I__3195 (
            .O(N__27309),
            .I(N__27286));
    InMux I__3194 (
            .O(N__27308),
            .I(N__27283));
    Span4Mux_h I__3193 (
            .O(N__27305),
            .I(N__27280));
    Span4Mux_h I__3192 (
            .O(N__27302),
            .I(N__27277));
    LocalMux I__3191 (
            .O(N__27297),
            .I(N__27272));
    Span4Mux_h I__3190 (
            .O(N__27292),
            .I(N__27272));
    LocalMux I__3189 (
            .O(N__27289),
            .I(N__27269));
    LocalMux I__3188 (
            .O(N__27286),
            .I(byte_transmit_counter_5));
    LocalMux I__3187 (
            .O(N__27283),
            .I(byte_transmit_counter_5));
    Odrv4 I__3186 (
            .O(N__27280),
            .I(byte_transmit_counter_5));
    Odrv4 I__3185 (
            .O(N__27277),
            .I(byte_transmit_counter_5));
    Odrv4 I__3184 (
            .O(N__27272),
            .I(byte_transmit_counter_5));
    Odrv12 I__3183 (
            .O(N__27269),
            .I(byte_transmit_counter_5));
    InMux I__3182 (
            .O(N__27256),
            .I(N__27250));
    InMux I__3181 (
            .O(N__27255),
            .I(N__27250));
    LocalMux I__3180 (
            .O(N__27250),
            .I(r_Tx_Data_1));
    CascadeMux I__3179 (
            .O(N__27247),
            .I(N__27242));
    CascadeMux I__3178 (
            .O(N__27246),
            .I(N__27239));
    InMux I__3177 (
            .O(N__27245),
            .I(N__27232));
    InMux I__3176 (
            .O(N__27242),
            .I(N__27232));
    InMux I__3175 (
            .O(N__27239),
            .I(N__27232));
    LocalMux I__3174 (
            .O(N__27232),
            .I(data_in_0_7));
    CascadeMux I__3173 (
            .O(N__27229),
            .I(N__27225));
    InMux I__3172 (
            .O(N__27228),
            .I(N__27222));
    InMux I__3171 (
            .O(N__27225),
            .I(N__27219));
    LocalMux I__3170 (
            .O(N__27222),
            .I(N__27214));
    LocalMux I__3169 (
            .O(N__27219),
            .I(N__27214));
    Odrv4 I__3168 (
            .O(N__27214),
            .I(data_out_frame_5_3));
    InMux I__3167 (
            .O(N__27211),
            .I(N__27207));
    InMux I__3166 (
            .O(N__27210),
            .I(N__27204));
    LocalMux I__3165 (
            .O(N__27207),
            .I(N__27201));
    LocalMux I__3164 (
            .O(N__27204),
            .I(data_out_frame_6_3));
    Odrv12 I__3163 (
            .O(N__27201),
            .I(data_out_frame_6_3));
    CascadeMux I__3162 (
            .O(N__27196),
            .I(N__27193));
    InMux I__3161 (
            .O(N__27193),
            .I(N__27190));
    LocalMux I__3160 (
            .O(N__27190),
            .I(N__27187));
    Span4Mux_h I__3159 (
            .O(N__27187),
            .I(N__27184));
    Odrv4 I__3158 (
            .O(N__27184),
            .I(\c0.n5 ));
    CascadeMux I__3157 (
            .O(N__27181),
            .I(N__27177));
    CascadeMux I__3156 (
            .O(N__27180),
            .I(N__27174));
    InMux I__3155 (
            .O(N__27177),
            .I(N__27171));
    InMux I__3154 (
            .O(N__27174),
            .I(N__27168));
    LocalMux I__3153 (
            .O(N__27171),
            .I(N__27165));
    LocalMux I__3152 (
            .O(N__27168),
            .I(N__27160));
    Span4Mux_h I__3151 (
            .O(N__27165),
            .I(N__27160));
    Odrv4 I__3150 (
            .O(N__27160),
            .I(data_out_frame_5_5));
    InMux I__3149 (
            .O(N__27157),
            .I(N__27153));
    InMux I__3148 (
            .O(N__27156),
            .I(N__27150));
    LocalMux I__3147 (
            .O(N__27153),
            .I(N__27147));
    LocalMux I__3146 (
            .O(N__27150),
            .I(data_out_frame_11_0));
    Odrv4 I__3145 (
            .O(N__27147),
            .I(data_out_frame_11_0));
    CascadeMux I__3144 (
            .O(N__27142),
            .I(\c0.n24165_cascade_ ));
    InMux I__3143 (
            .O(N__27139),
            .I(N__27136));
    LocalMux I__3142 (
            .O(N__27136),
            .I(\c0.n24168 ));
    CascadeMux I__3141 (
            .O(N__27133),
            .I(N__27130));
    InMux I__3140 (
            .O(N__27130),
            .I(N__27127));
    LocalMux I__3139 (
            .O(N__27127),
            .I(\c0.n11_adj_4218 ));
    CascadeMux I__3138 (
            .O(N__27124),
            .I(N__27120));
    InMux I__3137 (
            .O(N__27123),
            .I(N__27115));
    InMux I__3136 (
            .O(N__27120),
            .I(N__27115));
    LocalMux I__3135 (
            .O(N__27115),
            .I(data_out_frame_11_5));
    InMux I__3134 (
            .O(N__27112),
            .I(N__27109));
    LocalMux I__3133 (
            .O(N__27109),
            .I(N__27105));
    InMux I__3132 (
            .O(N__27108),
            .I(N__27102));
    Span4Mux_v I__3131 (
            .O(N__27105),
            .I(N__27099));
    LocalMux I__3130 (
            .O(N__27102),
            .I(data_out_frame_9_5));
    Odrv4 I__3129 (
            .O(N__27099),
            .I(data_out_frame_9_5));
    CascadeMux I__3128 (
            .O(N__27094),
            .I(\c0.n24141_cascade_ ));
    CascadeMux I__3127 (
            .O(N__27091),
            .I(N__27088));
    InMux I__3126 (
            .O(N__27088),
            .I(N__27082));
    InMux I__3125 (
            .O(N__27087),
            .I(N__27082));
    LocalMux I__3124 (
            .O(N__27082),
            .I(data_out_frame_8_5));
    InMux I__3123 (
            .O(N__27079),
            .I(N__27076));
    LocalMux I__3122 (
            .O(N__27076),
            .I(N__27073));
    Odrv4 I__3121 (
            .O(N__27073),
            .I(\c0.n24144 ));
    CascadeMux I__3120 (
            .O(N__27070),
            .I(N__27067));
    InMux I__3119 (
            .O(N__27067),
            .I(N__27063));
    InMux I__3118 (
            .O(N__27066),
            .I(N__27060));
    LocalMux I__3117 (
            .O(N__27063),
            .I(r_Tx_Data_7));
    LocalMux I__3116 (
            .O(N__27060),
            .I(r_Tx_Data_7));
    InMux I__3115 (
            .O(N__27055),
            .I(N__27051));
    InMux I__3114 (
            .O(N__27054),
            .I(N__27048));
    LocalMux I__3113 (
            .O(N__27051),
            .I(r_Tx_Data_3));
    LocalMux I__3112 (
            .O(N__27048),
            .I(r_Tx_Data_3));
    InMux I__3111 (
            .O(N__27043),
            .I(N__27037));
    InMux I__3110 (
            .O(N__27042),
            .I(N__27029));
    InMux I__3109 (
            .O(N__27041),
            .I(N__27029));
    InMux I__3108 (
            .O(N__27040),
            .I(N__27029));
    LocalMux I__3107 (
            .O(N__27037),
            .I(N__27026));
    InMux I__3106 (
            .O(N__27036),
            .I(N__27023));
    LocalMux I__3105 (
            .O(N__27029),
            .I(r_Bit_Index_2_adj_4551));
    Odrv4 I__3104 (
            .O(N__27026),
            .I(r_Bit_Index_2_adj_4551));
    LocalMux I__3103 (
            .O(N__27023),
            .I(r_Bit_Index_2_adj_4551));
    InMux I__3102 (
            .O(N__27016),
            .I(N__27013));
    LocalMux I__3101 (
            .O(N__27013),
            .I(N__27010));
    Span4Mux_h I__3100 (
            .O(N__27010),
            .I(N__27006));
    InMux I__3099 (
            .O(N__27009),
            .I(N__27003));
    Span4Mux_h I__3098 (
            .O(N__27006),
            .I(N__27000));
    LocalMux I__3097 (
            .O(N__27003),
            .I(N__26997));
    Odrv4 I__3096 (
            .O(N__27000),
            .I(n4_adj_4554));
    Odrv4 I__3095 (
            .O(N__26997),
            .I(n4_adj_4554));
    CascadeMux I__3094 (
            .O(N__26992),
            .I(n24189_cascade_));
    CascadeMux I__3093 (
            .O(N__26989),
            .I(N__26984));
    InMux I__3092 (
            .O(N__26988),
            .I(N__26979));
    InMux I__3091 (
            .O(N__26987),
            .I(N__26979));
    InMux I__3090 (
            .O(N__26984),
            .I(N__26975));
    LocalMux I__3089 (
            .O(N__26979),
            .I(N__26972));
    CascadeMux I__3088 (
            .O(N__26978),
            .I(N__26967));
    LocalMux I__3087 (
            .O(N__26975),
            .I(N__26963));
    Span4Mux_h I__3086 (
            .O(N__26972),
            .I(N__26960));
    InMux I__3085 (
            .O(N__26971),
            .I(N__26953));
    InMux I__3084 (
            .O(N__26970),
            .I(N__26953));
    InMux I__3083 (
            .O(N__26967),
            .I(N__26953));
    InMux I__3082 (
            .O(N__26966),
            .I(N__26950));
    Span4Mux_v I__3081 (
            .O(N__26963),
            .I(N__26947));
    Odrv4 I__3080 (
            .O(N__26960),
            .I(r_Bit_Index_1_adj_4552));
    LocalMux I__3079 (
            .O(N__26953),
            .I(r_Bit_Index_1_adj_4552));
    LocalMux I__3078 (
            .O(N__26950),
            .I(r_Bit_Index_1_adj_4552));
    Odrv4 I__3077 (
            .O(N__26947),
            .I(r_Bit_Index_1_adj_4552));
    InMux I__3076 (
            .O(N__26938),
            .I(N__26935));
    LocalMux I__3075 (
            .O(N__26935),
            .I(\c0.n6_adj_4392 ));
    InMux I__3074 (
            .O(N__26932),
            .I(N__26928));
    InMux I__3073 (
            .O(N__26931),
            .I(N__26925));
    LocalMux I__3072 (
            .O(N__26928),
            .I(N__26922));
    LocalMux I__3071 (
            .O(N__26925),
            .I(N__26917));
    Span4Mux_h I__3070 (
            .O(N__26922),
            .I(N__26917));
    Odrv4 I__3069 (
            .O(N__26917),
            .I(\c0.byte_transmit_counter_6 ));
    CascadeMux I__3068 (
            .O(N__26914),
            .I(\c0.n23574_cascade_ ));
    InMux I__3067 (
            .O(N__26911),
            .I(N__26907));
    InMux I__3066 (
            .O(N__26910),
            .I(N__26904));
    LocalMux I__3065 (
            .O(N__26907),
            .I(N__26901));
    LocalMux I__3064 (
            .O(N__26904),
            .I(\c0.byte_transmit_counter_7 ));
    Odrv12 I__3063 (
            .O(N__26901),
            .I(\c0.byte_transmit_counter_7 ));
    CascadeMux I__3062 (
            .O(N__26896),
            .I(\c0.n38_adj_4387_cascade_ ));
    CascadeMux I__3061 (
            .O(N__26893),
            .I(N__26890));
    InMux I__3060 (
            .O(N__26890),
            .I(N__26886));
    InMux I__3059 (
            .O(N__26889),
            .I(N__26883));
    LocalMux I__3058 (
            .O(N__26886),
            .I(N__26880));
    LocalMux I__3057 (
            .O(N__26883),
            .I(data_out_frame_5_2));
    Odrv4 I__3056 (
            .O(N__26880),
            .I(data_out_frame_5_2));
    InMux I__3055 (
            .O(N__26875),
            .I(N__26870));
    CascadeMux I__3054 (
            .O(N__26874),
            .I(N__26867));
    InMux I__3053 (
            .O(N__26873),
            .I(N__26860));
    LocalMux I__3052 (
            .O(N__26870),
            .I(N__26857));
    InMux I__3051 (
            .O(N__26867),
            .I(N__26854));
    InMux I__3050 (
            .O(N__26866),
            .I(N__26851));
    InMux I__3049 (
            .O(N__26865),
            .I(N__26848));
    CascadeMux I__3048 (
            .O(N__26864),
            .I(N__26845));
    CascadeMux I__3047 (
            .O(N__26863),
            .I(N__26842));
    LocalMux I__3046 (
            .O(N__26860),
            .I(N__26839));
    Span4Mux_v I__3045 (
            .O(N__26857),
            .I(N__26834));
    LocalMux I__3044 (
            .O(N__26854),
            .I(N__26834));
    LocalMux I__3043 (
            .O(N__26851),
            .I(N__26831));
    LocalMux I__3042 (
            .O(N__26848),
            .I(N__26828));
    InMux I__3041 (
            .O(N__26845),
            .I(N__26825));
    InMux I__3040 (
            .O(N__26842),
            .I(N__26822));
    Span4Mux_h I__3039 (
            .O(N__26839),
            .I(N__26819));
    Span4Mux_v I__3038 (
            .O(N__26834),
            .I(N__26814));
    Span4Mux_v I__3037 (
            .O(N__26831),
            .I(N__26814));
    Span4Mux_h I__3036 (
            .O(N__26828),
            .I(N__26811));
    LocalMux I__3035 (
            .O(N__26825),
            .I(N__26806));
    LocalMux I__3034 (
            .O(N__26822),
            .I(N__26806));
    Odrv4 I__3033 (
            .O(N__26819),
            .I(n23768));
    Odrv4 I__3032 (
            .O(N__26814),
            .I(n23768));
    Odrv4 I__3031 (
            .O(N__26811),
            .I(n23768));
    Odrv12 I__3030 (
            .O(N__26806),
            .I(n23768));
    CascadeMux I__3029 (
            .O(N__26797),
            .I(N__26793));
    CascadeMux I__3028 (
            .O(N__26796),
            .I(N__26785));
    InMux I__3027 (
            .O(N__26793),
            .I(N__26776));
    InMux I__3026 (
            .O(N__26792),
            .I(N__26771));
    InMux I__3025 (
            .O(N__26791),
            .I(N__26771));
    InMux I__3024 (
            .O(N__26790),
            .I(N__26766));
    InMux I__3023 (
            .O(N__26789),
            .I(N__26766));
    InMux I__3022 (
            .O(N__26788),
            .I(N__26761));
    InMux I__3021 (
            .O(N__26785),
            .I(N__26761));
    InMux I__3020 (
            .O(N__26784),
            .I(N__26756));
    InMux I__3019 (
            .O(N__26783),
            .I(N__26756));
    InMux I__3018 (
            .O(N__26782),
            .I(N__26749));
    InMux I__3017 (
            .O(N__26781),
            .I(N__26749));
    InMux I__3016 (
            .O(N__26780),
            .I(N__26749));
    InMux I__3015 (
            .O(N__26779),
            .I(N__26746));
    LocalMux I__3014 (
            .O(N__26776),
            .I(N__26739));
    LocalMux I__3013 (
            .O(N__26771),
            .I(N__26736));
    LocalMux I__3012 (
            .O(N__26766),
            .I(N__26733));
    LocalMux I__3011 (
            .O(N__26761),
            .I(N__26730));
    LocalMux I__3010 (
            .O(N__26756),
            .I(N__26723));
    LocalMux I__3009 (
            .O(N__26749),
            .I(N__26723));
    LocalMux I__3008 (
            .O(N__26746),
            .I(N__26723));
    InMux I__3007 (
            .O(N__26745),
            .I(N__26720));
    InMux I__3006 (
            .O(N__26744),
            .I(N__26715));
    InMux I__3005 (
            .O(N__26743),
            .I(N__26715));
    InMux I__3004 (
            .O(N__26742),
            .I(N__26712));
    Span4Mux_h I__3003 (
            .O(N__26739),
            .I(N__26709));
    Span4Mux_h I__3002 (
            .O(N__26736),
            .I(N__26704));
    Span4Mux_h I__3001 (
            .O(N__26733),
            .I(N__26704));
    Span4Mux_h I__3000 (
            .O(N__26730),
            .I(N__26701));
    Span4Mux_v I__2999 (
            .O(N__26723),
            .I(N__26696));
    LocalMux I__2998 (
            .O(N__26720),
            .I(N__26696));
    LocalMux I__2997 (
            .O(N__26715),
            .I(byte_transmit_counter_4));
    LocalMux I__2996 (
            .O(N__26712),
            .I(byte_transmit_counter_4));
    Odrv4 I__2995 (
            .O(N__26709),
            .I(byte_transmit_counter_4));
    Odrv4 I__2994 (
            .O(N__26704),
            .I(byte_transmit_counter_4));
    Odrv4 I__2993 (
            .O(N__26701),
            .I(byte_transmit_counter_4));
    Odrv4 I__2992 (
            .O(N__26696),
            .I(byte_transmit_counter_4));
    InMux I__2991 (
            .O(N__26683),
            .I(N__26680));
    LocalMux I__2990 (
            .O(N__26680),
            .I(n23864));
    InMux I__2989 (
            .O(N__26677),
            .I(N__26674));
    LocalMux I__2988 (
            .O(N__26674),
            .I(N__26670));
    InMux I__2987 (
            .O(N__26673),
            .I(N__26667));
    Span4Mux_h I__2986 (
            .O(N__26670),
            .I(N__26664));
    LocalMux I__2985 (
            .O(N__26667),
            .I(data_out_frame_5_6));
    Odrv4 I__2984 (
            .O(N__26664),
            .I(data_out_frame_5_6));
    InMux I__2983 (
            .O(N__26659),
            .I(N__26655));
    InMux I__2982 (
            .O(N__26658),
            .I(N__26652));
    LocalMux I__2981 (
            .O(N__26655),
            .I(N__26649));
    LocalMux I__2980 (
            .O(N__26652),
            .I(data_out_frame_13_3));
    Odrv4 I__2979 (
            .O(N__26649),
            .I(data_out_frame_13_3));
    InMux I__2978 (
            .O(N__26644),
            .I(N__26641));
    LocalMux I__2977 (
            .O(N__26641),
            .I(n2184));
    InMux I__2976 (
            .O(N__26638),
            .I(N__26635));
    LocalMux I__2975 (
            .O(N__26635),
            .I(n2182));
    InMux I__2974 (
            .O(N__26632),
            .I(N__26629));
    LocalMux I__2973 (
            .O(N__26629),
            .I(n2176));
    InMux I__2972 (
            .O(N__26626),
            .I(N__26623));
    LocalMux I__2971 (
            .O(N__26623),
            .I(N__26619));
    InMux I__2970 (
            .O(N__26622),
            .I(N__26616));
    Span4Mux_v I__2969 (
            .O(N__26619),
            .I(N__26613));
    LocalMux I__2968 (
            .O(N__26616),
            .I(data_out_frame_29_3));
    Odrv4 I__2967 (
            .O(N__26613),
            .I(data_out_frame_29_3));
    CascadeMux I__2966 (
            .O(N__26608),
            .I(N__26604));
    InMux I__2965 (
            .O(N__26607),
            .I(N__26601));
    InMux I__2964 (
            .O(N__26604),
            .I(N__26598));
    LocalMux I__2963 (
            .O(N__26601),
            .I(N__26595));
    LocalMux I__2962 (
            .O(N__26598),
            .I(data_out_frame_28_3));
    Odrv12 I__2961 (
            .O(N__26595),
            .I(data_out_frame_28_3));
    InMux I__2960 (
            .O(N__26590),
            .I(N__26587));
    LocalMux I__2959 (
            .O(N__26587),
            .I(N__26584));
    Odrv4 I__2958 (
            .O(N__26584),
            .I(\c0.n26 ));
    InMux I__2957 (
            .O(N__26581),
            .I(N__26578));
    LocalMux I__2956 (
            .O(N__26578),
            .I(n2175));
    InMux I__2955 (
            .O(N__26575),
            .I(N__26572));
    LocalMux I__2954 (
            .O(N__26572),
            .I(N__26568));
    InMux I__2953 (
            .O(N__26571),
            .I(N__26565));
    Span4Mux_h I__2952 (
            .O(N__26568),
            .I(N__26562));
    LocalMux I__2951 (
            .O(N__26565),
            .I(data_out_frame_7_5));
    Odrv4 I__2950 (
            .O(N__26562),
            .I(data_out_frame_7_5));
    CascadeMux I__2949 (
            .O(N__26557),
            .I(N__26554));
    InMux I__2948 (
            .O(N__26554),
            .I(N__26551));
    LocalMux I__2947 (
            .O(N__26551),
            .I(N__26548));
    Span4Mux_h I__2946 (
            .O(N__26548),
            .I(N__26545));
    Odrv4 I__2945 (
            .O(N__26545),
            .I(\c0.n5_adj_4346 ));
    InMux I__2944 (
            .O(N__26542),
            .I(N__26538));
    InMux I__2943 (
            .O(N__26541),
            .I(N__26535));
    LocalMux I__2942 (
            .O(N__26538),
            .I(N__26532));
    LocalMux I__2941 (
            .O(N__26535),
            .I(N__26527));
    Span4Mux_v I__2940 (
            .O(N__26532),
            .I(N__26527));
    Odrv4 I__2939 (
            .O(N__26527),
            .I(data_out_frame_9_7));
    IoInMux I__2938 (
            .O(N__26524),
            .I(N__26521));
    LocalMux I__2937 (
            .O(N__26521),
            .I(N__26518));
    IoSpan4Mux I__2936 (
            .O(N__26518),
            .I(N__26514));
    InMux I__2935 (
            .O(N__26517),
            .I(N__26511));
    Span4Mux_s0_h I__2934 (
            .O(N__26514),
            .I(N__26508));
    LocalMux I__2933 (
            .O(N__26511),
            .I(N__26505));
    Span4Mux_s3_v I__2932 (
            .O(N__26508),
            .I(N__26500));
    Span4Mux_s3_v I__2931 (
            .O(N__26505),
            .I(N__26500));
    Sp12to4 I__2930 (
            .O(N__26500),
            .I(N__26497));
    Span12Mux_s10_h I__2929 (
            .O(N__26497),
            .I(N__26494));
    Span12Mux_v I__2928 (
            .O(N__26494),
            .I(N__26490));
    InMux I__2927 (
            .O(N__26493),
            .I(N__26487));
    Odrv12 I__2926 (
            .O(N__26490),
            .I(tx_o));
    LocalMux I__2925 (
            .O(N__26487),
            .I(tx_o));
    InMux I__2924 (
            .O(N__26482),
            .I(N__26478));
    InMux I__2923 (
            .O(N__26481),
            .I(N__26475));
    LocalMux I__2922 (
            .O(N__26478),
            .I(N__26472));
    LocalMux I__2921 (
            .O(N__26475),
            .I(N__26467));
    Span4Mux_h I__2920 (
            .O(N__26472),
            .I(N__26467));
    Odrv4 I__2919 (
            .O(N__26467),
            .I(\c0.data_out_frame_29__7__N_850 ));
    InMux I__2918 (
            .O(N__26464),
            .I(N__26461));
    LocalMux I__2917 (
            .O(N__26461),
            .I(N__26457));
    InMux I__2916 (
            .O(N__26460),
            .I(N__26454));
    Span4Mux_v I__2915 (
            .O(N__26457),
            .I(N__26451));
    LocalMux I__2914 (
            .O(N__26454),
            .I(data_out_frame_11_4));
    Odrv4 I__2913 (
            .O(N__26451),
            .I(data_out_frame_11_4));
    InMux I__2912 (
            .O(N__26446),
            .I(N__26443));
    LocalMux I__2911 (
            .O(N__26443),
            .I(N__26440));
    Span4Mux_h I__2910 (
            .O(N__26440),
            .I(N__26437));
    Odrv4 I__2909 (
            .O(N__26437),
            .I(\c0.n23881 ));
    InMux I__2908 (
            .O(N__26434),
            .I(N__26431));
    LocalMux I__2907 (
            .O(N__26431),
            .I(n2189));
    CascadeMux I__2906 (
            .O(N__26428),
            .I(N__26424));
    CascadeMux I__2905 (
            .O(N__26427),
            .I(N__26420));
    InMux I__2904 (
            .O(N__26424),
            .I(N__26414));
    InMux I__2903 (
            .O(N__26423),
            .I(N__26411));
    InMux I__2902 (
            .O(N__26420),
            .I(N__26408));
    InMux I__2901 (
            .O(N__26419),
            .I(N__26403));
    InMux I__2900 (
            .O(N__26418),
            .I(N__26403));
    InMux I__2899 (
            .O(N__26417),
            .I(N__26400));
    LocalMux I__2898 (
            .O(N__26414),
            .I(N__26397));
    LocalMux I__2897 (
            .O(N__26411),
            .I(N__26394));
    LocalMux I__2896 (
            .O(N__26408),
            .I(N__26389));
    LocalMux I__2895 (
            .O(N__26403),
            .I(N__26389));
    LocalMux I__2894 (
            .O(N__26400),
            .I(encoder1_position_16));
    Odrv4 I__2893 (
            .O(N__26397),
            .I(encoder1_position_16));
    Odrv4 I__2892 (
            .O(N__26394),
            .I(encoder1_position_16));
    Odrv4 I__2891 (
            .O(N__26389),
            .I(encoder1_position_16));
    InMux I__2890 (
            .O(N__26380),
            .I(N__26374));
    InMux I__2889 (
            .O(N__26379),
            .I(N__26374));
    LocalMux I__2888 (
            .O(N__26374),
            .I(data_out_frame_10_4));
    InMux I__2887 (
            .O(N__26371),
            .I(N__26368));
    LocalMux I__2886 (
            .O(N__26368),
            .I(N__26365));
    Span4Mux_v I__2885 (
            .O(N__26365),
            .I(N__26361));
    InMux I__2884 (
            .O(N__26364),
            .I(N__26358));
    Span4Mux_v I__2883 (
            .O(N__26361),
            .I(N__26355));
    LocalMux I__2882 (
            .O(N__26358),
            .I(data_out_frame_7_2));
    Odrv4 I__2881 (
            .O(N__26355),
            .I(data_out_frame_7_2));
    InMux I__2880 (
            .O(N__26350),
            .I(N__26347));
    LocalMux I__2879 (
            .O(N__26347),
            .I(n2188));
    InMux I__2878 (
            .O(N__26344),
            .I(N__26341));
    LocalMux I__2877 (
            .O(N__26341),
            .I(n2204));
    CascadeMux I__2876 (
            .O(N__26338),
            .I(\c0.n6_adj_4310_cascade_ ));
    InMux I__2875 (
            .O(N__26335),
            .I(N__26329));
    InMux I__2874 (
            .O(N__26334),
            .I(N__26329));
    LocalMux I__2873 (
            .O(N__26329),
            .I(\c0.n22037 ));
    InMux I__2872 (
            .O(N__26326),
            .I(N__26321));
    InMux I__2871 (
            .O(N__26325),
            .I(N__26315));
    InMux I__2870 (
            .O(N__26324),
            .I(N__26315));
    LocalMux I__2869 (
            .O(N__26321),
            .I(N__26312));
    InMux I__2868 (
            .O(N__26320),
            .I(N__26307));
    LocalMux I__2867 (
            .O(N__26315),
            .I(N__26304));
    Span4Mux_v I__2866 (
            .O(N__26312),
            .I(N__26301));
    InMux I__2865 (
            .O(N__26311),
            .I(N__26298));
    InMux I__2864 (
            .O(N__26310),
            .I(N__26295));
    LocalMux I__2863 (
            .O(N__26307),
            .I(N__26292));
    Span4Mux_h I__2862 (
            .O(N__26304),
            .I(N__26289));
    Odrv4 I__2861 (
            .O(N__26301),
            .I(encoder1_position_15));
    LocalMux I__2860 (
            .O(N__26298),
            .I(encoder1_position_15));
    LocalMux I__2859 (
            .O(N__26295),
            .I(encoder1_position_15));
    Odrv4 I__2858 (
            .O(N__26292),
            .I(encoder1_position_15));
    Odrv4 I__2857 (
            .O(N__26289),
            .I(encoder1_position_15));
    CascadeMux I__2856 (
            .O(N__26278),
            .I(N__26275));
    InMux I__2855 (
            .O(N__26275),
            .I(N__26269));
    InMux I__2854 (
            .O(N__26274),
            .I(N__26269));
    LocalMux I__2853 (
            .O(N__26269),
            .I(data_out_frame_12_7));
    InMux I__2852 (
            .O(N__26266),
            .I(N__26263));
    LocalMux I__2851 (
            .O(N__26263),
            .I(N__26260));
    Span4Mux_h I__2850 (
            .O(N__26260),
            .I(N__26257));
    Odrv4 I__2849 (
            .O(N__26257),
            .I(\c0.n11_adj_4360 ));
    InMux I__2848 (
            .O(N__26254),
            .I(N__26251));
    LocalMux I__2847 (
            .O(N__26251),
            .I(n2197));
    InMux I__2846 (
            .O(N__26248),
            .I(N__26245));
    LocalMux I__2845 (
            .O(N__26245),
            .I(N__26242));
    Odrv4 I__2844 (
            .O(N__26242),
            .I(\c0.n5_adj_4227 ));
    InMux I__2843 (
            .O(N__26239),
            .I(N__26233));
    InMux I__2842 (
            .O(N__26238),
            .I(N__26233));
    LocalMux I__2841 (
            .O(N__26233),
            .I(data_out_frame_7_4));
    InMux I__2840 (
            .O(N__26230),
            .I(N__26227));
    LocalMux I__2839 (
            .O(N__26227),
            .I(\c0.n22116 ));
    CascadeMux I__2838 (
            .O(N__26224),
            .I(N__26221));
    InMux I__2837 (
            .O(N__26221),
            .I(N__26218));
    LocalMux I__2836 (
            .O(N__26218),
            .I(N__26215));
    Odrv4 I__2835 (
            .O(N__26215),
            .I(\c0.n6_adj_4308 ));
    InMux I__2834 (
            .O(N__26212),
            .I(N__26208));
    InMux I__2833 (
            .O(N__26211),
            .I(N__26205));
    LocalMux I__2832 (
            .O(N__26208),
            .I(N__26200));
    LocalMux I__2831 (
            .O(N__26205),
            .I(N__26200));
    Odrv4 I__2830 (
            .O(N__26200),
            .I(data_out_frame_13_0));
    CascadeMux I__2829 (
            .O(N__26197),
            .I(N__26194));
    InMux I__2828 (
            .O(N__26194),
            .I(N__26191));
    LocalMux I__2827 (
            .O(N__26191),
            .I(N__26188));
    Span4Mux_v I__2826 (
            .O(N__26188),
            .I(N__26185));
    Span4Mux_v I__2825 (
            .O(N__26185),
            .I(N__26182));
    Odrv4 I__2824 (
            .O(N__26182),
            .I(\c0.n11_adj_4424 ));
    CascadeMux I__2823 (
            .O(N__26179),
            .I(\c0.n6_adj_4335_cascade_ ));
    CascadeMux I__2822 (
            .O(N__26176),
            .I(\c0.n21229_cascade_ ));
    InMux I__2821 (
            .O(N__26173),
            .I(N__26170));
    LocalMux I__2820 (
            .O(N__26170),
            .I(N__26167));
    Span4Mux_v I__2819 (
            .O(N__26167),
            .I(N__26164));
    Odrv4 I__2818 (
            .O(N__26164),
            .I(n2193));
    InMux I__2817 (
            .O(N__26161),
            .I(N__26158));
    LocalMux I__2816 (
            .O(N__26158),
            .I(N__26155));
    Odrv4 I__2815 (
            .O(N__26155),
            .I(\c0.n6_adj_4309 ));
    CascadeMux I__2814 (
            .O(N__26152),
            .I(N__26149));
    InMux I__2813 (
            .O(N__26149),
            .I(N__26145));
    InMux I__2812 (
            .O(N__26148),
            .I(N__26142));
    LocalMux I__2811 (
            .O(N__26145),
            .I(data_out_frame_29_2));
    LocalMux I__2810 (
            .O(N__26142),
            .I(data_out_frame_29_2));
    InMux I__2809 (
            .O(N__26137),
            .I(N__26134));
    LocalMux I__2808 (
            .O(N__26134),
            .I(N__26131));
    Span4Mux_v I__2807 (
            .O(N__26131),
            .I(N__26128));
    Odrv4 I__2806 (
            .O(N__26128),
            .I(n2196));
    CascadeMux I__2805 (
            .O(N__26125),
            .I(\c0.n13079_cascade_ ));
    CascadeMux I__2804 (
            .O(N__26122),
            .I(\c0.n21305_cascade_ ));
    InMux I__2803 (
            .O(N__26119),
            .I(N__26116));
    LocalMux I__2802 (
            .O(N__26116),
            .I(\c0.data_out_frame_28_2 ));
    InMux I__2801 (
            .O(N__26113),
            .I(N__26110));
    LocalMux I__2800 (
            .O(N__26110),
            .I(N__26107));
    Odrv4 I__2799 (
            .O(N__26107),
            .I(\c0.n6_adj_4515 ));
    CascadeMux I__2798 (
            .O(N__26104),
            .I(\c0.n12532_cascade_ ));
    CascadeMux I__2797 (
            .O(N__26101),
            .I(\c0.n22126_cascade_ ));
    InMux I__2796 (
            .O(N__26098),
            .I(N__26095));
    LocalMux I__2795 (
            .O(N__26095),
            .I(N__26092));
    Span4Mux_v I__2794 (
            .O(N__26092),
            .I(N__26089));
    Odrv4 I__2793 (
            .O(N__26089),
            .I(\c0.data_out_frame_28_4 ));
    InMux I__2792 (
            .O(N__26086),
            .I(N__26082));
    InMux I__2791 (
            .O(N__26085),
            .I(N__26079));
    LocalMux I__2790 (
            .O(N__26082),
            .I(N__26076));
    LocalMux I__2789 (
            .O(N__26079),
            .I(\quad_counter1.a_delay_counter_12 ));
    Odrv4 I__2788 (
            .O(N__26076),
            .I(\quad_counter1.a_delay_counter_12 ));
    InMux I__2787 (
            .O(N__26071),
            .I(N__26067));
    InMux I__2786 (
            .O(N__26070),
            .I(N__26064));
    LocalMux I__2785 (
            .O(N__26067),
            .I(\quad_counter1.a_delay_counter_13 ));
    LocalMux I__2784 (
            .O(N__26064),
            .I(\quad_counter1.a_delay_counter_13 ));
    CascadeMux I__2783 (
            .O(N__26059),
            .I(N__26055));
    InMux I__2782 (
            .O(N__26058),
            .I(N__26052));
    InMux I__2781 (
            .O(N__26055),
            .I(N__26049));
    LocalMux I__2780 (
            .O(N__26052),
            .I(\quad_counter1.a_delay_counter_9 ));
    LocalMux I__2779 (
            .O(N__26049),
            .I(\quad_counter1.a_delay_counter_9 ));
    InMux I__2778 (
            .O(N__26044),
            .I(N__26040));
    InMux I__2777 (
            .O(N__26043),
            .I(N__26037));
    LocalMux I__2776 (
            .O(N__26040),
            .I(\quad_counter1.a_delay_counter_6 ));
    LocalMux I__2775 (
            .O(N__26037),
            .I(\quad_counter1.a_delay_counter_6 ));
    InMux I__2774 (
            .O(N__26032),
            .I(N__26029));
    LocalMux I__2773 (
            .O(N__26029),
            .I(N__26026));
    Span4Mux_v I__2772 (
            .O(N__26026),
            .I(N__26023));
    Odrv4 I__2771 (
            .O(N__26023),
            .I(\quad_counter1.n26 ));
    SRMux I__2770 (
            .O(N__26020),
            .I(N__26017));
    LocalMux I__2769 (
            .O(N__26017),
            .I(N__26013));
    SRMux I__2768 (
            .O(N__26016),
            .I(N__26010));
    Span4Mux_v I__2767 (
            .O(N__26013),
            .I(N__26005));
    LocalMux I__2766 (
            .O(N__26010),
            .I(N__26005));
    Sp12to4 I__2765 (
            .O(N__26005),
            .I(N__26001));
    InMux I__2764 (
            .O(N__26004),
            .I(N__25998));
    Odrv12 I__2763 (
            .O(N__26001),
            .I(a_delay_counter_15__N_4124_adj_4547));
    LocalMux I__2762 (
            .O(N__25998),
            .I(a_delay_counter_15__N_4124_adj_4547));
    InMux I__2761 (
            .O(N__25993),
            .I(N__25988));
    InMux I__2760 (
            .O(N__25992),
            .I(N__25983));
    InMux I__2759 (
            .O(N__25991),
            .I(N__25983));
    LocalMux I__2758 (
            .O(N__25988),
            .I(N__25980));
    LocalMux I__2757 (
            .O(N__25983),
            .I(N__25977));
    Span4Mux_h I__2756 (
            .O(N__25980),
            .I(N__25974));
    Span4Mux_v I__2755 (
            .O(N__25977),
            .I(N__25971));
    Odrv4 I__2754 (
            .O(N__25974),
            .I(quadA_delayed_adj_4542));
    Odrv4 I__2753 (
            .O(N__25971),
            .I(quadA_delayed_adj_4542));
    InMux I__2752 (
            .O(N__25966),
            .I(N__25960));
    InMux I__2751 (
            .O(N__25965),
            .I(N__25960));
    LocalMux I__2750 (
            .O(N__25960),
            .I(N__25956));
    InMux I__2749 (
            .O(N__25959),
            .I(N__25953));
    Span4Mux_v I__2748 (
            .O(N__25956),
            .I(N__25950));
    LocalMux I__2747 (
            .O(N__25953),
            .I(N__25947));
    Span4Mux_h I__2746 (
            .O(N__25950),
            .I(N__25943));
    Span4Mux_v I__2745 (
            .O(N__25947),
            .I(N__25940));
    InMux I__2744 (
            .O(N__25946),
            .I(N__25937));
    Span4Mux_h I__2743 (
            .O(N__25943),
            .I(N__25934));
    Sp12to4 I__2742 (
            .O(N__25940),
            .I(N__25929));
    LocalMux I__2741 (
            .O(N__25937),
            .I(N__25929));
    Sp12to4 I__2740 (
            .O(N__25934),
            .I(N__25924));
    Span12Mux_h I__2739 (
            .O(N__25929),
            .I(N__25924));
    Odrv12 I__2738 (
            .O(N__25924),
            .I(PIN_12_c));
    CascadeMux I__2737 (
            .O(N__25921),
            .I(a_delay_counter_15__N_4124_adj_4547_cascade_));
    InMux I__2736 (
            .O(N__25918),
            .I(N__25915));
    LocalMux I__2735 (
            .O(N__25915),
            .I(N__25912));
    Span4Mux_h I__2734 (
            .O(N__25912),
            .I(N__25909));
    Odrv4 I__2733 (
            .O(N__25909),
            .I(n9818));
    CEMux I__2732 (
            .O(N__25906),
            .I(N__25901));
    CEMux I__2731 (
            .O(N__25905),
            .I(N__25898));
    InMux I__2730 (
            .O(N__25904),
            .I(N__25895));
    LocalMux I__2729 (
            .O(N__25901),
            .I(n14228));
    LocalMux I__2728 (
            .O(N__25898),
            .I(n14228));
    LocalMux I__2727 (
            .O(N__25895),
            .I(n14228));
    InMux I__2726 (
            .O(N__25888),
            .I(\quad_counter0.n19502 ));
    InMux I__2725 (
            .O(N__25885),
            .I(N__25882));
    LocalMux I__2724 (
            .O(N__25882),
            .I(\c0.n24_adj_4502 ));
    CascadeMux I__2723 (
            .O(N__25879),
            .I(\c0.n18_adj_4414_cascade_ ));
    InMux I__2722 (
            .O(N__25876),
            .I(N__25873));
    LocalMux I__2721 (
            .O(N__25873),
            .I(\c0.n13360 ));
    CascadeMux I__2720 (
            .O(N__25870),
            .I(\c0.n23550_cascade_ ));
    CascadeMux I__2719 (
            .O(N__25867),
            .I(\c0.n22_adj_4503_cascade_ ));
    InMux I__2718 (
            .O(N__25864),
            .I(N__25861));
    LocalMux I__2717 (
            .O(N__25861),
            .I(\c0.n26_adj_4504 ));
    InMux I__2716 (
            .O(N__25858),
            .I(N__25855));
    LocalMux I__2715 (
            .O(N__25855),
            .I(N__25852));
    Span4Mux_h I__2714 (
            .O(N__25852),
            .I(N__25849));
    Span4Mux_v I__2713 (
            .O(N__25849),
            .I(N__25846));
    Span4Mux_v I__2712 (
            .O(N__25846),
            .I(N__25843));
    Odrv4 I__2711 (
            .O(N__25843),
            .I(\c0.n26_adj_4517 ));
    InMux I__2710 (
            .O(N__25840),
            .I(\quad_counter0.n19493 ));
    InMux I__2709 (
            .O(N__25837),
            .I(\quad_counter0.n19494 ));
    InMux I__2708 (
            .O(N__25834),
            .I(bfn_10_25_0_));
    InMux I__2707 (
            .O(N__25831),
            .I(\quad_counter0.n19496 ));
    InMux I__2706 (
            .O(N__25828),
            .I(\quad_counter0.n19497 ));
    InMux I__2705 (
            .O(N__25825),
            .I(\quad_counter0.n19498 ));
    InMux I__2704 (
            .O(N__25822),
            .I(\quad_counter0.n19499 ));
    InMux I__2703 (
            .O(N__25819),
            .I(\quad_counter0.n19500 ));
    InMux I__2702 (
            .O(N__25816),
            .I(\quad_counter0.n19501 ));
    InMux I__2701 (
            .O(N__25813),
            .I(\quad_counter0.n19485 ));
    InMux I__2700 (
            .O(N__25810),
            .I(\quad_counter0.n19486 ));
    InMux I__2699 (
            .O(N__25807),
            .I(\quad_counter0.n19487 ));
    CEMux I__2698 (
            .O(N__25804),
            .I(N__25800));
    CEMux I__2697 (
            .O(N__25803),
            .I(N__25797));
    LocalMux I__2696 (
            .O(N__25800),
            .I(N__25793));
    LocalMux I__2695 (
            .O(N__25797),
            .I(N__25790));
    InMux I__2694 (
            .O(N__25796),
            .I(N__25787));
    Odrv4 I__2693 (
            .O(N__25793),
            .I(n14198));
    Odrv4 I__2692 (
            .O(N__25790),
            .I(n14198));
    LocalMux I__2691 (
            .O(N__25787),
            .I(n14198));
    SRMux I__2690 (
            .O(N__25780),
            .I(N__25777));
    LocalMux I__2689 (
            .O(N__25777),
            .I(N__25773));
    SRMux I__2688 (
            .O(N__25776),
            .I(N__25770));
    Span4Mux_h I__2687 (
            .O(N__25773),
            .I(N__25766));
    LocalMux I__2686 (
            .O(N__25770),
            .I(N__25763));
    InMux I__2685 (
            .O(N__25769),
            .I(N__25760));
    Odrv4 I__2684 (
            .O(N__25766),
            .I(b_delay_counter_15__N_4141));
    Odrv4 I__2683 (
            .O(N__25763),
            .I(b_delay_counter_15__N_4141));
    LocalMux I__2682 (
            .O(N__25760),
            .I(b_delay_counter_15__N_4141));
    InMux I__2681 (
            .O(N__25753),
            .I(bfn_10_24_0_));
    InMux I__2680 (
            .O(N__25750),
            .I(\quad_counter0.n19488 ));
    InMux I__2679 (
            .O(N__25747),
            .I(\quad_counter0.n19489 ));
    InMux I__2678 (
            .O(N__25744),
            .I(\quad_counter0.n19490 ));
    InMux I__2677 (
            .O(N__25741),
            .I(\quad_counter0.n19491 ));
    InMux I__2676 (
            .O(N__25738),
            .I(\quad_counter0.n19492 ));
    InMux I__2675 (
            .O(N__25735),
            .I(\quad_counter0.n19476 ));
    InMux I__2674 (
            .O(N__25732),
            .I(\quad_counter0.n19477 ));
    InMux I__2673 (
            .O(N__25729),
            .I(\quad_counter0.n19478 ));
    InMux I__2672 (
            .O(N__25726),
            .I(\quad_counter0.n19479 ));
    InMux I__2671 (
            .O(N__25723),
            .I(bfn_10_23_0_));
    InMux I__2670 (
            .O(N__25720),
            .I(\quad_counter0.n19481 ));
    InMux I__2669 (
            .O(N__25717),
            .I(\quad_counter0.n19482 ));
    InMux I__2668 (
            .O(N__25714),
            .I(\quad_counter0.n19483 ));
    InMux I__2667 (
            .O(N__25711),
            .I(\quad_counter0.n19484 ));
    CascadeMux I__2666 (
            .O(N__25708),
            .I(n24100_cascade_));
    InMux I__2665 (
            .O(N__25705),
            .I(N__25702));
    LocalMux I__2664 (
            .O(N__25702),
            .I(n16706));
    CascadeMux I__2663 (
            .O(N__25699),
            .I(\c0.tx.n23985_cascade_ ));
    CascadeMux I__2662 (
            .O(N__25696),
            .I(\c0.tx.n31_adj_4216_cascade_ ));
    InMux I__2661 (
            .O(N__25693),
            .I(N__25690));
    LocalMux I__2660 (
            .O(N__25690),
            .I(n187));
    InMux I__2659 (
            .O(N__25687),
            .I(bfn_10_22_0_));
    InMux I__2658 (
            .O(N__25684),
            .I(\quad_counter0.n19473 ));
    InMux I__2657 (
            .O(N__25681),
            .I(\quad_counter0.n19474 ));
    InMux I__2656 (
            .O(N__25678),
            .I(\quad_counter0.n19475 ));
    InMux I__2655 (
            .O(N__25675),
            .I(N__25672));
    LocalMux I__2654 (
            .O(N__25672),
            .I(N__25669));
    Span4Mux_h I__2653 (
            .O(N__25669),
            .I(N__25666));
    Span4Mux_v I__2652 (
            .O(N__25666),
            .I(N__25663));
    Odrv4 I__2651 (
            .O(N__25663),
            .I(n10_adj_4536));
    InMux I__2650 (
            .O(N__25660),
            .I(N__25657));
    LocalMux I__2649 (
            .O(N__25657),
            .I(\c0.n5_adj_4422 ));
    CascadeMux I__2648 (
            .O(N__25654),
            .I(N__25651));
    InMux I__2647 (
            .O(N__25651),
            .I(N__25648));
    LocalMux I__2646 (
            .O(N__25648),
            .I(\c0.n24059 ));
    CascadeMux I__2645 (
            .O(N__25645),
            .I(\c0.n23850_cascade_ ));
    CascadeMux I__2644 (
            .O(N__25642),
            .I(n23852_cascade_));
    CascadeMux I__2643 (
            .O(N__25639),
            .I(N__25630));
    InMux I__2642 (
            .O(N__25638),
            .I(N__25627));
    InMux I__2641 (
            .O(N__25637),
            .I(N__25623));
    InMux I__2640 (
            .O(N__25636),
            .I(N__25620));
    InMux I__2639 (
            .O(N__25635),
            .I(N__25617));
    InMux I__2638 (
            .O(N__25634),
            .I(N__25614));
    InMux I__2637 (
            .O(N__25633),
            .I(N__25611));
    InMux I__2636 (
            .O(N__25630),
            .I(N__25608));
    LocalMux I__2635 (
            .O(N__25627),
            .I(N__25604));
    InMux I__2634 (
            .O(N__25626),
            .I(N__25601));
    LocalMux I__2633 (
            .O(N__25623),
            .I(N__25596));
    LocalMux I__2632 (
            .O(N__25620),
            .I(N__25596));
    LocalMux I__2631 (
            .O(N__25617),
            .I(N__25591));
    LocalMux I__2630 (
            .O(N__25614),
            .I(N__25591));
    LocalMux I__2629 (
            .O(N__25611),
            .I(N__25586));
    LocalMux I__2628 (
            .O(N__25608),
            .I(N__25583));
    InMux I__2627 (
            .O(N__25607),
            .I(N__25580));
    Span4Mux_h I__2626 (
            .O(N__25604),
            .I(N__25577));
    LocalMux I__2625 (
            .O(N__25601),
            .I(N__25570));
    Span4Mux_v I__2624 (
            .O(N__25596),
            .I(N__25570));
    Span4Mux_v I__2623 (
            .O(N__25591),
            .I(N__25570));
    InMux I__2622 (
            .O(N__25590),
            .I(N__25565));
    InMux I__2621 (
            .O(N__25589),
            .I(N__25565));
    Span4Mux_v I__2620 (
            .O(N__25586),
            .I(N__25558));
    Span4Mux_v I__2619 (
            .O(N__25583),
            .I(N__25558));
    LocalMux I__2618 (
            .O(N__25580),
            .I(N__25558));
    Odrv4 I__2617 (
            .O(N__25577),
            .I(byte_transmit_counter_3));
    Odrv4 I__2616 (
            .O(N__25570),
            .I(byte_transmit_counter_3));
    LocalMux I__2615 (
            .O(N__25565),
            .I(byte_transmit_counter_3));
    Odrv4 I__2614 (
            .O(N__25558),
            .I(byte_transmit_counter_3));
    CascadeMux I__2613 (
            .O(N__25549),
            .I(n10_adj_4537_cascade_));
    InMux I__2612 (
            .O(N__25546),
            .I(N__25543));
    LocalMux I__2611 (
            .O(N__25543),
            .I(n24110));
    CascadeMux I__2610 (
            .O(N__25540),
            .I(N__25536));
    InMux I__2609 (
            .O(N__25539),
            .I(N__25531));
    InMux I__2608 (
            .O(N__25536),
            .I(N__25531));
    LocalMux I__2607 (
            .O(N__25531),
            .I(r_Tx_Data_0));
    InMux I__2606 (
            .O(N__25528),
            .I(N__25525));
    LocalMux I__2605 (
            .O(N__25525),
            .I(n24195));
    InMux I__2604 (
            .O(N__25522),
            .I(N__25518));
    InMux I__2603 (
            .O(N__25521),
            .I(N__25515));
    LocalMux I__2602 (
            .O(N__25518),
            .I(N__25512));
    LocalMux I__2601 (
            .O(N__25515),
            .I(r_Tx_Data_5));
    Odrv12 I__2600 (
            .O(N__25512),
            .I(r_Tx_Data_5));
    InMux I__2599 (
            .O(N__25507),
            .I(N__25504));
    LocalMux I__2598 (
            .O(N__25504),
            .I(N__25500));
    InMux I__2597 (
            .O(N__25503),
            .I(N__25497));
    Span4Mux_v I__2596 (
            .O(N__25500),
            .I(N__25494));
    LocalMux I__2595 (
            .O(N__25497),
            .I(r_Tx_Data_4));
    Odrv4 I__2594 (
            .O(N__25494),
            .I(r_Tx_Data_4));
    InMux I__2593 (
            .O(N__25489),
            .I(N__25486));
    LocalMux I__2592 (
            .O(N__25486),
            .I(n10_adj_4533));
    InMux I__2591 (
            .O(N__25483),
            .I(N__25479));
    InMux I__2590 (
            .O(N__25482),
            .I(N__25476));
    LocalMux I__2589 (
            .O(N__25479),
            .I(data_out_frame_9_2));
    LocalMux I__2588 (
            .O(N__25476),
            .I(data_out_frame_9_2));
    CascadeMux I__2587 (
            .O(N__25471),
            .I(\c0.n24180_cascade_ ));
    InMux I__2586 (
            .O(N__25468),
            .I(N__25465));
    LocalMux I__2585 (
            .O(N__25465),
            .I(n24106));
    CascadeMux I__2584 (
            .O(N__25462),
            .I(N__25459));
    InMux I__2583 (
            .O(N__25459),
            .I(N__25453));
    InMux I__2582 (
            .O(N__25458),
            .I(N__25453));
    LocalMux I__2581 (
            .O(N__25453),
            .I(data_out_frame_7_0));
    InMux I__2580 (
            .O(N__25450),
            .I(N__25444));
    InMux I__2579 (
            .O(N__25449),
            .I(N__25444));
    LocalMux I__2578 (
            .O(N__25444),
            .I(data_out_frame_6_0));
    InMux I__2577 (
            .O(N__25441),
            .I(bfn_10_17_0_));
    InMux I__2576 (
            .O(N__25438),
            .I(N__25435));
    LocalMux I__2575 (
            .O(N__25435),
            .I(N__25432));
    Odrv4 I__2574 (
            .O(N__25432),
            .I(n2174));
    InMux I__2573 (
            .O(N__25429),
            .I(N__25426));
    LocalMux I__2572 (
            .O(N__25426),
            .I(N__25422));
    InMux I__2571 (
            .O(N__25425),
            .I(N__25419));
    Span4Mux_h I__2570 (
            .O(N__25422),
            .I(N__25416));
    LocalMux I__2569 (
            .O(N__25419),
            .I(data_out_frame_0_4));
    Odrv4 I__2568 (
            .O(N__25416),
            .I(data_out_frame_0_4));
    InMux I__2567 (
            .O(N__25411),
            .I(N__25407));
    InMux I__2566 (
            .O(N__25410),
            .I(N__25404));
    LocalMux I__2565 (
            .O(N__25407),
            .I(data_out_frame_13_5));
    LocalMux I__2564 (
            .O(N__25404),
            .I(data_out_frame_13_5));
    InMux I__2563 (
            .O(N__25399),
            .I(N__25393));
    InMux I__2562 (
            .O(N__25398),
            .I(N__25393));
    LocalMux I__2561 (
            .O(N__25393),
            .I(data_out_frame_9_3));
    InMux I__2560 (
            .O(N__25390),
            .I(N__25387));
    LocalMux I__2559 (
            .O(N__25387),
            .I(\c0.n24171 ));
    InMux I__2558 (
            .O(N__25384),
            .I(N__25381));
    LocalMux I__2557 (
            .O(N__25381),
            .I(\c0.n24174 ));
    InMux I__2556 (
            .O(N__25378),
            .I(N__25375));
    LocalMux I__2555 (
            .O(N__25375),
            .I(\c0.n23856 ));
    InMux I__2554 (
            .O(N__25372),
            .I(N__25369));
    LocalMux I__2553 (
            .O(N__25369),
            .I(N__25366));
    Odrv4 I__2552 (
            .O(N__25366),
            .I(n24108));
    CascadeMux I__2551 (
            .O(N__25363),
            .I(n23858_cascade_));
    InMux I__2550 (
            .O(N__25360),
            .I(bfn_10_16_0_));
    InMux I__2549 (
            .O(N__25357),
            .I(\quad_counter1.n19572 ));
    InMux I__2548 (
            .O(N__25354),
            .I(\quad_counter1.n19573 ));
    InMux I__2547 (
            .O(N__25351),
            .I(N__25348));
    LocalMux I__2546 (
            .O(N__25348),
            .I(N__25345));
    Odrv12 I__2545 (
            .O(N__25345),
            .I(n2179));
    InMux I__2544 (
            .O(N__25342),
            .I(\quad_counter1.n19574 ));
    InMux I__2543 (
            .O(N__25339),
            .I(\quad_counter1.n19575 ));
    InMux I__2542 (
            .O(N__25336),
            .I(N__25333));
    LocalMux I__2541 (
            .O(N__25333),
            .I(n2177));
    InMux I__2540 (
            .O(N__25330),
            .I(\quad_counter1.n19576 ));
    InMux I__2539 (
            .O(N__25327),
            .I(\quad_counter1.n19577 ));
    InMux I__2538 (
            .O(N__25324),
            .I(\quad_counter1.n19578 ));
    CascadeMux I__2537 (
            .O(N__25321),
            .I(N__25303));
    CascadeMux I__2536 (
            .O(N__25320),
            .I(N__25299));
    CascadeMux I__2535 (
            .O(N__25319),
            .I(N__25295));
    CascadeMux I__2534 (
            .O(N__25318),
            .I(N__25290));
    CascadeMux I__2533 (
            .O(N__25317),
            .I(N__25286));
    CascadeMux I__2532 (
            .O(N__25316),
            .I(N__25282));
    CascadeMux I__2531 (
            .O(N__25315),
            .I(N__25278));
    CascadeMux I__2530 (
            .O(N__25314),
            .I(N__25275));
    CascadeMux I__2529 (
            .O(N__25313),
            .I(N__25271));
    CascadeMux I__2528 (
            .O(N__25312),
            .I(N__25267));
    CascadeMux I__2527 (
            .O(N__25311),
            .I(N__25263));
    CascadeMux I__2526 (
            .O(N__25310),
            .I(N__25258));
    CascadeMux I__2525 (
            .O(N__25309),
            .I(N__25255));
    CascadeMux I__2524 (
            .O(N__25308),
            .I(N__25252));
    CascadeMux I__2523 (
            .O(N__25307),
            .I(N__25247));
    InMux I__2522 (
            .O(N__25306),
            .I(N__25243));
    InMux I__2521 (
            .O(N__25303),
            .I(N__25230));
    InMux I__2520 (
            .O(N__25302),
            .I(N__25230));
    InMux I__2519 (
            .O(N__25299),
            .I(N__25230));
    InMux I__2518 (
            .O(N__25298),
            .I(N__25230));
    InMux I__2517 (
            .O(N__25295),
            .I(N__25230));
    InMux I__2516 (
            .O(N__25294),
            .I(N__25230));
    InMux I__2515 (
            .O(N__25293),
            .I(N__25213));
    InMux I__2514 (
            .O(N__25290),
            .I(N__25213));
    InMux I__2513 (
            .O(N__25289),
            .I(N__25213));
    InMux I__2512 (
            .O(N__25286),
            .I(N__25213));
    InMux I__2511 (
            .O(N__25285),
            .I(N__25213));
    InMux I__2510 (
            .O(N__25282),
            .I(N__25213));
    InMux I__2509 (
            .O(N__25281),
            .I(N__25213));
    InMux I__2508 (
            .O(N__25278),
            .I(N__25213));
    InMux I__2507 (
            .O(N__25275),
            .I(N__25196));
    InMux I__2506 (
            .O(N__25274),
            .I(N__25196));
    InMux I__2505 (
            .O(N__25271),
            .I(N__25196));
    InMux I__2504 (
            .O(N__25270),
            .I(N__25196));
    InMux I__2503 (
            .O(N__25267),
            .I(N__25196));
    InMux I__2502 (
            .O(N__25266),
            .I(N__25196));
    InMux I__2501 (
            .O(N__25263),
            .I(N__25196));
    InMux I__2500 (
            .O(N__25262),
            .I(N__25196));
    InMux I__2499 (
            .O(N__25261),
            .I(N__25187));
    InMux I__2498 (
            .O(N__25258),
            .I(N__25187));
    InMux I__2497 (
            .O(N__25255),
            .I(N__25187));
    InMux I__2496 (
            .O(N__25252),
            .I(N__25187));
    CascadeMux I__2495 (
            .O(N__25251),
            .I(N__25183));
    CascadeMux I__2494 (
            .O(N__25250),
            .I(N__25180));
    InMux I__2493 (
            .O(N__25247),
            .I(N__25174));
    InMux I__2492 (
            .O(N__25246),
            .I(N__25174));
    LocalMux I__2491 (
            .O(N__25243),
            .I(N__25165));
    LocalMux I__2490 (
            .O(N__25230),
            .I(N__25165));
    LocalMux I__2489 (
            .O(N__25213),
            .I(N__25165));
    LocalMux I__2488 (
            .O(N__25196),
            .I(N__25165));
    LocalMux I__2487 (
            .O(N__25187),
            .I(N__25162));
    InMux I__2486 (
            .O(N__25186),
            .I(N__25153));
    InMux I__2485 (
            .O(N__25183),
            .I(N__25153));
    InMux I__2484 (
            .O(N__25180),
            .I(N__25153));
    InMux I__2483 (
            .O(N__25179),
            .I(N__25153));
    LocalMux I__2482 (
            .O(N__25174),
            .I(N__25150));
    Span4Mux_v I__2481 (
            .O(N__25165),
            .I(N__25143));
    Span4Mux_h I__2480 (
            .O(N__25162),
            .I(N__25143));
    LocalMux I__2479 (
            .O(N__25153),
            .I(N__25143));
    Span4Mux_v I__2478 (
            .O(N__25150),
            .I(N__25140));
    Span4Mux_v I__2477 (
            .O(N__25143),
            .I(N__25137));
    Odrv4 I__2476 (
            .O(N__25140),
            .I(\quad_counter1.n2140 ));
    Odrv4 I__2475 (
            .O(N__25137),
            .I(\quad_counter1.n2140 ));
    InMux I__2474 (
            .O(N__25132),
            .I(N__25129));
    LocalMux I__2473 (
            .O(N__25129),
            .I(N__25126));
    Odrv12 I__2472 (
            .O(N__25126),
            .I(n2191));
    InMux I__2471 (
            .O(N__25123),
            .I(\quad_counter1.n19562 ));
    InMux I__2470 (
            .O(N__25120),
            .I(N__25117));
    LocalMux I__2469 (
            .O(N__25117),
            .I(n2190));
    InMux I__2468 (
            .O(N__25114),
            .I(bfn_10_15_0_));
    InMux I__2467 (
            .O(N__25111),
            .I(\quad_counter1.n19564 ));
    InMux I__2466 (
            .O(N__25108),
            .I(\quad_counter1.n19565 ));
    InMux I__2465 (
            .O(N__25105),
            .I(N__25102));
    LocalMux I__2464 (
            .O(N__25102),
            .I(N__25099));
    Odrv4 I__2463 (
            .O(N__25099),
            .I(n2187));
    InMux I__2462 (
            .O(N__25096),
            .I(\quad_counter1.n19566 ));
    InMux I__2461 (
            .O(N__25093),
            .I(\quad_counter1.n19567 ));
    InMux I__2460 (
            .O(N__25090),
            .I(\quad_counter1.n19568 ));
    InMux I__2459 (
            .O(N__25087),
            .I(\quad_counter1.n19569 ));
    InMux I__2458 (
            .O(N__25084),
            .I(N__25081));
    LocalMux I__2457 (
            .O(N__25081),
            .I(N__25078));
    Odrv12 I__2456 (
            .O(N__25078),
            .I(n2183));
    InMux I__2455 (
            .O(N__25075),
            .I(\quad_counter1.n19570 ));
    InMux I__2454 (
            .O(N__25072),
            .I(N__25069));
    LocalMux I__2453 (
            .O(N__25069),
            .I(N__25066));
    Odrv4 I__2452 (
            .O(N__25066),
            .I(n2200));
    InMux I__2451 (
            .O(N__25063),
            .I(\quad_counter1.n19553 ));
    InMux I__2450 (
            .O(N__25060),
            .I(N__25057));
    LocalMux I__2449 (
            .O(N__25057),
            .I(n2199));
    InMux I__2448 (
            .O(N__25054),
            .I(\quad_counter1.n19554 ));
    InMux I__2447 (
            .O(N__25051),
            .I(bfn_10_14_0_));
    InMux I__2446 (
            .O(N__25048),
            .I(\quad_counter1.n19556 ));
    InMux I__2445 (
            .O(N__25045),
            .I(\quad_counter1.n19557 ));
    InMux I__2444 (
            .O(N__25042),
            .I(\quad_counter1.n19558 ));
    InMux I__2443 (
            .O(N__25039),
            .I(\quad_counter1.n19559 ));
    InMux I__2442 (
            .O(N__25036),
            .I(\quad_counter1.n19560 ));
    InMux I__2441 (
            .O(N__25033),
            .I(\quad_counter1.n19561 ));
    CascadeMux I__2440 (
            .O(N__25030),
            .I(\c0.n22048_cascade_ ));
    CascadeMux I__2439 (
            .O(N__25027),
            .I(N__25022));
    InMux I__2438 (
            .O(N__25026),
            .I(N__25018));
    InMux I__2437 (
            .O(N__25025),
            .I(N__25011));
    InMux I__2436 (
            .O(N__25022),
            .I(N__25011));
    InMux I__2435 (
            .O(N__25021),
            .I(N__25011));
    LocalMux I__2434 (
            .O(N__25018),
            .I(encoder1_position_0));
    LocalMux I__2433 (
            .O(N__25011),
            .I(encoder1_position_0));
    CascadeMux I__2432 (
            .O(N__25006),
            .I(N__25003));
    InMux I__2431 (
            .O(N__25003),
            .I(N__25000));
    LocalMux I__2430 (
            .O(N__25000),
            .I(N__24997));
    Odrv4 I__2429 (
            .O(N__24997),
            .I(\quad_counter1.count_direction ));
    InMux I__2428 (
            .O(N__24994),
            .I(N__24991));
    LocalMux I__2427 (
            .O(N__24991),
            .I(n2205));
    InMux I__2426 (
            .O(N__24988),
            .I(\quad_counter1.n19548 ));
    InMux I__2425 (
            .O(N__24985),
            .I(\quad_counter1.n19549 ));
    InMux I__2424 (
            .O(N__24982),
            .I(N__24979));
    LocalMux I__2423 (
            .O(N__24979),
            .I(N__24976));
    Odrv4 I__2422 (
            .O(N__24976),
            .I(n2203));
    InMux I__2421 (
            .O(N__24973),
            .I(\quad_counter1.n19550 ));
    InMux I__2420 (
            .O(N__24970),
            .I(N__24967));
    LocalMux I__2419 (
            .O(N__24967),
            .I(N__24964));
    Odrv4 I__2418 (
            .O(N__24964),
            .I(n2202));
    InMux I__2417 (
            .O(N__24961),
            .I(\quad_counter1.n19551 ));
    InMux I__2416 (
            .O(N__24958),
            .I(\quad_counter1.n19552 ));
    CascadeMux I__2415 (
            .O(N__24955),
            .I(N__24950));
    InMux I__2414 (
            .O(N__24954),
            .I(N__24947));
    InMux I__2413 (
            .O(N__24953),
            .I(N__24942));
    InMux I__2412 (
            .O(N__24950),
            .I(N__24942));
    LocalMux I__2411 (
            .O(N__24947),
            .I(N__24939));
    LocalMux I__2410 (
            .O(N__24942),
            .I(N__24934));
    Span4Mux_h I__2409 (
            .O(N__24939),
            .I(N__24931));
    InMux I__2408 (
            .O(N__24938),
            .I(N__24926));
    InMux I__2407 (
            .O(N__24937),
            .I(N__24926));
    Odrv12 I__2406 (
            .O(N__24934),
            .I(A_filtered_adj_4538));
    Odrv4 I__2405 (
            .O(N__24931),
            .I(A_filtered_adj_4538));
    LocalMux I__2404 (
            .O(N__24926),
            .I(A_filtered_adj_4538));
    InMux I__2403 (
            .O(N__24919),
            .I(N__24915));
    InMux I__2402 (
            .O(N__24918),
            .I(N__24912));
    LocalMux I__2401 (
            .O(N__24915),
            .I(N__24906));
    LocalMux I__2400 (
            .O(N__24912),
            .I(N__24906));
    InMux I__2399 (
            .O(N__24911),
            .I(N__24903));
    Odrv4 I__2398 (
            .O(N__24906),
            .I(\quad_counter1.B_delayed ));
    LocalMux I__2397 (
            .O(N__24903),
            .I(\quad_counter1.B_delayed ));
    InMux I__2396 (
            .O(N__24898),
            .I(N__24895));
    LocalMux I__2395 (
            .O(N__24895),
            .I(N__24892));
    Odrv4 I__2394 (
            .O(N__24892),
            .I(n39_adj_4545));
    InMux I__2393 (
            .O(N__24889),
            .I(N__24884));
    CascadeMux I__2392 (
            .O(N__24888),
            .I(N__24881));
    InMux I__2391 (
            .O(N__24887),
            .I(N__24878));
    LocalMux I__2390 (
            .O(N__24884),
            .I(N__24875));
    InMux I__2389 (
            .O(N__24881),
            .I(N__24872));
    LocalMux I__2388 (
            .O(N__24878),
            .I(N__24869));
    Span4Mux_h I__2387 (
            .O(N__24875),
            .I(N__24866));
    LocalMux I__2386 (
            .O(N__24872),
            .I(a_delay_counter_0_adj_4540));
    Odrv12 I__2385 (
            .O(N__24869),
            .I(a_delay_counter_0_adj_4540));
    Odrv4 I__2384 (
            .O(N__24866),
            .I(a_delay_counter_0_adj_4540));
    CascadeMux I__2383 (
            .O(N__24859),
            .I(N__24855));
    InMux I__2382 (
            .O(N__24858),
            .I(N__24852));
    InMux I__2381 (
            .O(N__24855),
            .I(N__24849));
    LocalMux I__2380 (
            .O(N__24852),
            .I(\quad_counter1.a_delay_counter_10 ));
    LocalMux I__2379 (
            .O(N__24849),
            .I(\quad_counter1.a_delay_counter_10 ));
    InMux I__2378 (
            .O(N__24844),
            .I(\quad_counter1.n19527 ));
    InMux I__2377 (
            .O(N__24841),
            .I(N__24837));
    InMux I__2376 (
            .O(N__24840),
            .I(N__24834));
    LocalMux I__2375 (
            .O(N__24837),
            .I(\quad_counter1.a_delay_counter_11 ));
    LocalMux I__2374 (
            .O(N__24834),
            .I(\quad_counter1.a_delay_counter_11 ));
    InMux I__2373 (
            .O(N__24829),
            .I(\quad_counter1.n19528 ));
    InMux I__2372 (
            .O(N__24826),
            .I(\quad_counter1.n19529 ));
    InMux I__2371 (
            .O(N__24823),
            .I(\quad_counter1.n19530 ));
    InMux I__2370 (
            .O(N__24820),
            .I(N__24816));
    InMux I__2369 (
            .O(N__24819),
            .I(N__24813));
    LocalMux I__2368 (
            .O(N__24816),
            .I(\quad_counter1.a_delay_counter_14 ));
    LocalMux I__2367 (
            .O(N__24813),
            .I(\quad_counter1.a_delay_counter_14 ));
    InMux I__2366 (
            .O(N__24808),
            .I(\quad_counter1.n19531 ));
    InMux I__2365 (
            .O(N__24805),
            .I(\quad_counter1.n19532 ));
    InMux I__2364 (
            .O(N__24802),
            .I(N__24798));
    InMux I__2363 (
            .O(N__24801),
            .I(N__24795));
    LocalMux I__2362 (
            .O(N__24798),
            .I(\quad_counter1.a_delay_counter_15 ));
    LocalMux I__2361 (
            .O(N__24795),
            .I(\quad_counter1.a_delay_counter_15 ));
    CascadeMux I__2360 (
            .O(N__24790),
            .I(N__24786));
    CascadeMux I__2359 (
            .O(N__24789),
            .I(N__24783));
    InMux I__2358 (
            .O(N__24786),
            .I(N__24780));
    InMux I__2357 (
            .O(N__24783),
            .I(N__24777));
    LocalMux I__2356 (
            .O(N__24780),
            .I(N__24774));
    LocalMux I__2355 (
            .O(N__24777),
            .I(data_out_frame_11_6));
    Odrv4 I__2354 (
            .O(N__24774),
            .I(data_out_frame_11_6));
    InMux I__2353 (
            .O(N__24769),
            .I(N__24765));
    InMux I__2352 (
            .O(N__24768),
            .I(N__24762));
    LocalMux I__2351 (
            .O(N__24765),
            .I(N__24757));
    LocalMux I__2350 (
            .O(N__24762),
            .I(N__24757));
    Odrv4 I__2349 (
            .O(N__24757),
            .I(\quad_counter1.a_delay_counter_1 ));
    InMux I__2348 (
            .O(N__24754),
            .I(\quad_counter1.n19518 ));
    CascadeMux I__2347 (
            .O(N__24751),
            .I(N__24747));
    InMux I__2346 (
            .O(N__24750),
            .I(N__24744));
    InMux I__2345 (
            .O(N__24747),
            .I(N__24741));
    LocalMux I__2344 (
            .O(N__24744),
            .I(\quad_counter1.a_delay_counter_2 ));
    LocalMux I__2343 (
            .O(N__24741),
            .I(\quad_counter1.a_delay_counter_2 ));
    InMux I__2342 (
            .O(N__24736),
            .I(\quad_counter1.n19519 ));
    InMux I__2341 (
            .O(N__24733),
            .I(N__24729));
    InMux I__2340 (
            .O(N__24732),
            .I(N__24726));
    LocalMux I__2339 (
            .O(N__24729),
            .I(\quad_counter1.a_delay_counter_3 ));
    LocalMux I__2338 (
            .O(N__24726),
            .I(\quad_counter1.a_delay_counter_3 ));
    InMux I__2337 (
            .O(N__24721),
            .I(\quad_counter1.n19520 ));
    CascadeMux I__2336 (
            .O(N__24718),
            .I(N__24714));
    InMux I__2335 (
            .O(N__24717),
            .I(N__24711));
    InMux I__2334 (
            .O(N__24714),
            .I(N__24708));
    LocalMux I__2333 (
            .O(N__24711),
            .I(\quad_counter1.a_delay_counter_4 ));
    LocalMux I__2332 (
            .O(N__24708),
            .I(\quad_counter1.a_delay_counter_4 ));
    InMux I__2331 (
            .O(N__24703),
            .I(\quad_counter1.n19521 ));
    InMux I__2330 (
            .O(N__24700),
            .I(N__24696));
    InMux I__2329 (
            .O(N__24699),
            .I(N__24693));
    LocalMux I__2328 (
            .O(N__24696),
            .I(\quad_counter1.a_delay_counter_5 ));
    LocalMux I__2327 (
            .O(N__24693),
            .I(\quad_counter1.a_delay_counter_5 ));
    InMux I__2326 (
            .O(N__24688),
            .I(\quad_counter1.n19522 ));
    InMux I__2325 (
            .O(N__24685),
            .I(\quad_counter1.n19523 ));
    InMux I__2324 (
            .O(N__24682),
            .I(N__24678));
    InMux I__2323 (
            .O(N__24681),
            .I(N__24675));
    LocalMux I__2322 (
            .O(N__24678),
            .I(N__24672));
    LocalMux I__2321 (
            .O(N__24675),
            .I(\quad_counter1.a_delay_counter_7 ));
    Odrv4 I__2320 (
            .O(N__24672),
            .I(\quad_counter1.a_delay_counter_7 ));
    InMux I__2319 (
            .O(N__24667),
            .I(\quad_counter1.n19524 ));
    InMux I__2318 (
            .O(N__24664),
            .I(N__24660));
    InMux I__2317 (
            .O(N__24663),
            .I(N__24657));
    LocalMux I__2316 (
            .O(N__24660),
            .I(N__24654));
    LocalMux I__2315 (
            .O(N__24657),
            .I(\quad_counter1.a_delay_counter_8 ));
    Odrv4 I__2314 (
            .O(N__24654),
            .I(\quad_counter1.a_delay_counter_8 ));
    InMux I__2313 (
            .O(N__24649),
            .I(bfn_10_10_0_));
    InMux I__2312 (
            .O(N__24646),
            .I(\quad_counter1.n19526 ));
    InMux I__2311 (
            .O(N__24643),
            .I(N__24640));
    LocalMux I__2310 (
            .O(N__24640),
            .I(N__24636));
    InMux I__2309 (
            .O(N__24639),
            .I(N__24633));
    Span4Mux_h I__2308 (
            .O(N__24636),
            .I(N__24630));
    LocalMux I__2307 (
            .O(N__24633),
            .I(r_Tx_Data_6));
    Odrv4 I__2306 (
            .O(N__24630),
            .I(r_Tx_Data_6));
    InMux I__2305 (
            .O(N__24625),
            .I(N__24622));
    LocalMux I__2304 (
            .O(N__24622),
            .I(N__24618));
    InMux I__2303 (
            .O(N__24621),
            .I(N__24615));
    Span4Mux_h I__2302 (
            .O(N__24618),
            .I(N__24612));
    LocalMux I__2301 (
            .O(N__24615),
            .I(r_Tx_Data_2));
    Odrv4 I__2300 (
            .O(N__24612),
            .I(r_Tx_Data_2));
    CascadeMux I__2299 (
            .O(N__24607),
            .I(b_delay_counter_15__N_4141_cascade_));
    InMux I__2298 (
            .O(N__24604),
            .I(bfn_10_9_0_));
    InMux I__2297 (
            .O(N__24601),
            .I(N__24597));
    InMux I__2296 (
            .O(N__24600),
            .I(N__24594));
    LocalMux I__2295 (
            .O(N__24597),
            .I(data_out_frame_0_2));
    LocalMux I__2294 (
            .O(N__24594),
            .I(data_out_frame_0_2));
    InMux I__2293 (
            .O(N__24589),
            .I(N__24586));
    LocalMux I__2292 (
            .O(N__24586),
            .I(\c0.n6_adj_4521 ));
    CascadeMux I__2291 (
            .O(N__24583),
            .I(\c0.n23859_cascade_ ));
    CascadeMux I__2290 (
            .O(N__24580),
            .I(n23861_cascade_));
    CascadeMux I__2289 (
            .O(N__24577),
            .I(N__24574));
    InMux I__2288 (
            .O(N__24574),
            .I(N__24571));
    LocalMux I__2287 (
            .O(N__24571),
            .I(N__24568));
    Odrv4 I__2286 (
            .O(N__24568),
            .I(n10_adj_4534));
    CascadeMux I__2285 (
            .O(N__24565),
            .I(N__24562));
    InMux I__2284 (
            .O(N__24562),
            .I(N__24559));
    LocalMux I__2283 (
            .O(N__24559),
            .I(\c0.n5_adj_4522 ));
    CascadeMux I__2282 (
            .O(N__24556),
            .I(N__24553));
    InMux I__2281 (
            .O(N__24553),
            .I(N__24547));
    InMux I__2280 (
            .O(N__24552),
            .I(N__24547));
    LocalMux I__2279 (
            .O(N__24547),
            .I(data_out_frame_6_2));
    InMux I__2278 (
            .O(N__24544),
            .I(N__24541));
    LocalMux I__2277 (
            .O(N__24541),
            .I(\c0.n24007 ));
    InMux I__2276 (
            .O(N__24538),
            .I(N__24535));
    LocalMux I__2275 (
            .O(N__24535),
            .I(\c0.n6 ));
    CascadeMux I__2274 (
            .O(N__24532),
            .I(N__24529));
    InMux I__2273 (
            .O(N__24529),
            .I(N__24526));
    LocalMux I__2272 (
            .O(N__24526),
            .I(\c0.n11_adj_4348 ));
    InMux I__2271 (
            .O(N__24523),
            .I(N__24520));
    LocalMux I__2270 (
            .O(N__24520),
            .I(N__24517));
    Odrv4 I__2269 (
            .O(N__24517),
            .I(n24102));
    InMux I__2268 (
            .O(N__24514),
            .I(N__24511));
    LocalMux I__2267 (
            .O(N__24511),
            .I(\c0.n24047 ));
    InMux I__2266 (
            .O(N__24508),
            .I(N__24505));
    LocalMux I__2265 (
            .O(N__24505),
            .I(\c0.n5_adj_4358 ));
    CascadeMux I__2264 (
            .O(N__24502),
            .I(N__24499));
    InMux I__2263 (
            .O(N__24499),
            .I(N__24493));
    InMux I__2262 (
            .O(N__24498),
            .I(N__24493));
    LocalMux I__2261 (
            .O(N__24493),
            .I(data_out_frame_6_7));
    InMux I__2260 (
            .O(N__24490),
            .I(N__24486));
    InMux I__2259 (
            .O(N__24489),
            .I(N__24483));
    LocalMux I__2258 (
            .O(N__24486),
            .I(data_out_frame_0_3));
    LocalMux I__2257 (
            .O(N__24483),
            .I(data_out_frame_0_3));
    InMux I__2256 (
            .O(N__24478),
            .I(N__24475));
    LocalMux I__2255 (
            .O(N__24475),
            .I(N__24472));
    Odrv4 I__2254 (
            .O(N__24472),
            .I(\c0.n24011 ));
    InMux I__2253 (
            .O(N__24469),
            .I(N__24466));
    LocalMux I__2252 (
            .O(N__24466),
            .I(\c0.n11_adj_4355 ));
    InMux I__2251 (
            .O(N__24463),
            .I(N__24460));
    LocalMux I__2250 (
            .O(N__24460),
            .I(n23846));
    CascadeMux I__2249 (
            .O(N__24457),
            .I(n24114_cascade_));
    InMux I__2248 (
            .O(N__24454),
            .I(N__24451));
    LocalMux I__2247 (
            .O(N__24451),
            .I(N__24448));
    Span4Mux_h I__2246 (
            .O(N__24448),
            .I(N__24445));
    Odrv4 I__2245 (
            .O(N__24445),
            .I(n10));
    InMux I__2244 (
            .O(N__24442),
            .I(N__24439));
    LocalMux I__2243 (
            .O(N__24439),
            .I(N__24436));
    Span4Mux_h I__2242 (
            .O(N__24436),
            .I(N__24433));
    Odrv4 I__2241 (
            .O(N__24433),
            .I(\c0.n23895 ));
    CascadeMux I__2240 (
            .O(N__24430),
            .I(\c0.n24051_cascade_ ));
    InMux I__2239 (
            .O(N__24427),
            .I(N__24424));
    LocalMux I__2238 (
            .O(N__24424),
            .I(\c0.n23844 ));
    InMux I__2237 (
            .O(N__24421),
            .I(N__24418));
    LocalMux I__2236 (
            .O(N__24418),
            .I(N__24415));
    Odrv4 I__2235 (
            .O(N__24415),
            .I(\c0.n23847 ));
    InMux I__2234 (
            .O(N__24412),
            .I(N__24409));
    LocalMux I__2233 (
            .O(N__24409),
            .I(n24112));
    CascadeMux I__2232 (
            .O(N__24406),
            .I(n23849_cascade_));
    InMux I__2231 (
            .O(N__24403),
            .I(N__24399));
    InMux I__2230 (
            .O(N__24402),
            .I(N__24396));
    LocalMux I__2229 (
            .O(N__24399),
            .I(N__24393));
    LocalMux I__2228 (
            .O(N__24396),
            .I(data_out_frame_10_3));
    Odrv4 I__2227 (
            .O(N__24393),
            .I(data_out_frame_10_3));
    CascadeMux I__2226 (
            .O(N__24388),
            .I(\c0.n24159_cascade_ ));
    InMux I__2225 (
            .O(N__24385),
            .I(N__24382));
    LocalMux I__2224 (
            .O(N__24382),
            .I(N__24379));
    Odrv4 I__2223 (
            .O(N__24379),
            .I(\c0.n24162 ));
    InMux I__2222 (
            .O(N__24376),
            .I(N__24373));
    LocalMux I__2221 (
            .O(N__24373),
            .I(N__24370));
    Odrv12 I__2220 (
            .O(N__24370),
            .I(n26));
    CascadeMux I__2219 (
            .O(N__24367),
            .I(n24118_cascade_));
    CascadeMux I__2218 (
            .O(N__24364),
            .I(\c0.n23950_cascade_ ));
    CascadeMux I__2217 (
            .O(N__24361),
            .I(\c0.n24147_cascade_ ));
    InMux I__2216 (
            .O(N__24358),
            .I(N__24355));
    LocalMux I__2215 (
            .O(N__24355),
            .I(N__24352));
    Odrv4 I__2214 (
            .O(N__24352),
            .I(\c0.n23882 ));
    InMux I__2213 (
            .O(N__24349),
            .I(N__24346));
    LocalMux I__2212 (
            .O(N__24346),
            .I(n24150));
    CascadeMux I__2211 (
            .O(N__24343),
            .I(n24097_cascade_));
    InMux I__2210 (
            .O(N__24340),
            .I(N__24337));
    LocalMux I__2209 (
            .O(N__24337),
            .I(n24117));
    InMux I__2208 (
            .O(N__24334),
            .I(\quad_counter1.n19517 ));
    InMux I__2207 (
            .O(N__24331),
            .I(N__24327));
    InMux I__2206 (
            .O(N__24330),
            .I(N__24324));
    LocalMux I__2205 (
            .O(N__24327),
            .I(N__24321));
    LocalMux I__2204 (
            .O(N__24324),
            .I(\quad_counter1.b_delay_counter_15 ));
    Odrv4 I__2203 (
            .O(N__24321),
            .I(\quad_counter1.b_delay_counter_15 ));
    CascadeMux I__2202 (
            .O(N__24316),
            .I(N__24312));
    CEMux I__2201 (
            .O(N__24315),
            .I(N__24308));
    InMux I__2200 (
            .O(N__24312),
            .I(N__24305));
    CEMux I__2199 (
            .O(N__24311),
            .I(N__24302));
    LocalMux I__2198 (
            .O(N__24308),
            .I(N__24299));
    LocalMux I__2197 (
            .O(N__24305),
            .I(N__24294));
    LocalMux I__2196 (
            .O(N__24302),
            .I(N__24294));
    Span4Mux_h I__2195 (
            .O(N__24299),
            .I(N__24291));
    Span4Mux_h I__2194 (
            .O(N__24294),
            .I(N__24288));
    Odrv4 I__2193 (
            .O(N__24291),
            .I(n14377));
    Odrv4 I__2192 (
            .O(N__24288),
            .I(n14377));
    SRMux I__2191 (
            .O(N__24283),
            .I(N__24279));
    SRMux I__2190 (
            .O(N__24282),
            .I(N__24275));
    LocalMux I__2189 (
            .O(N__24279),
            .I(N__24272));
    InMux I__2188 (
            .O(N__24278),
            .I(N__24268));
    LocalMux I__2187 (
            .O(N__24275),
            .I(N__24265));
    Span4Mux_v I__2186 (
            .O(N__24272),
            .I(N__24262));
    InMux I__2185 (
            .O(N__24271),
            .I(N__24259));
    LocalMux I__2184 (
            .O(N__24268),
            .I(b_delay_counter_15__N_4141_adj_4548));
    Odrv12 I__2183 (
            .O(N__24265),
            .I(b_delay_counter_15__N_4141_adj_4548));
    Odrv4 I__2182 (
            .O(N__24262),
            .I(b_delay_counter_15__N_4141_adj_4548));
    LocalMux I__2181 (
            .O(N__24259),
            .I(b_delay_counter_15__N_4141_adj_4548));
    InMux I__2180 (
            .O(N__24250),
            .I(N__24247));
    LocalMux I__2179 (
            .O(N__24247),
            .I(\quad_counter1.A_delayed ));
    InMux I__2178 (
            .O(N__24244),
            .I(N__24240));
    InMux I__2177 (
            .O(N__24243),
            .I(N__24237));
    LocalMux I__2176 (
            .O(N__24240),
            .I(N__24233));
    LocalMux I__2175 (
            .O(N__24237),
            .I(N__24230));
    InMux I__2174 (
            .O(N__24236),
            .I(N__24227));
    Span4Mux_h I__2173 (
            .O(N__24233),
            .I(N__24224));
    Odrv12 I__2172 (
            .O(N__24230),
            .I(B_filtered_adj_4539));
    LocalMux I__2171 (
            .O(N__24227),
            .I(B_filtered_adj_4539));
    Odrv4 I__2170 (
            .O(N__24224),
            .I(B_filtered_adj_4539));
    CascadeMux I__2169 (
            .O(N__24217),
            .I(count_enable_adj_4544_cascade_));
    InMux I__2168 (
            .O(N__24214),
            .I(N__24208));
    InMux I__2167 (
            .O(N__24213),
            .I(N__24208));
    LocalMux I__2166 (
            .O(N__24208),
            .I(data_out_frame_10_6));
    InMux I__2165 (
            .O(N__24205),
            .I(N__24202));
    LocalMux I__2164 (
            .O(N__24202),
            .I(N__24198));
    InMux I__2163 (
            .O(N__24201),
            .I(N__24195));
    Span4Mux_h I__2162 (
            .O(N__24198),
            .I(N__24192));
    LocalMux I__2161 (
            .O(N__24195),
            .I(\quad_counter1.b_delay_counter_7 ));
    Odrv4 I__2160 (
            .O(N__24192),
            .I(\quad_counter1.b_delay_counter_7 ));
    InMux I__2159 (
            .O(N__24187),
            .I(\quad_counter1.n19509 ));
    CascadeMux I__2158 (
            .O(N__24184),
            .I(N__24181));
    InMux I__2157 (
            .O(N__24181),
            .I(N__24177));
    InMux I__2156 (
            .O(N__24180),
            .I(N__24174));
    LocalMux I__2155 (
            .O(N__24177),
            .I(N__24171));
    LocalMux I__2154 (
            .O(N__24174),
            .I(\quad_counter1.b_delay_counter_8 ));
    Odrv4 I__2153 (
            .O(N__24171),
            .I(\quad_counter1.b_delay_counter_8 ));
    InMux I__2152 (
            .O(N__24166),
            .I(bfn_9_11_0_));
    InMux I__2151 (
            .O(N__24163),
            .I(N__24160));
    LocalMux I__2150 (
            .O(N__24160),
            .I(N__24156));
    InMux I__2149 (
            .O(N__24159),
            .I(N__24153));
    Span4Mux_v I__2148 (
            .O(N__24156),
            .I(N__24150));
    LocalMux I__2147 (
            .O(N__24153),
            .I(\quad_counter1.b_delay_counter_9 ));
    Odrv4 I__2146 (
            .O(N__24150),
            .I(\quad_counter1.b_delay_counter_9 ));
    InMux I__2145 (
            .O(N__24145),
            .I(\quad_counter1.n19511 ));
    InMux I__2144 (
            .O(N__24142),
            .I(N__24138));
    InMux I__2143 (
            .O(N__24141),
            .I(N__24135));
    LocalMux I__2142 (
            .O(N__24138),
            .I(N__24132));
    LocalMux I__2141 (
            .O(N__24135),
            .I(\quad_counter1.b_delay_counter_10 ));
    Odrv4 I__2140 (
            .O(N__24132),
            .I(\quad_counter1.b_delay_counter_10 ));
    InMux I__2139 (
            .O(N__24127),
            .I(\quad_counter1.n19512 ));
    InMux I__2138 (
            .O(N__24124),
            .I(N__24120));
    InMux I__2137 (
            .O(N__24123),
            .I(N__24117));
    LocalMux I__2136 (
            .O(N__24120),
            .I(N__24114));
    LocalMux I__2135 (
            .O(N__24117),
            .I(\quad_counter1.b_delay_counter_11 ));
    Odrv12 I__2134 (
            .O(N__24114),
            .I(\quad_counter1.b_delay_counter_11 ));
    InMux I__2133 (
            .O(N__24109),
            .I(\quad_counter1.n19513 ));
    CascadeMux I__2132 (
            .O(N__24106),
            .I(N__24103));
    InMux I__2131 (
            .O(N__24103),
            .I(N__24099));
    InMux I__2130 (
            .O(N__24102),
            .I(N__24096));
    LocalMux I__2129 (
            .O(N__24099),
            .I(N__24093));
    LocalMux I__2128 (
            .O(N__24096),
            .I(\quad_counter1.b_delay_counter_12 ));
    Odrv4 I__2127 (
            .O(N__24093),
            .I(\quad_counter1.b_delay_counter_12 ));
    InMux I__2126 (
            .O(N__24088),
            .I(\quad_counter1.n19514 ));
    InMux I__2125 (
            .O(N__24085),
            .I(N__24082));
    LocalMux I__2124 (
            .O(N__24082),
            .I(N__24078));
    InMux I__2123 (
            .O(N__24081),
            .I(N__24075));
    Span4Mux_h I__2122 (
            .O(N__24078),
            .I(N__24072));
    LocalMux I__2121 (
            .O(N__24075),
            .I(\quad_counter1.b_delay_counter_13 ));
    Odrv4 I__2120 (
            .O(N__24072),
            .I(\quad_counter1.b_delay_counter_13 ));
    InMux I__2119 (
            .O(N__24067),
            .I(\quad_counter1.n19515 ));
    InMux I__2118 (
            .O(N__24064),
            .I(N__24060));
    InMux I__2117 (
            .O(N__24063),
            .I(N__24057));
    LocalMux I__2116 (
            .O(N__24060),
            .I(N__24054));
    LocalMux I__2115 (
            .O(N__24057),
            .I(\quad_counter1.b_delay_counter_14 ));
    Odrv4 I__2114 (
            .O(N__24054),
            .I(\quad_counter1.b_delay_counter_14 ));
    InMux I__2113 (
            .O(N__24049),
            .I(\quad_counter1.n19516 ));
    InMux I__2112 (
            .O(N__24046),
            .I(N__24043));
    LocalMux I__2111 (
            .O(N__24043),
            .I(N__24038));
    InMux I__2110 (
            .O(N__24042),
            .I(N__24033));
    InMux I__2109 (
            .O(N__24041),
            .I(N__24033));
    Odrv4 I__2108 (
            .O(N__24038),
            .I(b_delay_counter_0_adj_4541));
    LocalMux I__2107 (
            .O(N__24033),
            .I(b_delay_counter_0_adj_4541));
    InMux I__2106 (
            .O(N__24028),
            .I(N__24025));
    LocalMux I__2105 (
            .O(N__24025),
            .I(N__24022));
    Odrv12 I__2104 (
            .O(N__24022),
            .I(n187_adj_4546));
    InMux I__2103 (
            .O(N__24019),
            .I(bfn_9_10_0_));
    InMux I__2102 (
            .O(N__24016),
            .I(N__24013));
    LocalMux I__2101 (
            .O(N__24013),
            .I(N__24009));
    InMux I__2100 (
            .O(N__24012),
            .I(N__24006));
    Span4Mux_h I__2099 (
            .O(N__24009),
            .I(N__24003));
    LocalMux I__2098 (
            .O(N__24006),
            .I(\quad_counter1.b_delay_counter_1 ));
    Odrv4 I__2097 (
            .O(N__24003),
            .I(\quad_counter1.b_delay_counter_1 ));
    InMux I__2096 (
            .O(N__23998),
            .I(\quad_counter1.n19503 ));
    CascadeMux I__2095 (
            .O(N__23995),
            .I(N__23992));
    InMux I__2094 (
            .O(N__23992),
            .I(N__23989));
    LocalMux I__2093 (
            .O(N__23989),
            .I(N__23985));
    InMux I__2092 (
            .O(N__23988),
            .I(N__23982));
    Span4Mux_h I__2091 (
            .O(N__23985),
            .I(N__23979));
    LocalMux I__2090 (
            .O(N__23982),
            .I(\quad_counter1.b_delay_counter_2 ));
    Odrv4 I__2089 (
            .O(N__23979),
            .I(\quad_counter1.b_delay_counter_2 ));
    InMux I__2088 (
            .O(N__23974),
            .I(\quad_counter1.n19504 ));
    InMux I__2087 (
            .O(N__23971),
            .I(N__23967));
    InMux I__2086 (
            .O(N__23970),
            .I(N__23964));
    LocalMux I__2085 (
            .O(N__23967),
            .I(N__23961));
    LocalMux I__2084 (
            .O(N__23964),
            .I(\quad_counter1.b_delay_counter_3 ));
    Odrv4 I__2083 (
            .O(N__23961),
            .I(\quad_counter1.b_delay_counter_3 ));
    InMux I__2082 (
            .O(N__23956),
            .I(\quad_counter1.n19505 ));
    CascadeMux I__2081 (
            .O(N__23953),
            .I(N__23950));
    InMux I__2080 (
            .O(N__23950),
            .I(N__23946));
    InMux I__2079 (
            .O(N__23949),
            .I(N__23943));
    LocalMux I__2078 (
            .O(N__23946),
            .I(N__23940));
    LocalMux I__2077 (
            .O(N__23943),
            .I(\quad_counter1.b_delay_counter_4 ));
    Odrv4 I__2076 (
            .O(N__23940),
            .I(\quad_counter1.b_delay_counter_4 ));
    InMux I__2075 (
            .O(N__23935),
            .I(\quad_counter1.n19506 ));
    InMux I__2074 (
            .O(N__23932),
            .I(N__23929));
    LocalMux I__2073 (
            .O(N__23929),
            .I(N__23925));
    InMux I__2072 (
            .O(N__23928),
            .I(N__23922));
    Span4Mux_v I__2071 (
            .O(N__23925),
            .I(N__23919));
    LocalMux I__2070 (
            .O(N__23922),
            .I(\quad_counter1.b_delay_counter_5 ));
    Odrv4 I__2069 (
            .O(N__23919),
            .I(\quad_counter1.b_delay_counter_5 ));
    InMux I__2068 (
            .O(N__23914),
            .I(\quad_counter1.n19507 ));
    InMux I__2067 (
            .O(N__23911),
            .I(N__23908));
    LocalMux I__2066 (
            .O(N__23908),
            .I(N__23904));
    InMux I__2065 (
            .O(N__23907),
            .I(N__23901));
    Span4Mux_h I__2064 (
            .O(N__23904),
            .I(N__23898));
    LocalMux I__2063 (
            .O(N__23901),
            .I(\quad_counter1.b_delay_counter_6 ));
    Odrv4 I__2062 (
            .O(N__23898),
            .I(\quad_counter1.b_delay_counter_6 ));
    InMux I__2061 (
            .O(N__23893),
            .I(\quad_counter1.n19508 ));
    SRMux I__2060 (
            .O(N__23890),
            .I(N__23887));
    LocalMux I__2059 (
            .O(N__23887),
            .I(N__23884));
    Sp12to4 I__2058 (
            .O(N__23884),
            .I(N__23881));
    Odrv12 I__2057 (
            .O(N__23881),
            .I(\c0.n21322 ));
    InMux I__2056 (
            .O(N__23878),
            .I(N__23875));
    LocalMux I__2055 (
            .O(N__23875),
            .I(N__23872));
    Span4Mux_v I__2054 (
            .O(N__23872),
            .I(N__23868));
    InMux I__2053 (
            .O(N__23871),
            .I(N__23865));
    Sp12to4 I__2052 (
            .O(N__23868),
            .I(N__23860));
    LocalMux I__2051 (
            .O(N__23865),
            .I(N__23860));
    Span12Mux_h I__2050 (
            .O(N__23860),
            .I(N__23857));
    Odrv12 I__2049 (
            .O(N__23857),
            .I(rx_i));
    InMux I__2048 (
            .O(N__23854),
            .I(N__23851));
    LocalMux I__2047 (
            .O(N__23851),
            .I(\quad_counter1.n27 ));
    CascadeMux I__2046 (
            .O(N__23848),
            .I(\quad_counter1.n28_cascade_ ));
    InMux I__2045 (
            .O(N__23845),
            .I(N__23842));
    LocalMux I__2044 (
            .O(N__23842),
            .I(\quad_counter1.n25 ));
    CascadeMux I__2043 (
            .O(N__23839),
            .I(n9818_cascade_));
    InMux I__2042 (
            .O(N__23836),
            .I(\c0.n19616 ));
    InMux I__2041 (
            .O(N__23833),
            .I(\c0.n19617 ));
    InMux I__2040 (
            .O(N__23830),
            .I(\c0.n19618 ));
    CascadeMux I__2039 (
            .O(N__23827),
            .I(n23768_cascade_));
    CascadeMux I__2038 (
            .O(N__23824),
            .I(n23897_cascade_));
    CascadeMux I__2037 (
            .O(N__23821),
            .I(n10_adj_4532_cascade_));
    CascadeMux I__2036 (
            .O(N__23818),
            .I(\quad_counter1.n26_adj_4207_cascade_ ));
    InMux I__2035 (
            .O(N__23815),
            .I(N__23812));
    LocalMux I__2034 (
            .O(N__23812),
            .I(\quad_counter1.n25_adj_4209 ));
    InMux I__2033 (
            .O(N__23809),
            .I(N__23806));
    LocalMux I__2032 (
            .O(N__23806),
            .I(N__23803));
    Odrv4 I__2031 (
            .O(N__23803),
            .I(n12907));
    CascadeMux I__2030 (
            .O(N__23800),
            .I(N__23795));
    InMux I__2029 (
            .O(N__23799),
            .I(N__23790));
    InMux I__2028 (
            .O(N__23798),
            .I(N__23790));
    InMux I__2027 (
            .O(N__23795),
            .I(N__23787));
    LocalMux I__2026 (
            .O(N__23790),
            .I(N__23784));
    LocalMux I__2025 (
            .O(N__23787),
            .I(quadB_delayed_adj_4543));
    Odrv4 I__2024 (
            .O(N__23784),
            .I(quadB_delayed_adj_4543));
    InMux I__2023 (
            .O(N__23779),
            .I(N__23773));
    InMux I__2022 (
            .O(N__23778),
            .I(N__23773));
    LocalMux I__2021 (
            .O(N__23773),
            .I(N__23768));
    InMux I__2020 (
            .O(N__23772),
            .I(N__23763));
    InMux I__2019 (
            .O(N__23771),
            .I(N__23763));
    Span4Mux_v I__2018 (
            .O(N__23768),
            .I(N__23760));
    LocalMux I__2017 (
            .O(N__23763),
            .I(N__23757));
    Sp12to4 I__2016 (
            .O(N__23760),
            .I(N__23752));
    Sp12to4 I__2015 (
            .O(N__23757),
            .I(N__23752));
    Span12Mux_v I__2014 (
            .O(N__23752),
            .I(N__23749));
    Odrv12 I__2013 (
            .O(N__23749),
            .I(PIN_13_c));
    CascadeMux I__2012 (
            .O(N__23746),
            .I(n12907_cascade_));
    InMux I__2011 (
            .O(N__23743),
            .I(N__23740));
    LocalMux I__2010 (
            .O(N__23740),
            .I(\quad_counter1.n27_adj_4208 ));
    InMux I__2009 (
            .O(N__23737),
            .I(N__23734));
    LocalMux I__2008 (
            .O(N__23734),
            .I(\quad_counter1.n28_adj_4206 ));
    InMux I__2007 (
            .O(N__23731),
            .I(\c0.n19612 ));
    InMux I__2006 (
            .O(N__23728),
            .I(\c0.n19613 ));
    InMux I__2005 (
            .O(N__23725),
            .I(\c0.n19614 ));
    InMux I__2004 (
            .O(N__23722),
            .I(\c0.n19615 ));
    IoInMux I__2003 (
            .O(N__23719),
            .I(N__23716));
    LocalMux I__2002 (
            .O(N__23716),
            .I(N__23713));
    IoSpan4Mux I__2001 (
            .O(N__23713),
            .I(N__23710));
    Span4Mux_s3_v I__2000 (
            .O(N__23710),
            .I(N__23707));
    Sp12to4 I__1999 (
            .O(N__23707),
            .I(N__23704));
    Span12Mux_v I__1998 (
            .O(N__23704),
            .I(N__23701));
    Span12Mux_v I__1997 (
            .O(N__23701),
            .I(N__23698));
    Odrv12 I__1996 (
            .O(N__23698),
            .I(CLK_c));
    IoInMux I__1995 (
            .O(N__23695),
            .I(N__23692));
    LocalMux I__1994 (
            .O(N__23692),
            .I(tx_enable));
    IoInMux I__1993 (
            .O(N__23689),
            .I(N__23686));
    LocalMux I__1992 (
            .O(N__23686),
            .I(GB_BUFFER_PIN_9_c_THRU_CO));
    IoInMux I__1991 (
            .O(N__23683),
            .I(N__23680));
    LocalMux I__1990 (
            .O(N__23680),
            .I(N__23677));
    Span12Mux_s2_v I__1989 (
            .O(N__23677),
            .I(N__23674));
    Span12Mux_v I__1988 (
            .O(N__23674),
            .I(N__23671));
    Odrv12 I__1987 (
            .O(N__23671),
            .I(LED_c));
    defparam IN_MUX_bfv_10_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_13_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(\quad_counter1.n19555 ),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(\quad_counter1.n19563 ),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(\quad_counter1.n19571 ),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(\quad_counter1.n19579 ),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(\quad_counter0.n19587 ),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\quad_counter0.n19595 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\quad_counter0.n19603 ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\quad_counter0.n19611 ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(\quad_counter1.n19510 ),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(\quad_counter1.n19525 ),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_10_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_23_0_ (
            .carryinitin(\quad_counter0.n19480 ),
            .carryinitout(bfn_10_23_0_));
    defparam IN_MUX_bfv_10_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_24_0_));
    defparam IN_MUX_bfv_10_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_25_0_ (
            .carryinitin(\quad_counter0.n19495 ),
            .carryinitout(bfn_10_25_0_));
    defparam IN_MUX_bfv_13_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_21_0_));
    defparam IN_MUX_bfv_13_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_22_0_ (
            .carryinitin(\c0.tx.n19547 ),
            .carryinitout(bfn_13_22_0_));
    defparam IN_MUX_bfv_20_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_24_0_));
    defparam IN_MUX_bfv_7_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_17_0_));
    defparam IN_MUX_bfv_19_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_1_0_));
    defparam IN_MUX_bfv_19_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_2_0_ (
            .carryinitin(\c0.n19442_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_2_0_));
    defparam IN_MUX_bfv_19_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_3_0_ (
            .carryinitin(\c0.n19443_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_3_0_));
    defparam IN_MUX_bfv_19_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_4_0_ (
            .carryinitin(\c0.n19444_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_4_0_));
    defparam IN_MUX_bfv_19_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_5_0_ (
            .carryinitin(\c0.n19445_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_5_0_));
    defparam IN_MUX_bfv_19_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_6_0_ (
            .carryinitin(\c0.n19446_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_6_0_));
    defparam IN_MUX_bfv_19_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_7_0_ (
            .carryinitin(\c0.n19447_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_7_0_));
    defparam IN_MUX_bfv_19_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_8_0_ (
            .carryinitin(\c0.n19448_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_8_0_));
    defparam IN_MUX_bfv_19_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_9_0_ (
            .carryinitin(\c0.n19449_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_9_0_));
    defparam IN_MUX_bfv_19_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_10_0_ (
            .carryinitin(\c0.n19450_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_10_0_));
    defparam IN_MUX_bfv_19_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_11_0_ (
            .carryinitin(\c0.n19451_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_11_0_));
    defparam IN_MUX_bfv_19_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_12_0_ (
            .carryinitin(\c0.n19452_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_12_0_));
    defparam IN_MUX_bfv_19_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_13_0_ (
            .carryinitin(\c0.n19453_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_13_0_));
    defparam IN_MUX_bfv_19_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_14_0_ (
            .carryinitin(\c0.n19454_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_14_0_));
    defparam IN_MUX_bfv_19_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_15_0_ (
            .carryinitin(\c0.n19455_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_15_0_));
    defparam IN_MUX_bfv_19_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_16_0_ (
            .carryinitin(\c0.n19456_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_16_0_));
    defparam IN_MUX_bfv_19_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_17_0_ (
            .carryinitin(\c0.n19457_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_17_0_));
    defparam IN_MUX_bfv_19_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_18_0_ (
            .carryinitin(\c0.n19458_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_18_0_));
    defparam IN_MUX_bfv_19_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_19_0_ (
            .carryinitin(\c0.n19459_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_19_0_));
    defparam IN_MUX_bfv_19_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_20_0_ (
            .carryinitin(\c0.n19460_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_20_0_));
    defparam IN_MUX_bfv_19_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_21_0_ (
            .carryinitin(\c0.n19461_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_21_0_));
    defparam IN_MUX_bfv_19_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_22_0_ (
            .carryinitin(\c0.n19462_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_22_0_));
    defparam IN_MUX_bfv_19_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_23_0_ (
            .carryinitin(\c0.n19463_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_23_0_));
    defparam IN_MUX_bfv_19_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_24_0_ (
            .carryinitin(\c0.n19464_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_24_0_));
    defparam IN_MUX_bfv_19_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_25_0_ (
            .carryinitin(\c0.n19465_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_25_0_));
    defparam IN_MUX_bfv_19_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_26_0_ (
            .carryinitin(\c0.n19466_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_26_0_));
    defparam IN_MUX_bfv_19_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_27_0_ (
            .carryinitin(\c0.n19467_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_27_0_));
    defparam IN_MUX_bfv_19_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_28_0_ (
            .carryinitin(\c0.n19468_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_28_0_));
    defparam IN_MUX_bfv_19_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_29_0_ (
            .carryinitin(\c0.n19469_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_29_0_));
    defparam IN_MUX_bfv_19_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_30_0_ (
            .carryinitin(\c0.n19470_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_30_0_));
    defparam IN_MUX_bfv_19_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_31_0_ (
            .carryinitin(\c0.n19471_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_31_0_));
    defparam IN_MUX_bfv_19_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_32_0_ (
            .carryinitin(\c0.n19472_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_32_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \c0.tx.i8_1_lut_LC_1_3_6 .C_ON=1'b0;
    defparam \c0.tx.i8_1_lut_LC_1_3_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i8_1_lut_LC_1_3_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx.i8_1_lut_LC_1_3_6  (
            .in0(N__26517),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(tx_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_PIN_9_c_THRU_LUT4_0_LC_1_19_1.C_ON=1'b0;
    defparam GB_BUFFER_PIN_9_c_THRU_LUT4_0_LC_1_19_1.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_PIN_9_c_THRU_LUT4_0_LC_1_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_PIN_9_c_THRU_LUT4_0_LC_1_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66880),
            .lcout(GB_BUFFER_PIN_9_c_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rx_i_I_0_1_lut_LC_5_9_1.C_ON=1'b0;
    defparam rx_i_I_0_1_lut_LC_5_9_1.SEQ_MODE=4'b0000;
    defparam rx_i_I_0_1_lut_LC_5_9_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 rx_i_I_0_1_lut_LC_5_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23871),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.quadB_delayed_62_LC_5_21_5 .C_ON=1'b0;
    defparam \quad_counter0.quadB_delayed_62_LC_5_21_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.quadB_delayed_62_LC_5_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.quadB_delayed_62_LC_5_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27574),
            .lcout(quadB_delayed),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66869),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i23_LC_6_21_7 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i23_LC_6_21_7 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i23_LC_6_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i23_LC_6_21_7  (
            .in0(_gnd_net_),
            .in1(N__37641),
            .in2(_gnd_net_),
            .in3(N__52868),
            .lcout(\c0.FRAME_MATCHER_state_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66867),
            .ce(),
            .sr(N__23890));
    defparam \c0.FRAME_MATCHER_state_i26_LC_6_22_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i26_LC_6_22_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i26_LC_6_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i26_LC_6_22_0  (
            .in0(_gnd_net_),
            .in1(N__37318),
            .in2(_gnd_net_),
            .in3(N__52891),
            .lcout(\c0.FRAME_MATCHER_state_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66870),
            .ce(),
            .sr(N__29245));
    defparam \quad_counter1.quadA_delayed_61_LC_7_7_0 .C_ON=1'b0;
    defparam \quad_counter1.quadA_delayed_61_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.quadA_delayed_61_LC_7_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter1.quadA_delayed_61_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25946),
            .lcout(quadA_delayed_adj_4542),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66695),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.B_65_LC_7_9_4 .C_ON=1'b0;
    defparam \quad_counter1.B_65_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.B_65_LC_7_9_4 .LUT_INIT=16'b1010101011101000;
    LogicCell40 \quad_counter1.B_65_LC_7_9_4  (
            .in0(N__24236),
            .in1(N__23771),
            .in2(N__23800),
            .in3(N__23809),
            .lcout(B_filtered_adj_4539),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66723),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.quadB_delayed_62_LC_7_9_5 .C_ON=1'b0;
    defparam \quad_counter1.quadB_delayed_62_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.quadB_delayed_62_LC_7_9_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \quad_counter1.quadB_delayed_62_LC_7_9_5  (
            .in0(N__23772),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(quadB_delayed_adj_4543),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66723),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i9_4_lut_adj_1169_LC_7_10_2 .C_ON=1'b0;
    defparam \quad_counter1.i9_4_lut_adj_1169_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i9_4_lut_adj_1169_LC_7_10_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \quad_counter1.i9_4_lut_adj_1169_LC_7_10_2  (
            .in0(N__24163),
            .in1(N__23971),
            .in2(N__23953),
            .in3(N__24041),
            .lcout(\quad_counter1.n25_adj_4209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.b_delay_counter__i0_LC_7_10_4 .C_ON=1'b0;
    defparam \quad_counter1.b_delay_counter__i0_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i0_LC_7_10_4 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \quad_counter1.b_delay_counter__i0_LC_7_10_4  (
            .in0(N__24028),
            .in1(N__24042),
            .in2(N__24316),
            .in3(N__24278),
            .lcout(b_delay_counter_0_adj_4541),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66737),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.quadB_I_0_79_2_lut_LC_7_11_0 .C_ON=1'b0;
    defparam \quad_counter1.quadB_I_0_79_2_lut_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.quadB_I_0_79_2_lut_LC_7_11_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \quad_counter1.quadB_I_0_79_2_lut_LC_7_11_0  (
            .in0(N__23798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23779),
            .lcout(b_delay_counter_15__N_4141_adj_4548),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i10_4_lut_adj_1167_LC_7_11_2 .C_ON=1'b0;
    defparam \quad_counter1.i10_4_lut_adj_1167_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i10_4_lut_adj_1167_LC_7_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i10_4_lut_adj_1167_LC_7_11_2  (
            .in0(N__24142),
            .in1(N__24124),
            .in2(N__24184),
            .in3(N__23911),
            .lcout(),
            .ltout(\quad_counter1.n26_adj_4207_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i15_4_lut_adj_1170_LC_7_11_3 .C_ON=1'b0;
    defparam \quad_counter1.i15_4_lut_adj_1170_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i15_4_lut_adj_1170_LC_7_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i15_4_lut_adj_1170_LC_7_11_3  (
            .in0(N__23737),
            .in1(N__23743),
            .in2(N__23818),
            .in3(N__23815),
            .lcout(n12907),
            .ltout(n12907_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_1918_LC_7_11_4.C_ON=1'b0;
    defparam i1_4_lut_adj_1918_LC_7_11_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_1918_LC_7_11_4.LUT_INIT=16'b1111111110010000;
    LogicCell40 i1_4_lut_adj_1918_LC_7_11_4 (
            .in0(N__23799),
            .in1(N__23778),
            .in2(N__23746),
            .in3(N__24271),
            .lcout(n14377),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i11_4_lut_adj_1168_LC_7_11_5 .C_ON=1'b0;
    defparam \quad_counter1.i11_4_lut_adj_1168_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i11_4_lut_adj_1168_LC_7_11_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i11_4_lut_adj_1168_LC_7_11_5  (
            .in0(N__24064),
            .in1(N__24205),
            .in2(N__24106),
            .in3(N__24331),
            .lcout(\quad_counter1.n27_adj_4208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i12_4_lut_adj_1166_LC_7_11_6 .C_ON=1'b0;
    defparam \quad_counter1.i12_4_lut_adj_1166_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i12_4_lut_adj_1166_LC_7_11_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \quad_counter1.i12_4_lut_adj_1166_LC_7_11_6  (
            .in0(N__24016),
            .in1(N__24085),
            .in2(N__23995),
            .in3(N__23932),
            .lcout(\quad_counter1.n28_adj_4206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1411__i0_LC_7_17_0 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1411__i0_LC_7_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1411__i0_LC_7_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1411__i0_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__39189),
            .in2(N__39720),
            .in3(_gnd_net_),
            .lcout(\c0.byte_transmit_counter_0 ),
            .ltout(),
            .carryin(bfn_7_17_0_),
            .carryout(\c0.n19612 ),
            .clk(N__66822),
            .ce(N__39220),
            .sr(N__39202));
    defparam \c0.byte_transmit_counter_1411__i1_LC_7_17_1 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1411__i1_LC_7_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1411__i1_LC_7_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1411__i1_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__36742),
            .in2(_gnd_net_),
            .in3(N__23731),
            .lcout(\c0.byte_transmit_counter_1 ),
            .ltout(),
            .carryin(\c0.n19612 ),
            .carryout(\c0.n19613 ),
            .clk(N__66822),
            .ce(N__39220),
            .sr(N__39202));
    defparam \c0.byte_transmit_counter_1411__i2_LC_7_17_2 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1411__i2_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1411__i2_LC_7_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1411__i2_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(N__33863),
            .in2(_gnd_net_),
            .in3(N__23728),
            .lcout(\c0.byte_transmit_counter_2 ),
            .ltout(),
            .carryin(\c0.n19613 ),
            .carryout(\c0.n19614 ),
            .clk(N__66822),
            .ce(N__39220),
            .sr(N__39202));
    defparam \c0.byte_transmit_counter_1411__i3_LC_7_17_3 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1411__i3_LC_7_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1411__i3_LC_7_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1411__i3_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(N__25626),
            .in2(_gnd_net_),
            .in3(N__23725),
            .lcout(byte_transmit_counter_3),
            .ltout(),
            .carryin(\c0.n19614 ),
            .carryout(\c0.n19615 ),
            .clk(N__66822),
            .ce(N__39220),
            .sr(N__39202));
    defparam \c0.byte_transmit_counter_1411__i4_LC_7_17_4 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1411__i4_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1411__i4_LC_7_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1411__i4_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(N__26742),
            .in2(_gnd_net_),
            .in3(N__23722),
            .lcout(byte_transmit_counter_4),
            .ltout(),
            .carryin(\c0.n19615 ),
            .carryout(\c0.n19616 ),
            .clk(N__66822),
            .ce(N__39220),
            .sr(N__39202));
    defparam \c0.byte_transmit_counter_1411__i5_LC_7_17_5 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1411__i5_LC_7_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1411__i5_LC_7_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1411__i5_LC_7_17_5  (
            .in0(_gnd_net_),
            .in1(N__27308),
            .in2(_gnd_net_),
            .in3(N__23836),
            .lcout(byte_transmit_counter_5),
            .ltout(),
            .carryin(\c0.n19616 ),
            .carryout(\c0.n19617 ),
            .clk(N__66822),
            .ce(N__39220),
            .sr(N__39202));
    defparam \c0.byte_transmit_counter_1411__i6_LC_7_17_6 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1411__i6_LC_7_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1411__i6_LC_7_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1411__i6_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(N__26931),
            .in2(_gnd_net_),
            .in3(N__23833),
            .lcout(\c0.byte_transmit_counter_6 ),
            .ltout(),
            .carryin(\c0.n19617 ),
            .carryout(\c0.n19618 ),
            .clk(N__66822),
            .ce(N__39220),
            .sr(N__39202));
    defparam \c0.byte_transmit_counter_1411__i7_LC_7_17_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1411__i7_LC_7_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1411__i7_LC_7_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1411__i7_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(N__26910),
            .in2(_gnd_net_),
            .in3(N__23830),
            .lcout(\c0.byte_transmit_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66822),
            .ce(N__39220),
            .sr(N__39202));
    defparam \c0.i2_3_lut_adj_1673_LC_7_18_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1673_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1673_LC_7_18_4 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \c0.i2_3_lut_adj_1673_LC_7_18_4  (
            .in0(N__36741),
            .in1(N__33854),
            .in2(_gnd_net_),
            .in3(N__25589),
            .lcout(n23768),
            .ltout(n23768_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20202_4_lut_LC_7_18_5 .C_ON=1'b0;
    defparam \c0.i20202_4_lut_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20202_4_lut_LC_7_18_5 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \c0.i20202_4_lut_LC_7_18_5  (
            .in0(N__29443),
            .in1(N__24442),
            .in2(N__23827),
            .in3(N__26743),
            .lcout(),
            .ltout(n23897_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_1913_LC_7_18_6.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_1913_LC_7_18_6.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_1913_LC_7_18_6.LUT_INIT=16'b1110010011110000;
    LogicCell40 i24_3_lut_4_lut_adj_1913_LC_7_18_6 (
            .in0(N__26744),
            .in1(N__24523),
            .in2(N__23824),
            .in3(N__25590),
            .lcout(),
            .ltout(n10_adj_4532_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i5_LC_7_18_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i5_LC_7_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i5_LC_7_18_7 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \c0.tx.r_Tx_Data_i5_LC_7_18_7  (
            .in0(N__29154),
            .in1(N__25521),
            .in2(N__23821),
            .in3(N__27309),
            .lcout(r_Tx_Data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66834),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i2_LC_7_19_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i2_LC_7_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i2_LC_7_19_6 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.tx.r_Tx_Data_i2_LC_7_19_6  (
            .in0(N__24621),
            .in1(N__27322),
            .in2(N__24577),
            .in3(N__29144),
            .lcout(r_Tx_Data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66846),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i6_LC_7_19_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i6_LC_7_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i6_LC_7_19_7 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \c0.tx.r_Tx_Data_i6_LC_7_19_7  (
            .in0(N__29145),
            .in1(N__24639),
            .in2(N__27334),
            .in3(N__24454),
            .lcout(r_Tx_Data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66846),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1517_LC_7_21_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1517_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1517_LC_7_21_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_1517_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__37640),
            .in2(_gnd_net_),
            .in3(N__40657),
            .lcout(\c0.n21322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_R_49_LC_9_8_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_R_49_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_R_49_LC_9_8_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.rx.r_Rx_Data_R_49_LC_9_8_1  (
            .in0(N__23878),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.rx.r_Rx_Data_R ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66681),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i26_3_lut_LC_9_8_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i26_3_lut_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i26_3_lut_LC_9_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_4_i26_3_lut_LC_9_8_6  (
            .in0(N__39838),
            .in1(N__26098),
            .in2(_gnd_net_),
            .in3(N__29254),
            .lcout(n26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__1__5428_LC_9_8_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__1__5428_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__1__5428_LC_9_8_7 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.data_out_frame_12__1__5428_LC_9_8_7  (
            .in0(N__34710),
            .in1(N__49179),
            .in2(N__32311),
            .in3(N__49040),
            .lcout(data_out_frame_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66681),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i9_4_lut_LC_9_9_0 .C_ON=1'b0;
    defparam \quad_counter1.i9_4_lut_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i9_4_lut_LC_9_9_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \quad_counter1.i9_4_lut_LC_9_9_0  (
            .in0(N__24699),
            .in1(N__24840),
            .in2(N__24718),
            .in3(N__24889),
            .lcout(\quad_counter1.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i11_4_lut_LC_9_9_1 .C_ON=1'b0;
    defparam \quad_counter1.i11_4_lut_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i11_4_lut_LC_9_9_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i11_4_lut_LC_9_9_1  (
            .in0(N__24819),
            .in1(N__24682),
            .in2(N__24859),
            .in3(N__24801),
            .lcout(\quad_counter1.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i12_4_lut_LC_9_9_2 .C_ON=1'b0;
    defparam \quad_counter1.i12_4_lut_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i12_4_lut_LC_9_9_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \quad_counter1.i12_4_lut_LC_9_9_2  (
            .in0(N__24732),
            .in1(N__24664),
            .in2(N__24751),
            .in3(N__24768),
            .lcout(),
            .ltout(\quad_counter1.n28_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i15_4_lut_LC_9_9_3 .C_ON=1'b0;
    defparam \quad_counter1.i15_4_lut_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i15_4_lut_LC_9_9_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i15_4_lut_LC_9_9_3  (
            .in0(N__26032),
            .in1(N__23854),
            .in2(N__23848),
            .in3(N__23845),
            .lcout(n9818),
            .ltout(n9818_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.A_63_LC_9_9_4 .C_ON=1'b0;
    defparam \quad_counter1.A_63_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.A_63_LC_9_9_4 .LUT_INIT=16'b1111111000001000;
    LogicCell40 \quad_counter1.A_63_LC_9_9_4  (
            .in0(N__25959),
            .in1(N__25993),
            .in2(N__23839),
            .in3(N__24938),
            .lcout(A_filtered_adj_4538),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66696),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1073_1_lut_2_lut_LC_9_9_6 .C_ON=1'b0;
    defparam \quad_counter1.i1073_1_lut_2_lut_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1073_1_lut_2_lut_LC_9_9_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \quad_counter1.i1073_1_lut_2_lut_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__24911),
            .in2(_gnd_net_),
            .in3(N__24937),
            .lcout(\quad_counter1.n2140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.B_delayed_68_LC_9_9_7 .C_ON=1'b0;
    defparam \quad_counter1.B_delayed_68_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.B_delayed_68_LC_9_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter1.B_delayed_68_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24243),
            .lcout(\quad_counter1.B_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66696),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_86_2_lut_LC_9_10_0 .C_ON=1'b1;
    defparam \quad_counter1.add_86_2_lut_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_86_2_lut_LC_9_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_86_2_lut_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__24046),
            .in2(_gnd_net_),
            .in3(N__24019),
            .lcout(n187_adj_4546),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\quad_counter1.n19503 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.b_delay_counter__i1_LC_9_10_1 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i1_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i1_LC_9_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i1_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__24012),
            .in2(_gnd_net_),
            .in3(N__23998),
            .lcout(\quad_counter1.b_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter1.n19503 ),
            .carryout(\quad_counter1.n19504 ),
            .clk(N__66709),
            .ce(N__24311),
            .sr(N__24283));
    defparam \quad_counter1.b_delay_counter__i2_LC_9_10_2 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i2_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i2_LC_9_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i2_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__23988),
            .in2(_gnd_net_),
            .in3(N__23974),
            .lcout(\quad_counter1.b_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter1.n19504 ),
            .carryout(\quad_counter1.n19505 ),
            .clk(N__66709),
            .ce(N__24311),
            .sr(N__24283));
    defparam \quad_counter1.b_delay_counter__i3_LC_9_10_3 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i3_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i3_LC_9_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i3_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__23970),
            .in2(_gnd_net_),
            .in3(N__23956),
            .lcout(\quad_counter1.b_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter1.n19505 ),
            .carryout(\quad_counter1.n19506 ),
            .clk(N__66709),
            .ce(N__24311),
            .sr(N__24283));
    defparam \quad_counter1.b_delay_counter__i4_LC_9_10_4 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i4_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i4_LC_9_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i4_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__23949),
            .in2(_gnd_net_),
            .in3(N__23935),
            .lcout(\quad_counter1.b_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter1.n19506 ),
            .carryout(\quad_counter1.n19507 ),
            .clk(N__66709),
            .ce(N__24311),
            .sr(N__24283));
    defparam \quad_counter1.b_delay_counter__i5_LC_9_10_5 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i5_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i5_LC_9_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i5_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__23928),
            .in2(_gnd_net_),
            .in3(N__23914),
            .lcout(\quad_counter1.b_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter1.n19507 ),
            .carryout(\quad_counter1.n19508 ),
            .clk(N__66709),
            .ce(N__24311),
            .sr(N__24283));
    defparam \quad_counter1.b_delay_counter__i6_LC_9_10_6 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i6_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i6_LC_9_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i6_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__23907),
            .in2(_gnd_net_),
            .in3(N__23893),
            .lcout(\quad_counter1.b_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter1.n19508 ),
            .carryout(\quad_counter1.n19509 ),
            .clk(N__66709),
            .ce(N__24311),
            .sr(N__24283));
    defparam \quad_counter1.b_delay_counter__i7_LC_9_10_7 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i7_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i7_LC_9_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i7_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__24201),
            .in2(_gnd_net_),
            .in3(N__24187),
            .lcout(\quad_counter1.b_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter1.n19509 ),
            .carryout(\quad_counter1.n19510 ),
            .clk(N__66709),
            .ce(N__24311),
            .sr(N__24283));
    defparam \quad_counter1.b_delay_counter__i8_LC_9_11_0 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i8_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i8_LC_9_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i8_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__24180),
            .in2(_gnd_net_),
            .in3(N__24166),
            .lcout(\quad_counter1.b_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\quad_counter1.n19511 ),
            .clk(N__66724),
            .ce(N__24315),
            .sr(N__24282));
    defparam \quad_counter1.b_delay_counter__i9_LC_9_11_1 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i9_LC_9_11_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i9_LC_9_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i9_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__24159),
            .in2(_gnd_net_),
            .in3(N__24145),
            .lcout(\quad_counter1.b_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter1.n19511 ),
            .carryout(\quad_counter1.n19512 ),
            .clk(N__66724),
            .ce(N__24315),
            .sr(N__24282));
    defparam \quad_counter1.b_delay_counter__i10_LC_9_11_2 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i10_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i10_LC_9_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i10_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__24141),
            .in2(_gnd_net_),
            .in3(N__24127),
            .lcout(\quad_counter1.b_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter1.n19512 ),
            .carryout(\quad_counter1.n19513 ),
            .clk(N__66724),
            .ce(N__24315),
            .sr(N__24282));
    defparam \quad_counter1.b_delay_counter__i11_LC_9_11_3 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i11_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i11_LC_9_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i11_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__24123),
            .in2(_gnd_net_),
            .in3(N__24109),
            .lcout(\quad_counter1.b_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter1.n19513 ),
            .carryout(\quad_counter1.n19514 ),
            .clk(N__66724),
            .ce(N__24315),
            .sr(N__24282));
    defparam \quad_counter1.b_delay_counter__i12_LC_9_11_4 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i12_LC_9_11_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i12_LC_9_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i12_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__24102),
            .in2(_gnd_net_),
            .in3(N__24088),
            .lcout(\quad_counter1.b_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter1.n19514 ),
            .carryout(\quad_counter1.n19515 ),
            .clk(N__66724),
            .ce(N__24315),
            .sr(N__24282));
    defparam \quad_counter1.b_delay_counter__i13_LC_9_11_5 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i13_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i13_LC_9_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i13_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__24081),
            .in2(_gnd_net_),
            .in3(N__24067),
            .lcout(\quad_counter1.b_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter1.n19515 ),
            .carryout(\quad_counter1.n19516 ),
            .clk(N__66724),
            .ce(N__24315),
            .sr(N__24282));
    defparam \quad_counter1.b_delay_counter__i14_LC_9_11_6 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i14_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i14_LC_9_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i14_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__24063),
            .in2(_gnd_net_),
            .in3(N__24049),
            .lcout(\quad_counter1.b_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter1.n19516 ),
            .carryout(\quad_counter1.n19517 ),
            .clk(N__66724),
            .ce(N__24315),
            .sr(N__24282));
    defparam \quad_counter1.b_delay_counter__i15_LC_9_11_7 .C_ON=1'b0;
    defparam \quad_counter1.b_delay_counter__i15_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i15_LC_9_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i15_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__24330),
            .in2(_gnd_net_),
            .in3(N__24334),
            .lcout(\quad_counter1.b_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66724),
            .ce(N__24315),
            .sr(N__24282));
    defparam \quad_counter1.A_delayed_67_LC_9_12_0 .C_ON=1'b0;
    defparam \quad_counter1.A_delayed_67_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.A_delayed_67_LC_9_12_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \quad_counter1.A_delayed_67_LC_9_12_0  (
            .in0(N__24953),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\quad_counter1.A_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20187_4_lut_LC_9_12_1 .C_ON=1'b0;
    defparam \c0.i20187_4_lut_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i20187_4_lut_LC_9_12_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.i20187_4_lut_LC_9_12_1  (
            .in0(N__26446),
            .in1(N__36902),
            .in2(N__34654),
            .in3(N__33976),
            .lcout(\c0.n23882 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__0__5421_LC_9_12_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__0__5421_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__0__5421_LC_9_12_2 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.data_out_frame_13__0__5421_LC_9_12_2  (
            .in0(N__26212),
            .in1(N__49565),
            .in2(N__25027),
            .in3(N__49020),
            .lcout(data_out_frame_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1406_LC_9_12_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1406_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1406_LC_9_12_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1406_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__25021),
            .in2(_gnd_net_),
            .in3(N__26320),
            .lcout(\c0.n6_adj_4308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i3_4_lut_LC_9_12_4 .C_ON=1'b0;
    defparam \quad_counter1.i3_4_lut_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i3_4_lut_LC_9_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \quad_counter1.i3_4_lut_LC_9_12_4  (
            .in0(N__24919),
            .in1(N__24250),
            .in2(N__24955),
            .in3(N__24244),
            .lcout(count_enable_adj_4544),
            .ltout(count_enable_adj_4544_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i0_LC_9_12_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i0_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i0_LC_9_12_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \quad_counter1.count_i0_i0_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__24994),
            .in2(N__24217),
            .in3(N__25025),
            .lcout(encoder1_position_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66738),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i6_LC_9_12_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i6_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i6_LC_9_12_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i6_LC_9_12_7  (
            .in0(N__25060),
            .in1(N__38356),
            .in2(_gnd_net_),
            .in3(N__34957),
            .lcout(encoder1_position_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__6__5439_LC_9_13_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__6__5439_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__6__5439_LC_9_13_3 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_10__6__5439_LC_9_13_3  (
            .in0(N__49273),
            .in1(N__49022),
            .in2(N__35530),
            .in3(N__24214),
            .lcout(data_out_frame_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66751),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20461_LC_9_13_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20461_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20461_LC_9_13_4 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_20461_LC_9_13_4  (
            .in0(N__24213),
            .in1(N__36834),
            .in2(N__24790),
            .in3(N__39781),
            .lcout(\c0.n24153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__5__5464_LC_9_13_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__5__5464_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__5__5464_LC_9_13_5 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_7__5__5464_LC_9_13_5  (
            .in0(N__49274),
            .in1(N__49023),
            .in2(N__36004),
            .in3(N__26571),
            .lcout(data_out_frame_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66751),
            .ce(),
            .sr(_gnd_net_));
    defparam i20420_4_lut_LC_9_13_6.C_ON=1'b0;
    defparam i20420_4_lut_LC_9_13_6.SEQ_MODE=4'b0000;
    defparam i20420_4_lut_LC_9_13_6.LUT_INIT=16'b0101110000001100;
    LogicCell40 i20420_4_lut_LC_9_13_6 (
            .in0(N__26875),
            .in1(N__24340),
            .in2(N__26797),
            .in3(N__24376),
            .lcout(),
            .ltout(n24118_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i4_LC_9_13_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i4_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i4_LC_9_13_7 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \c0.tx.r_Tx_Data_i4_LC_9_13_7  (
            .in0(N__29155),
            .in1(N__25503),
            .in2(N__24367),
            .in3(N__27338),
            .lcout(r_Tx_Data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66751),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20414_4_lut_LC_9_14_0 .C_ON=1'b0;
    defparam \c0.i20414_4_lut_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i20414_4_lut_LC_9_14_0 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \c0.i20414_4_lut_LC_9_14_0  (
            .in0(N__26266),
            .in1(N__33969),
            .in2(N__36910),
            .in3(N__24385),
            .lcout(n24112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20399_2_lut_LC_9_14_1 .C_ON=1'b0;
    defparam \c0.i20399_2_lut_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i20399_2_lut_LC_9_14_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.i20399_2_lut_LC_9_14_1  (
            .in0(N__39758),
            .in1(N__30115),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n23950_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_9_14_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_9_14_2 .LUT_INIT=16'b1011100011001100;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_LC_9_14_2  (
            .in0(N__26248),
            .in1(N__36906),
            .in2(N__24364),
            .in3(N__33970),
            .lcout(),
            .ltout(\c0.n24147_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n24147_bdd_4_lut_4_lut_LC_9_14_3 .C_ON=1'b0;
    defparam \c0.n24147_bdd_4_lut_4_lut_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.n24147_bdd_4_lut_4_lut_LC_9_14_3 .LUT_INIT=16'b1111000010100100;
    LogicCell40 \c0.n24147_bdd_4_lut_4_lut_LC_9_14_3  (
            .in0(N__39759),
            .in1(N__25429),
            .in2(N__24361),
            .in3(N__33938),
            .lcout(n24150),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20400_4_lut_LC_9_14_4 .C_ON=1'b0;
    defparam \c0.i20400_4_lut_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i20400_4_lut_LC_9_14_4 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.i20400_4_lut_LC_9_14_4  (
            .in0(N__24358),
            .in1(N__36907),
            .in2(N__30214),
            .in3(N__33971),
            .lcout(),
            .ltout(n24097_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20419_3_lut_LC_9_14_5.C_ON=1'b0;
    defparam i20419_3_lut_LC_9_14_5.SEQ_MODE=4'b0000;
    defparam i20419_3_lut_LC_9_14_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 i20419_3_lut_LC_9_14_5 (
            .in0(_gnd_net_),
            .in1(N__24349),
            .in2(N__24343),
            .in3(N__25638),
            .lcout(n24117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__3__5442_LC_9_14_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__3__5442_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__3__5442_LC_9_14_6 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_10__3__5442_LC_9_14_6  (
            .in0(N__49379),
            .in1(N__49013),
            .in2(N__30175),
            .in3(N__24402),
            .lcout(data_out_frame_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66766),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i15_LC_9_15_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i15_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i15_LC_9_15_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i15_LC_9_15_1  (
            .in0(N__38411),
            .in1(N__25120),
            .in2(_gnd_net_),
            .in3(N__26311),
            .lcout(encoder1_position_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66778),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20154_4_lut_LC_9_15_2 .C_ON=1'b0;
    defparam \c0.i20154_4_lut_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i20154_4_lut_LC_9_15_2 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \c0.i20154_4_lut_LC_9_15_2  (
            .in0(N__34753),
            .in1(N__24421),
            .in2(N__26874),
            .in3(N__26789),
            .lcout(),
            .ltout(n23849_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_1915_LC_9_15_3.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_1915_LC_9_15_3.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_1915_LC_9_15_3.LUT_INIT=16'b1110010011110000;
    LogicCell40 i24_3_lut_4_lut_adj_1915_LC_9_15_3 (
            .in0(N__26790),
            .in1(N__24412),
            .in2(N__24406),
            .in3(N__25634),
            .lcout(n10_adj_4536),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_9_15_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_9_15_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_9_15_4  (
            .in0(N__29887),
            .in1(N__28543),
            .in2(_gnd_net_),
            .in3(N__39773),
            .lcout(\c0.n11_adj_4355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i28_LC_9_15_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i28_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i28_LC_9_15_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter1.count_i0_i28_LC_9_15_6  (
            .in0(N__36495),
            .in1(N__25336),
            .in2(_gnd_net_),
            .in3(N__38412),
            .lcout(encoder1_position_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66778),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20151_4_lut_LC_9_16_0 .C_ON=1'b0;
    defparam \c0.i20151_4_lut_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i20151_4_lut_LC_9_16_0 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \c0.i20151_4_lut_LC_9_16_0  (
            .in0(N__26865),
            .in1(N__24427),
            .in2(N__26796),
            .in3(N__29311),
            .lcout(n23846),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20476_LC_9_16_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20476_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20476_LC_9_16_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_20476_LC_9_16_2  (
            .in0(N__24403),
            .in1(N__36862),
            .in2(N__28525),
            .in3(N__39772),
            .lcout(\c0.n24171 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20466_LC_9_16_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20466_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20466_LC_9_16_3 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_20466_LC_9_16_3  (
            .in0(N__39771),
            .in1(N__28708),
            .in2(N__36900),
            .in3(N__28740),
            .lcout(),
            .ltout(\c0.n24159_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n24159_bdd_4_lut_LC_9_16_4 .C_ON=1'b0;
    defparam \c0.n24159_bdd_4_lut_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.n24159_bdd_4_lut_LC_9_16_4 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n24159_bdd_4_lut_LC_9_16_4  (
            .in0(N__26542),
            .in1(N__36863),
            .in2(N__24388),
            .in3(N__28723),
            .lcout(\c0.n24162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20416_4_lut_LC_9_16_5 .C_ON=1'b0;
    defparam \c0.i20416_4_lut_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20416_4_lut_LC_9_16_5 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \c0.i20416_4_lut_LC_9_16_5  (
            .in0(N__24469),
            .in1(N__33942),
            .in2(N__36901),
            .in3(N__28555),
            .lcout(),
            .ltout(n24114_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_1916_LC_9_16_6.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_1916_LC_9_16_6.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_1916_LC_9_16_6.LUT_INIT=16'b1101100011001100;
    LogicCell40 i24_3_lut_4_lut_adj_1916_LC_9_16_6 (
            .in0(N__26788),
            .in1(N__24463),
            .in2(N__24457),
            .in3(N__25635),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20200_4_lut_LC_9_17_0 .C_ON=1'b0;
    defparam \c0.i20200_4_lut_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i20200_4_lut_LC_9_17_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.i20200_4_lut_LC_9_17_0  (
            .in0(N__33889),
            .in1(N__36761),
            .in2(N__26557),
            .in3(N__24514),
            .lcout(\c0.n23895 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_9_17_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_9_17_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_9_17_1  (
            .in0(N__25410),
            .in1(N__38020),
            .in2(_gnd_net_),
            .in3(N__39701),
            .lcout(\c0.n11_adj_4348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i31_LC_9_17_3 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i31_LC_9_17_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i31_LC_9_17_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i31_LC_9_17_3  (
            .in0(N__25438),
            .in1(N__38458),
            .in2(_gnd_net_),
            .in3(N__28771),
            .lcout(encoder1_position_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66800),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i18_LC_9_17_4 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i18_LC_9_17_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i18_LC_9_17_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i18_LC_9_17_4  (
            .in0(N__25105),
            .in1(N__38457),
            .in2(_gnd_net_),
            .in3(N__29032),
            .lcout(encoder1_position_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66800),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20355_3_lut_LC_9_17_5 .C_ON=1'b0;
    defparam \c0.i20355_3_lut_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20355_3_lut_LC_9_17_5 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \c0.i20355_3_lut_LC_9_17_5  (
            .in0(N__26677),
            .in1(N__33886),
            .in2(_gnd_net_),
            .in3(N__39700),
            .lcout(),
            .ltout(\c0.n24051_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20149_4_lut_LC_9_17_6 .C_ON=1'b0;
    defparam \c0.i20149_4_lut_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i20149_4_lut_LC_9_17_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \c0.i20149_4_lut_LC_9_17_6  (
            .in0(N__33888),
            .in1(N__39514),
            .in2(N__24430),
            .in3(N__36760),
            .lcout(\c0.n23844 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20152_4_lut_LC_9_17_7 .C_ON=1'b0;
    defparam \c0.i20152_4_lut_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i20152_4_lut_LC_9_17_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \c0.i20152_4_lut_LC_9_17_7  (
            .in0(N__36759),
            .in1(N__33887),
            .in2(N__33790),
            .in3(N__24508),
            .lcout(\c0.n23847 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20404_4_lut_LC_9_18_0 .C_ON=1'b0;
    defparam \c0.i20404_4_lut_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i20404_4_lut_LC_9_18_0 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.i20404_4_lut_LC_9_18_0  (
            .in0(N__36848),
            .in1(N__27079),
            .in2(N__24532),
            .in3(N__33948),
            .lcout(n24102),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_0__3__5522_LC_9_18_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_0__3__5522_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_0__3__5522_LC_9_18_1 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \c0.data_out_frame_0__3__5522_LC_9_18_1  (
            .in0(N__24490),
            .in1(N__37193),
            .in2(_gnd_net_),
            .in3(N__40170),
            .lcout(data_out_frame_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66810),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20351_4_lut_LC_9_18_3 .C_ON=1'b0;
    defparam \c0.i20351_4_lut_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i20351_4_lut_LC_9_18_3 .LUT_INIT=16'b1011000100000000;
    LogicCell40 \c0.i20351_4_lut_LC_9_18_3  (
            .in0(N__33946),
            .in1(N__36847),
            .in2(N__27181),
            .in3(N__39775),
            .lcout(\c0.n24047 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_9_18_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_9_18_4 .LUT_INIT=16'b1010000001000100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_9_18_4  (
            .in0(N__39776),
            .in1(N__24478),
            .in2(N__26893),
            .in3(N__33947),
            .lcout(\c0.n6_adj_4521 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_9_18_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_9_18_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_9_18_5  (
            .in0(N__33436),
            .in1(N__24498),
            .in2(_gnd_net_),
            .in3(N__39774),
            .lcout(\c0.n5_adj_4358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__7__5470_LC_9_18_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__7__5470_LC_9_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__7__5470_LC_9_18_6 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_out_frame_6__7__5470_LC_9_18_6  (
            .in0(N__48844),
            .in1(N__49447),
            .in2(N__24502),
            .in3(N__41646),
            .lcout(data_out_frame_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66810),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__3__5418_LC_9_18_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__3__5418_LC_9_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__3__5418_LC_9_18_7 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_13__3__5418_LC_9_18_7  (
            .in0(N__49446),
            .in1(N__48845),
            .in2(N__28357),
            .in3(N__26658),
            .lcout(data_out_frame_13_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66810),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20385_2_lut_LC_9_19_0 .C_ON=1'b0;
    defparam \c0.i20385_2_lut_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i20385_2_lut_LC_9_19_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i20385_2_lut_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__24489),
            .in2(_gnd_net_),
            .in3(N__36870),
            .lcout(\c0.n24007 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20389_2_lut_LC_9_19_1 .C_ON=1'b0;
    defparam \c0.i20389_2_lut_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i20389_2_lut_LC_9_19_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.i20389_2_lut_LC_9_19_1  (
            .in0(N__36871),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24600),
            .lcout(\c0.n24011 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20161_4_lut_LC_9_19_2 .C_ON=1'b0;
    defparam \c0.i20161_4_lut_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i20161_4_lut_LC_9_19_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \c0.i20161_4_lut_LC_9_19_2  (
            .in0(N__24538),
            .in1(N__36872),
            .in2(N__27196),
            .in3(N__33964),
            .lcout(\c0.n23856 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_0__2__5523_LC_9_19_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_0__2__5523_LC_9_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_0__2__5523_LC_9_19_3 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \c0.data_out_frame_0__2__5523_LC_9_19_3  (
            .in0(N__24601),
            .in1(N__37204),
            .in2(_gnd_net_),
            .in3(N__40169),
            .lcout(data_out_frame_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66823),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20164_4_lut_LC_9_19_4 .C_ON=1'b0;
    defparam \c0.i20164_4_lut_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i20164_4_lut_LC_9_19_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \c0.i20164_4_lut_LC_9_19_4  (
            .in0(N__24589),
            .in1(N__36873),
            .in2(N__24565),
            .in3(N__33965),
            .lcout(),
            .ltout(\c0.n23859_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20166_4_lut_LC_9_19_5 .C_ON=1'b0;
    defparam \c0.i20166_4_lut_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20166_4_lut_LC_9_19_5 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.i20166_4_lut_LC_9_19_5  (
            .in0(N__26866),
            .in1(N__25858),
            .in2(N__24583),
            .in3(N__26791),
            .lcout(),
            .ltout(n23861_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_1911_LC_9_19_6.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_1911_LC_9_19_6.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_1911_LC_9_19_6.LUT_INIT=16'b1110010011110000;
    LogicCell40 i24_3_lut_4_lut_adj_1911_LC_9_19_6 (
            .in0(N__26792),
            .in1(N__25468),
            .in2(N__24580),
            .in3(N__25636),
            .lcout(n10_adj_4534),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_9_20_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_9_20_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_9_20_0  (
            .in0(N__26371),
            .in1(N__24552),
            .in2(_gnd_net_),
            .in3(N__39779),
            .lcout(\c0.n5_adj_4522 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__2__5475_LC_9_20_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__2__5475_LC_9_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__2__5475_LC_9_20_1 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_6__2__5475_LC_9_20_1  (
            .in0(N__49548),
            .in1(N__49021),
            .in2(N__24556),
            .in3(N__40063),
            .lcout(data_out_frame_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66835),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20362_4_lut_LC_9_20_3 .C_ON=1'b0;
    defparam \c0.i20362_4_lut_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i20362_4_lut_LC_9_20_3 .LUT_INIT=16'b1000000010001010;
    LogicCell40 \c0.i20362_4_lut_LC_9_20_3  (
            .in0(N__39780),
            .in1(N__28984),
            .in2(N__33975),
            .in3(N__36882),
            .lcout(\c0.n24059 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_9_20_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_9_20_6 .LUT_INIT=16'b1111001100100010;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_9_20_6  (
            .in0(N__24544),
            .in1(N__33959),
            .in2(N__27229),
            .in3(N__39778),
            .lcout(\c0.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Bit_Index_2__bdd_4_lut_LC_9_20_7.C_ON=1'b0;
    defparam r_Bit_Index_2__bdd_4_lut_LC_9_20_7.SEQ_MODE=4'b0000;
    defparam r_Bit_Index_2__bdd_4_lut_LC_9_20_7.LUT_INIT=16'b1010111111000000;
    LogicCell40 r_Bit_Index_2__bdd_4_lut_LC_9_20_7 (
            .in0(N__24643),
            .in1(N__24625),
            .in2(N__26989),
            .in3(N__27036),
            .lcout(n24195),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i0_LC_9_22_0 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i0_LC_9_22_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i0_LC_9_22_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \quad_counter0.b_delay_counter__i0_LC_9_22_0  (
            .in0(N__25769),
            .in1(N__25796),
            .in2(N__27607),
            .in3(N__25693),
            .lcout(b_delay_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66856),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.quadA_delayed_61_LC_9_22_4 .C_ON=1'b0;
    defparam \quad_counter0.quadA_delayed_61_LC_9_22_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.quadA_delayed_61_LC_9_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.quadA_delayed_61_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27824),
            .lcout(quadA_delayed),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66856),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.quadB_I_0_79_2_lut_LC_9_22_6 .C_ON=1'b0;
    defparam \quad_counter0.quadB_I_0_79_2_lut_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.quadB_I_0_79_2_lut_LC_9_22_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \quad_counter0.quadB_I_0_79_2_lut_LC_9_22_6  (
            .in0(N__27579),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27530),
            .lcout(b_delay_counter_15__N_4141),
            .ltout(b_delay_counter_15__N_4141_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_1917_LC_9_22_7.C_ON=1'b0;
    defparam i1_4_lut_adj_1917_LC_9_22_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_1917_LC_9_22_7.LUT_INIT=16'b1111100111110000;
    LogicCell40 i1_4_lut_adj_1917_LC_9_22_7 (
            .in0(N__27531),
            .in1(N__27578),
            .in2(N__24607),
            .in3(N__27376),
            .lcout(n14198),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i4_LC_9_23_6 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i4_LC_9_23_6 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i4_LC_9_23_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i4_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(N__37789),
            .in2(_gnd_net_),
            .in3(N__52890),
            .lcout(\c0.FRAME_MATCHER_state_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66864),
            .ce(),
            .sr(N__34210));
    defparam \quad_counter0.quadA_I_0_73_2_lut_LC_9_24_0 .C_ON=1'b0;
    defparam \quad_counter0.quadA_I_0_73_2_lut_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.quadA_I_0_73_2_lut_LC_9_24_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \quad_counter0.quadA_I_0_73_2_lut_LC_9_24_0  (
            .in0(N__27825),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27789),
            .lcout(a_delay_counter_15__N_4124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1708_LC_10_8_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1708_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1708_LC_10_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1708_LC_10_8_2  (
            .in0(N__28338),
            .in1(N__29710),
            .in2(_gnd_net_),
            .in3(N__53368),
            .lcout(\c0.n13360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1803_LC_10_8_6 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1803_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1803_LC_10_8_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1803_LC_10_8_6  (
            .in0(N__29425),
            .in1(N__32592),
            .in2(N__32566),
            .in3(N__31636),
            .lcout(\c0.n24_adj_4502 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_85_2_lut_LC_10_9_0 .C_ON=1'b1;
    defparam \quad_counter1.add_85_2_lut_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_85_2_lut_LC_10_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_85_2_lut_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__24887),
            .in2(_gnd_net_),
            .in3(N__24604),
            .lcout(n39_adj_4545),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\quad_counter1.n19518 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.a_delay_counter__i1_LC_10_9_1 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i1_LC_10_9_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i1_LC_10_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i1_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__24769),
            .in2(_gnd_net_),
            .in3(N__24754),
            .lcout(\quad_counter1.a_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter1.n19518 ),
            .carryout(\quad_counter1.n19519 ),
            .clk(N__66672),
            .ce(N__25906),
            .sr(N__26020));
    defparam \quad_counter1.a_delay_counter__i2_LC_10_9_2 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i2_LC_10_9_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i2_LC_10_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i2_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__24750),
            .in2(_gnd_net_),
            .in3(N__24736),
            .lcout(\quad_counter1.a_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter1.n19519 ),
            .carryout(\quad_counter1.n19520 ),
            .clk(N__66672),
            .ce(N__25906),
            .sr(N__26020));
    defparam \quad_counter1.a_delay_counter__i3_LC_10_9_3 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i3_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i3_LC_10_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i3_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__24733),
            .in2(_gnd_net_),
            .in3(N__24721),
            .lcout(\quad_counter1.a_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter1.n19520 ),
            .carryout(\quad_counter1.n19521 ),
            .clk(N__66672),
            .ce(N__25906),
            .sr(N__26020));
    defparam \quad_counter1.a_delay_counter__i4_LC_10_9_4 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i4_LC_10_9_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i4_LC_10_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i4_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__24717),
            .in2(_gnd_net_),
            .in3(N__24703),
            .lcout(\quad_counter1.a_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter1.n19521 ),
            .carryout(\quad_counter1.n19522 ),
            .clk(N__66672),
            .ce(N__25906),
            .sr(N__26020));
    defparam \quad_counter1.a_delay_counter__i5_LC_10_9_5 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i5_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i5_LC_10_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i5_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__24700),
            .in2(_gnd_net_),
            .in3(N__24688),
            .lcout(\quad_counter1.a_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter1.n19522 ),
            .carryout(\quad_counter1.n19523 ),
            .clk(N__66672),
            .ce(N__25906),
            .sr(N__26020));
    defparam \quad_counter1.a_delay_counter__i6_LC_10_9_6 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i6_LC_10_9_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i6_LC_10_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i6_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__26044),
            .in2(_gnd_net_),
            .in3(N__24685),
            .lcout(\quad_counter1.a_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter1.n19523 ),
            .carryout(\quad_counter1.n19524 ),
            .clk(N__66672),
            .ce(N__25906),
            .sr(N__26020));
    defparam \quad_counter1.a_delay_counter__i7_LC_10_9_7 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i7_LC_10_9_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i7_LC_10_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i7_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__24681),
            .in2(_gnd_net_),
            .in3(N__24667),
            .lcout(\quad_counter1.a_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter1.n19524 ),
            .carryout(\quad_counter1.n19525 ),
            .clk(N__66672),
            .ce(N__25906),
            .sr(N__26020));
    defparam \quad_counter1.a_delay_counter__i8_LC_10_10_0 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i8_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i8_LC_10_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i8_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(N__24663),
            .in2(_gnd_net_),
            .in3(N__24649),
            .lcout(\quad_counter1.a_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\quad_counter1.n19526 ),
            .clk(N__66683),
            .ce(N__25905),
            .sr(N__26016));
    defparam \quad_counter1.a_delay_counter__i9_LC_10_10_1 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i9_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i9_LC_10_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i9_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__26058),
            .in2(_gnd_net_),
            .in3(N__24646),
            .lcout(\quad_counter1.a_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter1.n19526 ),
            .carryout(\quad_counter1.n19527 ),
            .clk(N__66683),
            .ce(N__25905),
            .sr(N__26016));
    defparam \quad_counter1.a_delay_counter__i10_LC_10_10_2 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i10_LC_10_10_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i10_LC_10_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i10_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__24858),
            .in2(_gnd_net_),
            .in3(N__24844),
            .lcout(\quad_counter1.a_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter1.n19527 ),
            .carryout(\quad_counter1.n19528 ),
            .clk(N__66683),
            .ce(N__25905),
            .sr(N__26016));
    defparam \quad_counter1.a_delay_counter__i11_LC_10_10_3 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i11_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i11_LC_10_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i11_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__24841),
            .in2(_gnd_net_),
            .in3(N__24829),
            .lcout(\quad_counter1.a_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter1.n19528 ),
            .carryout(\quad_counter1.n19529 ),
            .clk(N__66683),
            .ce(N__25905),
            .sr(N__26016));
    defparam \quad_counter1.a_delay_counter__i12_LC_10_10_4 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i12_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i12_LC_10_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i12_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__26085),
            .in2(_gnd_net_),
            .in3(N__24826),
            .lcout(\quad_counter1.a_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter1.n19529 ),
            .carryout(\quad_counter1.n19530 ),
            .clk(N__66683),
            .ce(N__25905),
            .sr(N__26016));
    defparam \quad_counter1.a_delay_counter__i13_LC_10_10_5 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i13_LC_10_10_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i13_LC_10_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i13_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__26071),
            .in2(_gnd_net_),
            .in3(N__24823),
            .lcout(\quad_counter1.a_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter1.n19530 ),
            .carryout(\quad_counter1.n19531 ),
            .clk(N__66683),
            .ce(N__25905),
            .sr(N__26016));
    defparam \quad_counter1.a_delay_counter__i14_LC_10_10_6 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i14_LC_10_10_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i14_LC_10_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i14_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__24820),
            .in2(_gnd_net_),
            .in3(N__24808),
            .lcout(\quad_counter1.a_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter1.n19531 ),
            .carryout(\quad_counter1.n19532 ),
            .clk(N__66683),
            .ce(N__25905),
            .sr(N__26016));
    defparam \quad_counter1.a_delay_counter__i15_LC_10_10_7 .C_ON=1'b0;
    defparam \quad_counter1.a_delay_counter__i15_LC_10_10_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i15_LC_10_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i15_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(N__24802),
            .in2(_gnd_net_),
            .in3(N__24805),
            .lcout(\quad_counter1.a_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66683),
            .ce(N__25905),
            .sr(N__26016));
    defparam \c0.i3_4_lut_adj_1403_LC_10_11_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1403_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1403_LC_10_11_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1403_LC_10_11_0  (
            .in0(N__35390),
            .in1(N__33085),
            .in2(N__28219),
            .in3(N__28426),
            .lcout(\c0.n10434 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__6__5431_LC_10_11_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__6__5431_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__6__5431_LC_10_11_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_out_frame_11__6__5431_LC_10_11_1  (
            .in0(N__49017),
            .in1(N__49358),
            .in2(N__24789),
            .in3(N__28481),
            .lcout(data_out_frame_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66698),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i3_LC_10_11_3 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i3_LC_10_11_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i3_LC_10_11_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \quad_counter1.count_i0_i3_LC_10_11_3  (
            .in0(N__24970),
            .in1(_gnd_net_),
            .in2(N__38410),
            .in3(N__28325),
            .lcout(encoder1_position_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66698),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__4__5433_LC_10_11_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__4__5433_LC_10_11_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__4__5433_LC_10_11_4 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_11__4__5433_LC_10_11_4  (
            .in0(N__49357),
            .in1(N__49018),
            .in2(N__38941),
            .in3(N__26460),
            .lcout(data_out_frame_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66698),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.A_filtered_I_0_2_lut_LC_10_11_5 .C_ON=1'b0;
    defparam \quad_counter1.A_filtered_I_0_2_lut_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.A_filtered_I_0_2_lut_LC_10_11_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \quad_counter1.A_filtered_I_0_2_lut_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(N__24954),
            .in2(_gnd_net_),
            .in3(N__24918),
            .lcout(\quad_counter1.count_direction ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.a_delay_counter__i0_LC_10_11_6 .C_ON=1'b0;
    defparam \quad_counter1.a_delay_counter__i0_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i0_LC_10_11_6 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \quad_counter1.a_delay_counter__i0_LC_10_11_6  (
            .in0(N__26004),
            .in1(N__24898),
            .in2(N__24888),
            .in3(N__25904),
            .lcout(a_delay_counter_0_adj_4540),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66698),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i5_LC_10_11_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i5_LC_10_11_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i5_LC_10_11_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i5_LC_10_11_7  (
            .in0(N__38377),
            .in1(N__25072),
            .in2(_gnd_net_),
            .in3(N__32700),
            .lcout(encoder1_position_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66698),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1628_LC_10_12_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1628_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1628_LC_10_12_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1628_LC_10_12_0  (
            .in0(N__31190),
            .in1(N__34348),
            .in2(N__32448),
            .in3(N__32552),
            .lcout(\c0.n20257 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i14_LC_10_12_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i14_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i14_LC_10_12_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter1.count_i0_i14_LC_10_12_1  (
            .in0(N__29640),
            .in1(N__38357),
            .in2(_gnd_net_),
            .in3(N__25132),
            .lcout(encoder1_position_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66711),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i2_LC_10_12_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i2_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i2_LC_10_12_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \quad_counter1.count_i0_i2_LC_10_12_2  (
            .in0(N__38360),
            .in1(_gnd_net_),
            .in2(N__35042),
            .in3(N__24982),
            .lcout(encoder1_position_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66711),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i26_LC_10_12_3 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i26_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i26_LC_10_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter1.count_i0_i26_LC_10_12_3  (
            .in0(N__35644),
            .in1(N__25351),
            .in2(_gnd_net_),
            .in3(N__38359),
            .lcout(encoder1_position_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66711),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1405_LC_10_12_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1405_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1405_LC_10_12_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1405_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(N__36459),
            .in2(_gnd_net_),
            .in3(N__29639),
            .lcout(\c0.n22116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1807_LC_10_12_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1807_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1807_LC_10_12_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1807_LC_10_12_5  (
            .in0(_gnd_net_),
            .in1(N__32784),
            .in2(_gnd_net_),
            .in3(N__35031),
            .lcout(),
            .ltout(\c0.n22048_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1810_LC_10_12_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1810_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1810_LC_10_12_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1810_LC_10_12_6  (
            .in0(N__31813),
            .in1(N__32498),
            .in2(N__25030),
            .in3(N__28321),
            .lcout(\c0.n20819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i22_LC_10_12_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i22_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i22_LC_10_12_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter1.count_i0_i22_LC_10_12_7  (
            .in0(N__28470),
            .in1(N__25084),
            .in2(_gnd_net_),
            .in3(N__38358),
            .lcout(encoder1_position_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66711),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_1_LC_10_13_0 .C_ON=1'b1;
    defparam \quad_counter1.add_611_1_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_1_LC_10_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \quad_counter1.add_611_1_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(N__25179),
            .in2(N__25308),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_13_0_),
            .carryout(\quad_counter1.n19548 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_2_lut_LC_10_13_1 .C_ON=1'b1;
    defparam \quad_counter1.add_611_2_lut_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_2_lut_LC_10_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_2_lut_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__25026),
            .in2(N__25006),
            .in3(N__24988),
            .lcout(n2205),
            .ltout(),
            .carryin(\quad_counter1.n19548 ),
            .carryout(\quad_counter1.n19549 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_3_lut_LC_10_13_2 .C_ON=1'b1;
    defparam \quad_counter1.add_611_3_lut_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_3_lut_LC_10_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_3_lut_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__32785),
            .in2(N__25309),
            .in3(N__24985),
            .lcout(n2204),
            .ltout(),
            .carryin(\quad_counter1.n19549 ),
            .carryout(\quad_counter1.n19550 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_4_lut_LC_10_13_3 .C_ON=1'b1;
    defparam \quad_counter1.add_611_4_lut_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_4_lut_LC_10_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_4_lut_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(N__35035),
            .in2(N__25250),
            .in3(N__24973),
            .lcout(n2203),
            .ltout(),
            .carryin(\quad_counter1.n19550 ),
            .carryout(\quad_counter1.n19551 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_5_lut_LC_10_13_4 .C_ON=1'b1;
    defparam \quad_counter1.add_611_5_lut_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_5_lut_LC_10_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_5_lut_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(N__28334),
            .in2(N__25310),
            .in3(N__24961),
            .lcout(n2202),
            .ltout(),
            .carryin(\quad_counter1.n19551 ),
            .carryout(\quad_counter1.n19552 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_6_lut_LC_10_13_5 .C_ON=1'b1;
    defparam \quad_counter1.add_611_6_lut_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_6_lut_LC_10_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_6_lut_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(N__35139),
            .in2(N__25251),
            .in3(N__24958),
            .lcout(n2201),
            .ltout(),
            .carryin(\quad_counter1.n19552 ),
            .carryout(\quad_counter1.n19553 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_7_lut_LC_10_13_6 .C_ON=1'b1;
    defparam \quad_counter1.add_611_7_lut_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_7_lut_LC_10_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_7_lut_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(N__25186),
            .in2(N__32734),
            .in3(N__25063),
            .lcout(n2200),
            .ltout(),
            .carryin(\quad_counter1.n19553 ),
            .carryout(\quad_counter1.n19554 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_8_lut_LC_10_13_7 .C_ON=1'b1;
    defparam \quad_counter1.add_611_8_lut_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_8_lut_LC_10_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_8_lut_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(N__25261),
            .in2(N__34966),
            .in3(N__25054),
            .lcout(n2199),
            .ltout(),
            .carryin(\quad_counter1.n19554 ),
            .carryout(\quad_counter1.n19555 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_9_lut_LC_10_14_0 .C_ON=1'b1;
    defparam \quad_counter1.add_611_9_lut_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_9_lut_LC_10_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_9_lut_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__25262),
            .in2(N__34929),
            .in3(N__25051),
            .lcout(n2198),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\quad_counter1.n19556 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_10_lut_LC_10_14_1 .C_ON=1'b1;
    defparam \quad_counter1.add_611_10_lut_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_10_lut_LC_10_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_10_lut_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__35381),
            .in2(N__25311),
            .in3(N__25048),
            .lcout(n2197),
            .ltout(),
            .carryin(\quad_counter1.n19556 ),
            .carryout(\quad_counter1.n19557 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_11_lut_LC_10_14_2 .C_ON=1'b1;
    defparam \quad_counter1.add_611_11_lut_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_11_lut_LC_10_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_11_lut_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__25266),
            .in2(N__32310),
            .in3(N__25045),
            .lcout(n2196),
            .ltout(),
            .carryin(\quad_counter1.n19557 ),
            .carryout(\quad_counter1.n19558 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_12_lut_LC_10_14_3 .C_ON=1'b1;
    defparam \quad_counter1.add_611_12_lut_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_12_lut_LC_10_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_12_lut_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(N__35220),
            .in2(N__25312),
            .in3(N__25042),
            .lcout(n2195),
            .ltout(),
            .carryin(\quad_counter1.n19558 ),
            .carryout(\quad_counter1.n19559 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_13_lut_LC_10_14_4 .C_ON=1'b1;
    defparam \quad_counter1.add_611_13_lut_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_13_lut_LC_10_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_13_lut_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__25270),
            .in2(N__32980),
            .in3(N__25039),
            .lcout(n2194),
            .ltout(),
            .carryin(\quad_counter1.n19559 ),
            .carryout(\quad_counter1.n19560 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_14_lut_LC_10_14_5 .C_ON=1'b1;
    defparam \quad_counter1.add_611_14_lut_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_14_lut_LC_10_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_14_lut_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(N__34635),
            .in2(N__25313),
            .in3(N__25036),
            .lcout(n2193),
            .ltout(),
            .carryin(\quad_counter1.n19560 ),
            .carryout(\quad_counter1.n19561 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_15_lut_LC_10_14_6 .C_ON=1'b1;
    defparam \quad_counter1.add_611_15_lut_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_15_lut_LC_10_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_15_lut_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__25274),
            .in2(N__38070),
            .in3(N__25033),
            .lcout(n2192),
            .ltout(),
            .carryin(\quad_counter1.n19561 ),
            .carryout(\quad_counter1.n19562 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_16_lut_LC_10_14_7 .C_ON=1'b1;
    defparam \quad_counter1.add_611_16_lut_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_16_lut_LC_10_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_16_lut_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__29655),
            .in2(N__25314),
            .in3(N__25123),
            .lcout(n2191),
            .ltout(),
            .carryin(\quad_counter1.n19562 ),
            .carryout(\quad_counter1.n19563 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_17_lut_LC_10_15_0 .C_ON=1'b1;
    defparam \quad_counter1.add_611_17_lut_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_17_lut_LC_10_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_17_lut_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__26310),
            .in2(N__25315),
            .in3(N__25114),
            .lcout(n2190),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\quad_counter1.n19564 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_18_lut_LC_10_15_1 .C_ON=1'b1;
    defparam \quad_counter1.add_611_18_lut_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_18_lut_LC_10_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_18_lut_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__25281),
            .in2(N__26427),
            .in3(N__25111),
            .lcout(n2189),
            .ltout(),
            .carryin(\quad_counter1.n19564 ),
            .carryout(\quad_counter1.n19565 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_19_lut_LC_10_15_2 .C_ON=1'b1;
    defparam \quad_counter1.add_611_19_lut_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_19_lut_LC_10_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_19_lut_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__37246),
            .in2(N__25316),
            .in3(N__25108),
            .lcout(n2188),
            .ltout(),
            .carryin(\quad_counter1.n19565 ),
            .carryout(\quad_counter1.n19566 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_20_lut_LC_10_15_3 .C_ON=1'b1;
    defparam \quad_counter1.add_611_20_lut_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_20_lut_LC_10_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_20_lut_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__25285),
            .in2(N__29049),
            .in3(N__25096),
            .lcout(n2187),
            .ltout(),
            .carryin(\quad_counter1.n19566 ),
            .carryout(\quad_counter1.n19567 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_21_lut_LC_10_15_4 .C_ON=1'b1;
    defparam \quad_counter1.add_611_21_lut_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_21_lut_LC_10_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_21_lut_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__30034),
            .in2(N__25317),
            .in3(N__25093),
            .lcout(n2186),
            .ltout(),
            .carryin(\quad_counter1.n19567 ),
            .carryout(\quad_counter1.n19568 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_22_lut_LC_10_15_5 .C_ON=1'b1;
    defparam \quad_counter1.add_611_22_lut_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_22_lut_LC_10_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_22_lut_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__25289),
            .in2(N__38934),
            .in3(N__25090),
            .lcout(n2185),
            .ltout(),
            .carryin(\quad_counter1.n19568 ),
            .carryout(\quad_counter1.n19569 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_23_lut_LC_10_15_6 .C_ON=1'b1;
    defparam \quad_counter1.add_611_23_lut_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_23_lut_LC_10_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_23_lut_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__28606),
            .in2(N__25318),
            .in3(N__25087),
            .lcout(n2184),
            .ltout(),
            .carryin(\quad_counter1.n19569 ),
            .carryout(\quad_counter1.n19570 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_24_lut_LC_10_15_7 .C_ON=1'b1;
    defparam \quad_counter1.add_611_24_lut_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_24_lut_LC_10_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_24_lut_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__25293),
            .in2(N__28487),
            .in3(N__25075),
            .lcout(n2183),
            .ltout(),
            .carryin(\quad_counter1.n19570 ),
            .carryout(\quad_counter1.n19571 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_25_lut_LC_10_16_0 .C_ON=1'b1;
    defparam \quad_counter1.add_611_25_lut_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_25_lut_LC_10_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_25_lut_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__25294),
            .in2(N__32900),
            .in3(N__25360),
            .lcout(n2182),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\quad_counter1.n19572 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_26_lut_LC_10_16_1 .C_ON=1'b1;
    defparam \quad_counter1.add_611_26_lut_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_26_lut_LC_10_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_26_lut_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__29958),
            .in2(N__25319),
            .in3(N__25357),
            .lcout(n2181),
            .ltout(),
            .carryin(\quad_counter1.n19572 ),
            .carryout(\quad_counter1.n19573 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_27_lut_LC_10_16_2 .C_ON=1'b1;
    defparam \quad_counter1.add_611_27_lut_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_27_lut_LC_10_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_27_lut_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(N__25298),
            .in2(N__33022),
            .in3(N__25354),
            .lcout(n2180),
            .ltout(),
            .carryin(\quad_counter1.n19573 ),
            .carryout(\quad_counter1.n19574 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_28_lut_LC_10_16_3 .C_ON=1'b1;
    defparam \quad_counter1.add_611_28_lut_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_28_lut_LC_10_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_28_lut_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__35645),
            .in2(N__25320),
            .in3(N__25342),
            .lcout(n2179),
            .ltout(),
            .carryin(\quad_counter1.n19574 ),
            .carryout(\quad_counter1.n19575 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_29_lut_LC_10_16_4 .C_ON=1'b1;
    defparam \quad_counter1.add_611_29_lut_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_29_lut_LC_10_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_29_lut_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(N__25302),
            .in2(N__30171),
            .in3(N__25339),
            .lcout(n2178),
            .ltout(),
            .carryin(\quad_counter1.n19575 ),
            .carryout(\quad_counter1.n19576 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_30_lut_LC_10_16_5 .C_ON=1'b1;
    defparam \quad_counter1.add_611_30_lut_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_30_lut_LC_10_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_30_lut_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(N__25246),
            .in2(N__36503),
            .in3(N__25330),
            .lcout(n2177),
            .ltout(),
            .carryin(\quad_counter1.n19576 ),
            .carryout(\quad_counter1.n19577 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_31_lut_LC_10_16_6 .C_ON=1'b1;
    defparam \quad_counter1.add_611_31_lut_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_31_lut_LC_10_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_31_lut_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__28954),
            .in2(N__25307),
            .in3(N__25327),
            .lcout(n2176),
            .ltout(),
            .carryin(\quad_counter1.n19577 ),
            .carryout(\quad_counter1.n19578 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_32_lut_LC_10_16_7 .C_ON=1'b1;
    defparam \quad_counter1.add_611_32_lut_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_32_lut_LC_10_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_611_32_lut_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(N__35517),
            .in2(N__25321),
            .in3(N__25324),
            .lcout(n2175),
            .ltout(),
            .carryin(\quad_counter1.n19578 ),
            .carryout(\quad_counter1.n19579 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_611_33_lut_LC_10_17_0 .C_ON=1'b0;
    defparam \quad_counter1.add_611_33_lut_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_611_33_lut_LC_10_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \quad_counter1.add_611_33_lut_LC_10_17_0  (
            .in0(N__25306),
            .in1(N__28770),
            .in2(_gnd_net_),
            .in3(N__25441),
            .lcout(n2174),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20410_4_lut_LC_10_17_1 .C_ON=1'b0;
    defparam \c0.i20410_4_lut_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i20410_4_lut_LC_10_17_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.i20410_4_lut_LC_10_17_1  (
            .in0(N__25384),
            .in1(N__36765),
            .in2(N__27133),
            .in3(N__33937),
            .lcout(n24108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__3__5450_LC_10_17_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__3__5450_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__3__5450_LC_10_17_2 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_9__3__5450_LC_10_17_2  (
            .in0(N__49412),
            .in1(N__49007),
            .in2(N__41704),
            .in3(N__25399),
            .lcout(data_out_frame_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66780),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_0__4__5521_LC_10_17_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_0__4__5521_LC_10_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_0__4__5521_LC_10_17_3 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \c0.data_out_frame_0__4__5521_LC_10_17_3  (
            .in0(N__25425),
            .in1(N__37203),
            .in2(_gnd_net_),
            .in3(N__40171),
            .lcout(data_out_frame_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66780),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1600_LC_10_17_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1600_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1600_LC_10_17_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i2_2_lut_adj_1600_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(N__26745),
            .in2(_gnd_net_),
            .in3(N__25607),
            .lcout(\c0.n6_adj_4392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__5__5416_LC_10_17_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__5__5416_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__5__5416_LC_10_17_6 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_frame_13__5__5416_LC_10_17_6  (
            .in0(N__49411),
            .in1(N__25411),
            .in2(N__32740),
            .in3(N__49008),
            .lcout(data_out_frame_13_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66780),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n24171_bdd_4_lut_LC_10_17_7 .C_ON=1'b0;
    defparam \c0.n24171_bdd_4_lut_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.n24171_bdd_4_lut_LC_10_17_7 .LUT_INIT=16'b1100101111001000;
    LogicCell40 \c0.n24171_bdd_4_lut_LC_10_17_7  (
            .in0(N__25398),
            .in1(N__25390),
            .in2(N__36833),
            .in3(N__34675),
            .lcout(\c0.n24174 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__0__5437_LC_10_18_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__0__5437_LC_10_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__0__5437_LC_10_18_0 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.data_out_frame_11__0__5437_LC_10_18_0  (
            .in0(N__27156),
            .in1(N__49448),
            .in2(N__26428),
            .in3(N__48847),
            .lcout(data_out_frame_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66792),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20163_4_lut_LC_10_18_2 .C_ON=1'b0;
    defparam \c0.i20163_4_lut_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i20163_4_lut_LC_10_18_2 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \c0.i20163_4_lut_LC_10_18_2  (
            .in0(N__26780),
            .in1(N__26590),
            .in2(N__26864),
            .in3(N__25378),
            .lcout(),
            .ltout(n23858_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_1912_LC_10_18_3.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_1912_LC_10_18_3.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_1912_LC_10_18_3.LUT_INIT=16'b1110001011110000;
    LogicCell40 i24_3_lut_4_lut_adj_1912_LC_10_18_3 (
            .in0(N__25372),
            .in1(N__26782),
            .in2(N__25363),
            .in3(N__25637),
            .lcout(n10_adj_4533),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__2__5451_LC_10_18_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__2__5451_LC_10_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__2__5451_LC_10_18_4 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_9__2__5451_LC_10_18_4  (
            .in0(N__49445),
            .in1(N__48846),
            .in2(N__53476),
            .in3(N__25483),
            .lcout(data_out_frame_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66792),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_LC_10_18_5.C_ON=1'b0;
    defparam i24_3_lut_4_lut_LC_10_18_5.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_LC_10_18_5.LUT_INIT=16'b1011101010001010;
    LogicCell40 i24_3_lut_4_lut_LC_10_18_5 (
            .in0(N__26683),
            .in1(N__26781),
            .in2(N__25639),
            .in3(N__28651),
            .lcout(n10_adj_4535),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_2__I_0_i4_3_lut_LC_10_18_6 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_2__I_0_i4_3_lut_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Bit_Index_2__I_0_i4_3_lut_LC_10_18_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Bit_Index_2__I_0_i4_3_lut_LC_10_18_6  (
            .in0(N__30432),
            .in1(N__25522),
            .in2(_gnd_net_),
            .in3(N__25507),
            .lcout(n4_adj_4554),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i3_LC_10_19_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i3_LC_10_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i3_LC_10_19_0 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \c0.tx.r_Tx_Data_i3_LC_10_19_0  (
            .in0(N__27055),
            .in1(N__25489),
            .in2(N__27342),
            .in3(N__29135),
            .lcout(r_Tx_Data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66802),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i5_3_lut_LC_10_19_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i5_3_lut_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i5_3_lut_LC_10_19_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_0_i5_3_lut_LC_10_19_1  (
            .in0(N__25458),
            .in1(N__25449),
            .in2(_gnd_net_),
            .in3(N__39777),
            .lcout(\c0.n5_adj_4422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n24177_bdd_4_lut_LC_10_19_3 .C_ON=1'b0;
    defparam \c0.n24177_bdd_4_lut_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.n24177_bdd_4_lut_LC_10_19_3 .LUT_INIT=16'b1010101011011000;
    LogicCell40 \c0.n24177_bdd_4_lut_LC_10_19_3  (
            .in0(N__28996),
            .in1(N__25482),
            .in2(N__39943),
            .in3(N__36896),
            .lcout(),
            .ltout(\c0.n24180_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20408_4_lut_LC_10_19_4 .C_ON=1'b0;
    defparam \c0.i20408_4_lut_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i20408_4_lut_LC_10_19_4 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.i20408_4_lut_LC_10_19_4  (
            .in0(N__36897),
            .in1(N__30097),
            .in2(N__25471),
            .in3(N__33963),
            .lcout(n24106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__0__5469_LC_10_19_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__0__5469_LC_10_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__0__5469_LC_10_19_5 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_7__0__5469_LC_10_19_5  (
            .in0(N__49415),
            .in1(N__48970),
            .in2(N__25462),
            .in3(N__39115),
            .lcout(data_out_frame_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66802),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__0__5477_LC_10_19_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__0__5477_LC_10_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__0__5477_LC_10_19_7 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_6__0__5477_LC_10_19_7  (
            .in0(N__49414),
            .in1(N__48969),
            .in2(N__39334),
            .in3(N__25450),
            .lcout(data_out_frame_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66802),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i7_LC_10_20_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i7_LC_10_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i7_LC_10_20_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.tx.r_Tx_Data_i7_LC_10_20_0  (
            .in0(N__27330),
            .in1(N__29153),
            .in2(N__27070),
            .in3(N__25675),
            .lcout(r_Tx_Data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66812),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20155_4_lut_LC_10_20_1 .C_ON=1'b0;
    defparam \c0.i20155_4_lut_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i20155_4_lut_LC_10_20_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.i20155_4_lut_LC_10_20_1  (
            .in0(N__25660),
            .in1(N__36899),
            .in2(N__25654),
            .in3(N__33967),
            .lcout(),
            .ltout(\c0.n23850_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20157_4_lut_LC_10_20_2 .C_ON=1'b0;
    defparam \c0.i20157_4_lut_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i20157_4_lut_LC_10_20_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \c0.i20157_4_lut_LC_10_20_2  (
            .in0(N__26783),
            .in1(N__26873),
            .in2(N__25645),
            .in3(N__28243),
            .lcout(),
            .ltout(n23852_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_1914_LC_10_20_3.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_1914_LC_10_20_3.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_1914_LC_10_20_3.LUT_INIT=16'b1110001011110000;
    LogicCell40 i24_3_lut_4_lut_adj_1914_LC_10_20_3 (
            .in0(N__25546),
            .in1(N__26784),
            .in2(N__25642),
            .in3(N__25633),
            .lcout(),
            .ltout(n10_adj_4537_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i0_LC_10_20_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i0_LC_10_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i0_LC_10_20_4 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \c0.tx.r_Tx_Data_i0_LC_10_20_4  (
            .in0(N__27329),
            .in1(N__29152),
            .in2(N__25549),
            .in3(N__25539),
            .lcout(r_Tx_Data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66812),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20412_4_lut_LC_10_20_5 .C_ON=1'b0;
    defparam \c0.i20412_4_lut_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20412_4_lut_LC_10_20_5 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.i20412_4_lut_LC_10_20_5  (
            .in0(N__27139),
            .in1(N__36898),
            .in2(N__26197),
            .in3(N__33966),
            .lcout(n24110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n24195_bdd_4_lut_LC_10_20_7.C_ON=1'b0;
    defparam n24195_bdd_4_lut_LC_10_20_7.SEQ_MODE=4'b0000;
    defparam n24195_bdd_4_lut_LC_10_20_7.LUT_INIT=16'b1110111001010000;
    LogicCell40 n24195_bdd_4_lut_LC_10_20_7 (
            .in0(N__26966),
            .in1(N__27009),
            .in2(N__25540),
            .in3(N__25528),
            .lcout(n24198),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i0_LC_10_21_0 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i0_LC_10_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i0_LC_10_21_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i0_LC_10_21_0  (
            .in0(N__30929),
            .in1(N__41485),
            .in2(_gnd_net_),
            .in3(N__30910),
            .lcout(\c0.tx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66824),
            .ce(),
            .sr(_gnd_net_));
    defparam i13175_3_lut_LC_10_21_2.C_ON=1'b0;
    defparam i13175_3_lut_LC_10_21_2.SEQ_MODE=4'b0000;
    defparam i13175_3_lut_LC_10_21_2.LUT_INIT=16'b0110011010101010;
    LogicCell40 i13175_3_lut_LC_10_21_2 (
            .in0(N__27041),
            .in1(N__26987),
            .in2(_gnd_net_),
            .in3(N__29199),
            .lcout(n16706),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20402_4_lut_LC_10_21_3.C_ON=1'b0;
    defparam i20402_4_lut_LC_10_21_3.SEQ_MODE=4'b0000;
    defparam i20402_4_lut_LC_10_21_3.LUT_INIT=16'b0111010100000000;
    LogicCell40 i20402_4_lut_LC_10_21_3 (
            .in0(N__29200),
            .in1(N__30451),
            .in2(N__30736),
            .in3(N__27042),
            .lcout(),
            .ltout(n24100_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i2_LC_10_21_4 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i2_LC_10_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i2_LC_10_21_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \c0.tx.r_Bit_Index_i2_LC_10_21_4  (
            .in0(N__30452),
            .in1(N__30735),
            .in2(N__25708),
            .in3(N__25705),
            .lcout(r_Bit_Index_2_adj_4551),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66824),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i20364_4_lut_LC_10_21_5 .C_ON=1'b0;
    defparam \c0.tx.i20364_4_lut_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i20364_4_lut_LC_10_21_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx.i20364_4_lut_LC_10_21_5  (
            .in0(N__26988),
            .in1(N__27040),
            .in2(N__30661),
            .in3(N__30450),
            .lcout(),
            .ltout(\c0.tx.n23985_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i28_3_lut_LC_10_21_6 .C_ON=1'b0;
    defparam \c0.tx.i28_3_lut_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i28_3_lut_LC_10_21_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \c0.tx.i28_3_lut_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(N__39274),
            .in2(N__25699),
            .in3(N__30731),
            .lcout(),
            .ltout(\c0.tx.n31_adj_4216_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i0_LC_10_21_7 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i0_LC_10_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i0_LC_10_21_7 .LUT_INIT=16'b0001000001010100;
    LogicCell40 \c0.tx.r_SM_Main_i0_LC_10_21_7  (
            .in0(N__41484),
            .in1(N__33734),
            .in2(N__25696),
            .in3(N__30660),
            .lcout(\c0.tx.r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66824),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_2_lut_LC_10_22_0 .C_ON=1'b1;
    defparam \quad_counter0.add_86_2_lut_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_2_lut_LC_10_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_86_2_lut_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__27602),
            .in2(_gnd_net_),
            .in3(N__25687),
            .lcout(n187),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(\quad_counter0.n19473 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i1_LC_10_22_1 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i1_LC_10_22_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i1_LC_10_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i1_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__27481),
            .in2(_gnd_net_),
            .in3(N__25684),
            .lcout(\quad_counter0.b_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter0.n19473 ),
            .carryout(\quad_counter0.n19474 ),
            .clk(N__66836),
            .ce(N__25803),
            .sr(N__25776));
    defparam \quad_counter0.b_delay_counter__i2_LC_10_22_2 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i2_LC_10_22_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i2_LC_10_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i2_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(N__27468),
            .in2(_gnd_net_),
            .in3(N__25681),
            .lcout(\quad_counter0.b_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter0.n19474 ),
            .carryout(\quad_counter0.n19475 ),
            .clk(N__66836),
            .ce(N__25803),
            .sr(N__25776));
    defparam \quad_counter0.b_delay_counter__i3_LC_10_22_3 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i3_LC_10_22_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i3_LC_10_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i3_LC_10_22_3  (
            .in0(_gnd_net_),
            .in1(N__27646),
            .in2(_gnd_net_),
            .in3(N__25678),
            .lcout(\quad_counter0.b_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter0.n19475 ),
            .carryout(\quad_counter0.n19476 ),
            .clk(N__66836),
            .ce(N__25803),
            .sr(N__25776));
    defparam \quad_counter0.b_delay_counter__i4_LC_10_22_4 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i4_LC_10_22_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i4_LC_10_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i4_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(N__27621),
            .in2(_gnd_net_),
            .in3(N__25735),
            .lcout(\quad_counter0.b_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter0.n19476 ),
            .carryout(\quad_counter0.n19477 ),
            .clk(N__66836),
            .ce(N__25803),
            .sr(N__25776));
    defparam \quad_counter0.b_delay_counter__i5_LC_10_22_5 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i5_LC_10_22_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i5_LC_10_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i5_LC_10_22_5  (
            .in0(_gnd_net_),
            .in1(N__27454),
            .in2(_gnd_net_),
            .in3(N__25732),
            .lcout(\quad_counter0.b_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter0.n19477 ),
            .carryout(\quad_counter0.n19478 ),
            .clk(N__66836),
            .ce(N__25803),
            .sr(N__25776));
    defparam \quad_counter0.b_delay_counter__i6_LC_10_22_6 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i6_LC_10_22_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i6_LC_10_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i6_LC_10_22_6  (
            .in0(_gnd_net_),
            .in1(N__27403),
            .in2(_gnd_net_),
            .in3(N__25729),
            .lcout(\quad_counter0.b_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter0.n19478 ),
            .carryout(\quad_counter0.n19479 ),
            .clk(N__66836),
            .ce(N__25803),
            .sr(N__25776));
    defparam \quad_counter0.b_delay_counter__i7_LC_10_22_7 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i7_LC_10_22_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i7_LC_10_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i7_LC_10_22_7  (
            .in0(_gnd_net_),
            .in1(N__34101),
            .in2(_gnd_net_),
            .in3(N__25726),
            .lcout(\quad_counter0.b_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter0.n19479 ),
            .carryout(\quad_counter0.n19480 ),
            .clk(N__66836),
            .ce(N__25803),
            .sr(N__25776));
    defparam \quad_counter0.b_delay_counter__i8_LC_10_23_0 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i8_LC_10_23_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i8_LC_10_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i8_LC_10_23_0  (
            .in0(_gnd_net_),
            .in1(N__27417),
            .in2(_gnd_net_),
            .in3(N__25723),
            .lcout(\quad_counter0.b_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_10_23_0_),
            .carryout(\quad_counter0.n19481 ),
            .clk(N__66847),
            .ce(N__25804),
            .sr(N__25780));
    defparam \quad_counter0.b_delay_counter__i9_LC_10_23_1 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i9_LC_10_23_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i9_LC_10_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i9_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(N__27634),
            .in2(_gnd_net_),
            .in3(N__25720),
            .lcout(\quad_counter0.b_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter0.n19481 ),
            .carryout(\quad_counter0.n19482 ),
            .clk(N__66847),
            .ce(N__25804),
            .sr(N__25780));
    defparam \quad_counter0.b_delay_counter__i10_LC_10_23_2 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i10_LC_10_23_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i10_LC_10_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i10_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(N__27430),
            .in2(_gnd_net_),
            .in3(N__25717),
            .lcout(\quad_counter0.b_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter0.n19482 ),
            .carryout(\quad_counter0.n19483 ),
            .clk(N__66847),
            .ce(N__25804),
            .sr(N__25780));
    defparam \quad_counter0.b_delay_counter__i11_LC_10_23_3 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i11_LC_10_23_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i11_LC_10_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i11_LC_10_23_3  (
            .in0(_gnd_net_),
            .in1(N__27442),
            .in2(_gnd_net_),
            .in3(N__25714),
            .lcout(\quad_counter0.b_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter0.n19483 ),
            .carryout(\quad_counter0.n19484 ),
            .clk(N__66847),
            .ce(N__25804),
            .sr(N__25780));
    defparam \quad_counter0.b_delay_counter__i12_LC_10_23_4 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i12_LC_10_23_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i12_LC_10_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i12_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(N__34080),
            .in2(_gnd_net_),
            .in3(N__25711),
            .lcout(\quad_counter0.b_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter0.n19484 ),
            .carryout(\quad_counter0.n19485 ),
            .clk(N__66847),
            .ce(N__25804),
            .sr(N__25780));
    defparam \quad_counter0.b_delay_counter__i13_LC_10_23_5 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i13_LC_10_23_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i13_LC_10_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i13_LC_10_23_5  (
            .in0(_gnd_net_),
            .in1(N__27493),
            .in2(_gnd_net_),
            .in3(N__25813),
            .lcout(\quad_counter0.b_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter0.n19485 ),
            .carryout(\quad_counter0.n19486 ),
            .clk(N__66847),
            .ce(N__25804),
            .sr(N__25780));
    defparam \quad_counter0.b_delay_counter__i14_LC_10_23_6 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i14_LC_10_23_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i14_LC_10_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i14_LC_10_23_6  (
            .in0(_gnd_net_),
            .in1(N__34119),
            .in2(_gnd_net_),
            .in3(N__25810),
            .lcout(\quad_counter0.b_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter0.n19486 ),
            .carryout(\quad_counter0.n19487 ),
            .clk(N__66847),
            .ce(N__25804),
            .sr(N__25780));
    defparam \quad_counter0.b_delay_counter__i15_LC_10_23_7 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i15_LC_10_23_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i15_LC_10_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i15_LC_10_23_7  (
            .in0(_gnd_net_),
            .in1(N__34062),
            .in2(_gnd_net_),
            .in3(N__25807),
            .lcout(\quad_counter0.b_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66847),
            .ce(N__25804),
            .sr(N__25780));
    defparam \quad_counter0.add_85_2_lut_LC_10_24_0 .C_ON=1'b1;
    defparam \quad_counter0.add_85_2_lut_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_85_2_lut_LC_10_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_85_2_lut_LC_10_24_0  (
            .in0(_gnd_net_),
            .in1(N__27714),
            .in2(_gnd_net_),
            .in3(N__25753),
            .lcout(n39),
            .ltout(),
            .carryin(bfn_10_24_0_),
            .carryout(\quad_counter0.n19488 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_delay_counter__i1_LC_10_24_1 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i1_LC_10_24_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i1_LC_10_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i1_LC_10_24_1  (
            .in0(_gnd_net_),
            .in1(N__27919),
            .in2(_gnd_net_),
            .in3(N__25750),
            .lcout(\quad_counter0.a_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter0.n19488 ),
            .carryout(\quad_counter0.n19489 ),
            .clk(N__66857),
            .ce(N__27772),
            .sr(N__27747));
    defparam \quad_counter0.a_delay_counter__i2_LC_10_24_2 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i2_LC_10_24_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i2_LC_10_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i2_LC_10_24_2  (
            .in0(_gnd_net_),
            .in1(N__27933),
            .in2(_gnd_net_),
            .in3(N__25747),
            .lcout(\quad_counter0.a_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter0.n19489 ),
            .carryout(\quad_counter0.n19490 ),
            .clk(N__66857),
            .ce(N__27772),
            .sr(N__27747));
    defparam \quad_counter0.a_delay_counter__i3_LC_10_24_3 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i3_LC_10_24_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i3_LC_10_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i3_LC_10_24_3  (
            .in0(_gnd_net_),
            .in1(N__27958),
            .in2(_gnd_net_),
            .in3(N__25744),
            .lcout(\quad_counter0.a_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter0.n19490 ),
            .carryout(\quad_counter0.n19491 ),
            .clk(N__66857),
            .ce(N__27772),
            .sr(N__27747));
    defparam \quad_counter0.a_delay_counter__i4_LC_10_24_4 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i4_LC_10_24_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i4_LC_10_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i4_LC_10_24_4  (
            .in0(_gnd_net_),
            .in1(N__27882),
            .in2(_gnd_net_),
            .in3(N__25741),
            .lcout(\quad_counter0.a_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter0.n19491 ),
            .carryout(\quad_counter0.n19492 ),
            .clk(N__66857),
            .ce(N__27772),
            .sr(N__27747));
    defparam \quad_counter0.a_delay_counter__i5_LC_10_24_5 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i5_LC_10_24_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i5_LC_10_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i5_LC_10_24_5  (
            .in0(_gnd_net_),
            .in1(N__27907),
            .in2(_gnd_net_),
            .in3(N__25738),
            .lcout(\quad_counter0.a_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter0.n19492 ),
            .carryout(\quad_counter0.n19493 ),
            .clk(N__66857),
            .ce(N__27772),
            .sr(N__27747));
    defparam \quad_counter0.a_delay_counter__i6_LC_10_24_6 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i6_LC_10_24_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i6_LC_10_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i6_LC_10_24_6  (
            .in0(_gnd_net_),
            .in1(N__28098),
            .in2(_gnd_net_),
            .in3(N__25840),
            .lcout(\quad_counter0.a_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter0.n19493 ),
            .carryout(\quad_counter0.n19494 ),
            .clk(N__66857),
            .ce(N__27772),
            .sr(N__27747));
    defparam \quad_counter0.a_delay_counter__i7_LC_10_24_7 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i7_LC_10_24_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i7_LC_10_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i7_LC_10_24_7  (
            .in0(_gnd_net_),
            .in1(N__27672),
            .in2(_gnd_net_),
            .in3(N__25837),
            .lcout(\quad_counter0.a_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter0.n19494 ),
            .carryout(\quad_counter0.n19495 ),
            .clk(N__66857),
            .ce(N__27772),
            .sr(N__27747));
    defparam \quad_counter0.a_delay_counter__i8_LC_10_25_0 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i8_LC_10_25_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i8_LC_10_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i8_LC_10_25_0  (
            .in0(_gnd_net_),
            .in1(N__27946),
            .in2(_gnd_net_),
            .in3(N__25834),
            .lcout(\quad_counter0.a_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_10_25_0_),
            .carryout(\quad_counter0.n19496 ),
            .clk(N__66865),
            .ce(N__27768),
            .sr(N__27748));
    defparam \quad_counter0.a_delay_counter__i9_LC_10_25_1 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i9_LC_10_25_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i9_LC_10_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i9_LC_10_25_1  (
            .in0(_gnd_net_),
            .in1(N__28084),
            .in2(_gnd_net_),
            .in3(N__25831),
            .lcout(\quad_counter0.a_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter0.n19496 ),
            .carryout(\quad_counter0.n19497 ),
            .clk(N__66865),
            .ce(N__27768),
            .sr(N__27748));
    defparam \quad_counter0.a_delay_counter__i10_LC_10_25_2 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i10_LC_10_25_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i10_LC_10_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i10_LC_10_25_2  (
            .in0(_gnd_net_),
            .in1(N__27658),
            .in2(_gnd_net_),
            .in3(N__25828),
            .lcout(\quad_counter0.a_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter0.n19497 ),
            .carryout(\quad_counter0.n19498 ),
            .clk(N__66865),
            .ce(N__27768),
            .sr(N__27748));
    defparam \quad_counter0.a_delay_counter__i11_LC_10_25_3 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i11_LC_10_25_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i11_LC_10_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i11_LC_10_25_3  (
            .in0(_gnd_net_),
            .in1(N__27895),
            .in2(_gnd_net_),
            .in3(N__25825),
            .lcout(\quad_counter0.a_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter0.n19498 ),
            .carryout(\quad_counter0.n19499 ),
            .clk(N__66865),
            .ce(N__27768),
            .sr(N__27748));
    defparam \quad_counter0.a_delay_counter__i12_LC_10_25_4 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i12_LC_10_25_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i12_LC_10_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i12_LC_10_25_4  (
            .in0(_gnd_net_),
            .in1(N__28123),
            .in2(_gnd_net_),
            .in3(N__25822),
            .lcout(\quad_counter0.a_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter0.n19499 ),
            .carryout(\quad_counter0.n19500 ),
            .clk(N__66865),
            .ce(N__27768),
            .sr(N__27748));
    defparam \quad_counter0.a_delay_counter__i13_LC_10_25_5 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i13_LC_10_25_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i13_LC_10_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i13_LC_10_25_5  (
            .in0(_gnd_net_),
            .in1(N__28111),
            .in2(_gnd_net_),
            .in3(N__25819),
            .lcout(\quad_counter0.a_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter0.n19500 ),
            .carryout(\quad_counter0.n19501 ),
            .clk(N__66865),
            .ce(N__27768),
            .sr(N__27748));
    defparam \quad_counter0.a_delay_counter__i14_LC_10_25_6 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i14_LC_10_25_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i14_LC_10_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i14_LC_10_25_6  (
            .in0(_gnd_net_),
            .in1(N__27697),
            .in2(_gnd_net_),
            .in3(N__25816),
            .lcout(\quad_counter0.a_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter0.n19501 ),
            .carryout(\quad_counter0.n19502 ),
            .clk(N__66865),
            .ce(N__27768),
            .sr(N__27748));
    defparam \quad_counter0.a_delay_counter__i15_LC_10_25_7 .C_ON=1'b0;
    defparam \quad_counter0.a_delay_counter__i15_LC_10_25_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i15_LC_10_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i15_LC_10_25_7  (
            .in0(_gnd_net_),
            .in1(N__27685),
            .in2(_gnd_net_),
            .in3(N__25888),
            .lcout(\quad_counter0.a_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66865),
            .ce(N__27768),
            .sr(N__27748));
    defparam \c0.i1_2_lut_3_lut_adj_1876_LC_11_7_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1876_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1876_LC_11_7_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1876_LC_11_7_5  (
            .in0(N__31485),
            .in1(N__29564),
            .in2(_gnd_net_),
            .in3(N__34426),
            .lcout(\c0.n22317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_LC_11_8_0 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_LC_11_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i4_2_lut_3_lut_LC_11_8_0  (
            .in0(N__32792),
            .in1(N__35057),
            .in2(_gnd_net_),
            .in3(N__29788),
            .lcout(),
            .ltout(\c0.n18_adj_4414_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1805_LC_11_8_1 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1805_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1805_LC_11_8_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1805_LC_11_8_1  (
            .in0(N__31489),
            .in1(N__25885),
            .in2(N__25879),
            .in3(N__28189),
            .lcout(\c0.n26_adj_4504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1396_LC_11_8_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1396_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1396_LC_11_8_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_3_lut_adj_1396_LC_11_8_3  (
            .in0(N__32565),
            .in1(N__32516),
            .in2(_gnd_net_),
            .in3(N__34828),
            .lcout(),
            .ltout(\c0.n23550_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1804_LC_11_8_4 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1804_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1804_LC_11_8_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_1804_LC_11_8_4  (
            .in0(N__25876),
            .in1(N__34476),
            .in2(N__25870),
            .in3(N__31798),
            .lcout(),
            .ltout(\c0.n22_adj_4503_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__1__5292_LC_11_8_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__1__5292_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__1__5292_LC_11_8_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_29__1__5292_LC_11_8_5  (
            .in0(N__28012),
            .in1(N__29292),
            .in2(N__25867),
            .in3(N__25864),
            .lcout(\c0.data_out_frame_29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66659),
            .ce(N__40953),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_11_9_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_11_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_11_9_0  (
            .in0(N__26148),
            .in1(N__26119),
            .in2(_gnd_net_),
            .in3(N__39835),
            .lcout(\c0.n26_adj_4517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1408_LC_11_9_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1408_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1408_LC_11_9_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_3_lut_adj_1408_LC_11_9_1  (
            .in0(N__32039),
            .in1(N__32790),
            .in2(_gnd_net_),
            .in3(N__31964),
            .lcout(\c0.n10462 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1400_LC_11_9_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1400_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1400_LC_11_9_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1400_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__31927),
            .in2(_gnd_net_),
            .in3(N__32115),
            .lcout(),
            .ltout(\c0.n21305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__2__5299_LC_11_9_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__2__5299_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__2__5299_LC_11_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_28__2__5299_LC_11_9_3  (
            .in0(N__26113),
            .in1(N__28035),
            .in2(N__26122),
            .in3(N__29562),
            .lcout(\c0.data_out_frame_28_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66664),
            .ce(N__40951),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1889_LC_11_9_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1889_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1889_LC_11_9_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1889_LC_11_9_4  (
            .in0(N__32149),
            .in1(N__29353),
            .in2(_gnd_net_),
            .in3(N__32206),
            .lcout(\c0.n6_adj_4515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1870_LC_11_9_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1870_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1870_LC_11_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1870_LC_11_9_5  (
            .in0(N__28171),
            .in1(N__32791),
            .in2(N__32046),
            .in3(N__32517),
            .lcout(\c0.n12532 ),
            .ltout(\c0.n12532_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1641_LC_11_9_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1641_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1641_LC_11_9_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1641_LC_11_9_6  (
            .in0(N__29423),
            .in1(_gnd_net_),
            .in2(N__26104),
            .in3(N__32205),
            .lcout(\c0.n22126 ),
            .ltout(\c0.n22126_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__4__5297_LC_11_9_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__4__5297_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__4__5297_LC_11_9_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.data_out_frame_28__4__5297_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__31840),
            .in2(N__26101),
            .in3(N__34850),
            .lcout(\c0.data_out_frame_28_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66664),
            .ce(N__40951),
            .sr(_gnd_net_));
    defparam \quad_counter1.i10_4_lut_LC_11_10_0 .C_ON=1'b0;
    defparam \quad_counter1.i10_4_lut_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i10_4_lut_LC_11_10_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i10_4_lut_LC_11_10_0  (
            .in0(N__26086),
            .in1(N__26070),
            .in2(N__26059),
            .in3(N__26043),
            .lcout(\quad_counter1.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.quadA_I_0_73_2_lut_LC_11_10_1 .C_ON=1'b0;
    defparam \quad_counter1.quadA_I_0_73_2_lut_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.quadA_I_0_73_2_lut_LC_11_10_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \quad_counter1.quadA_I_0_73_2_lut_LC_11_10_1  (
            .in0(N__25966),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25991),
            .lcout(a_delay_counter_15__N_4124_adj_4547),
            .ltout(a_delay_counter_15__N_4124_adj_4547_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_11_10_2.C_ON=1'b0;
    defparam i1_4_lut_LC_11_10_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_11_10_2.LUT_INIT=16'b1111100111110000;
    LogicCell40 i1_4_lut_LC_11_10_2 (
            .in0(N__25992),
            .in1(N__25965),
            .in2(N__25921),
            .in3(N__25918),
            .lcout(n14228),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_2_lut_LC_11_10_5 .C_ON=1'b0;
    defparam \c0.i14_2_lut_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i14_2_lut_LC_11_10_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i14_2_lut_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__41913),
            .in2(_gnd_net_),
            .in3(N__43079),
            .lcout(\c0.n161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__2__5291_LC_11_10_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__2__5291_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__2__5291_LC_11_10_6 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.data_out_frame_29__2__5291_LC_11_10_6  (
            .in0(N__28269),
            .in1(N__49410),
            .in2(N__26152),
            .in3(N__49019),
            .lcout(data_out_frame_29_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66673),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1724_LC_11_10_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1724_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1724_LC_11_10_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1724_LC_11_10_7  (
            .in0(N__31926),
            .in1(N__32116),
            .in2(N__29377),
            .in3(N__32148),
            .lcout(data_out_frame_28__3__N_1881),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_rx_data_ready_prev_5283_LC_11_11_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_rx_data_ready_prev_5283_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_rx_data_ready_prev_5283_LC_11_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.FRAME_MATCHER_rx_data_ready_prev_5283_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43110),
            .lcout(\c0.FRAME_MATCHER_rx_data_ready_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66684),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_52_LC_11_11_2 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_52_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_DV_52_LC_11_11_2 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \c0.rx.r_Rx_DV_52_LC_11_11_2  (
            .in0(N__57028),
            .in1(N__43111),
            .in2(N__54343),
            .in3(N__56950),
            .lcout(rx_data_ready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66684),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i9_LC_11_11_3 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i9_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i9_LC_11_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i9_LC_11_11_3  (
            .in0(N__38505),
            .in1(N__26137),
            .in2(_gnd_net_),
            .in3(N__32286),
            .lcout(encoder1_position_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66684),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__3__5290_LC_11_11_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__3__5290_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__3__5290_LC_11_11_4 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \c0.data_out_frame_29__3__5290_LC_11_11_4  (
            .in0(N__49569),
            .in1(N__26622),
            .in2(N__49047),
            .in3(N__29293),
            .lcout(data_out_frame_29_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66684),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1454_LC_11_11_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1454_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1454_LC_11_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1454_LC_11_11_5  (
            .in0(N__26482),
            .in1(N__35149),
            .in2(N__28965),
            .in3(N__38870),
            .lcout(\c0.n13079 ),
            .ltout(\c0.n13079_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1413_LC_11_11_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1413_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1413_LC_11_11_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1413_LC_11_11_6  (
            .in0(N__35911),
            .in1(N__26161),
            .in2(N__26125),
            .in3(N__35723),
            .lcout(\c0.n21056 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i3_LC_11_11_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i3_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i3_LC_11_11_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i3_LC_11_11_7  (
            .in0(N__43109),
            .in1(N__30611),
            .in2(_gnd_net_),
            .in3(N__30338),
            .lcout(data_in_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66684),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1407_LC_11_12_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1407_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1407_LC_11_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1407_LC_11_12_0  (
            .in0(N__26335),
            .in1(N__26230),
            .in2(N__26224),
            .in3(N__35839),
            .lcout(\c0.n20175 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_11_12_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_11_12_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_11_12_2  (
            .in0(N__39822),
            .in1(N__26211),
            .in2(_gnd_net_),
            .in3(N__35341),
            .lcout(\c0.n11_adj_4424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1485_LC_11_12_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1485_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1485_LC_11_12_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_1485_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__26334),
            .in2(_gnd_net_),
            .in3(N__35449),
            .lcout(),
            .ltout(\c0.n6_adj_4335_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1486_LC_11_12_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1486_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1486_LC_11_12_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_4_lut_adj_1486_LC_11_12_4  (
            .in0(N__35030),
            .in1(N__28678),
            .in2(N__26179),
            .in3(N__26423),
            .lcout(\c0.n21229 ),
            .ltout(\c0.n21229_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1685_LC_11_12_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1685_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1685_LC_11_12_5 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1685_LC_11_12_5  (
            .in0(N__28311),
            .in1(_gnd_net_),
            .in2(N__26176),
            .in3(N__31256),
            .lcout(\c0.n21152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i12_LC_11_12_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i12_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i12_LC_11_12_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter1.count_i0_i12_LC_11_12_7  (
            .in0(N__34631),
            .in1(N__26173),
            .in2(_gnd_net_),
            .in3(N__38395),
            .lcout(encoder1_position_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66699),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1705_LC_11_13_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1705_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1705_LC_11_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1705_LC_11_13_0  (
            .in0(N__33163),
            .in1(N__26325),
            .in2(N__28786),
            .in3(N__26419),
            .lcout(\c0.n6_adj_4309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__5__5448_LC_11_13_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__5__5448_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__5__5448_LC_11_13_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_9__5__5448_LC_11_13_1  (
            .in0(N__49561),
            .in1(N__48968),
            .in2(N__36082),
            .in3(N__27108),
            .lcout(data_out_frame_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1429_LC_11_13_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1429_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1429_LC_11_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1429_LC_11_13_2  (
            .in0(N__33161),
            .in1(N__26418),
            .in2(_gnd_net_),
            .in3(N__26324),
            .lcout(\c0.n22293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1483_LC_11_13_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1483_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1483_LC_11_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1483_LC_11_13_3  (
            .in0(N__28660),
            .in1(N__35445),
            .in2(N__37072),
            .in3(N__33160),
            .lcout(\c0.n20330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i1_LC_11_13_4 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i1_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i1_LC_11_13_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i1_LC_11_13_4  (
            .in0(N__38497),
            .in1(N__26344),
            .in2(_gnd_net_),
            .in3(N__32789),
            .lcout(encoder1_position_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1414_LC_11_13_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1414_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1414_LC_11_13_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1414_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__35519),
            .in2(_gnd_net_),
            .in3(N__33162),
            .lcout(),
            .ltout(\c0.n6_adj_4310_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1415_LC_11_13_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1415_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1415_LC_11_13_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1415_LC_11_13_6  (
            .in0(N__26481),
            .in1(N__38179),
            .in2(N__26338),
            .in3(N__38875),
            .lcout(\c0.n22037 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__7__5422_LC_11_14_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__7__5422_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__7__5422_LC_11_14_0 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_out_frame_12__7__5422_LC_11_14_0  (
            .in0(N__49002),
            .in1(N__49380),
            .in2(N__26278),
            .in3(N__26326),
            .lcout(data_out_frame_12_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66726),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_11_14_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_11_14_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_11_14_1  (
            .in0(N__32068),
            .in1(N__26274),
            .in2(_gnd_net_),
            .in3(N__39756),
            .lcout(\c0.n11_adj_4360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i8_LC_11_14_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i8_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i8_LC_11_14_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i8_LC_11_14_2  (
            .in0(N__38498),
            .in1(N__26254),
            .in2(_gnd_net_),
            .in3(N__35391),
            .lcout(encoder1_position_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66726),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_11_14_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_11_14_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_11_14_3  (
            .in0(N__26238),
            .in1(N__30388),
            .in2(_gnd_net_),
            .in3(N__39757),
            .lcout(\c0.n5_adj_4227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__4__5465_LC_11_14_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__4__5465_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__4__5465_LC_11_14_4 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_7__4__5465_LC_11_14_4  (
            .in0(N__49004),
            .in1(N__49382),
            .in2(N__36136),
            .in3(N__26239),
            .lcout(data_out_frame_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66726),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__3__5298_LC_11_14_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__3__5298_LC_11_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__3__5298_LC_11_14_6 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_out_frame_28__3__5298_LC_11_14_6  (
            .in0(N__49003),
            .in1(N__49381),
            .in2(N__26608),
            .in3(N__28065),
            .lcout(data_out_frame_28_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66726),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1849_LC_11_14_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1849_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1849_LC_11_14_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1849_LC_11_14_7  (
            .in0(N__39499),
            .in1(N__35418),
            .in2(N__35794),
            .in3(N__38586),
            .lcout(\c0.n10422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.encoder0_position_27__I_0_2_lut_LC_11_15_0 .C_ON=1'b0;
    defparam \c0.encoder0_position_27__I_0_2_lut_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.encoder0_position_27__I_0_2_lut_LC_11_15_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.encoder0_position_27__I_0_2_lut_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__33386),
            .in2(_gnd_net_),
            .in3(N__40056),
            .lcout(\c0.data_out_frame_29__7__N_850 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20186_3_lut_LC_11_15_1 .C_ON=1'b0;
    defparam \c0.i20186_3_lut_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i20186_3_lut_LC_11_15_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i20186_3_lut_LC_11_15_1  (
            .in0(N__26464),
            .in1(N__26379),
            .in2(_gnd_net_),
            .in3(N__39805),
            .lcout(\c0.n23881 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i16_LC_11_15_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i16_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i16_LC_11_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i16_LC_11_15_2  (
            .in0(N__38491),
            .in1(N__26434),
            .in2(_gnd_net_),
            .in3(N__26417),
            .lcout(encoder1_position_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66739),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__4__5441_LC_11_15_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__4__5441_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__4__5441_LC_11_15_3 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_frame_10__4__5441_LC_11_15_3  (
            .in0(N__49553),
            .in1(N__26380),
            .in2(N__36505),
            .in3(N__48939),
            .lcout(data_out_frame_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66739),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i11_LC_11_15_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i11_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i11_LC_11_15_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i11_LC_11_15_4  (
            .in0(N__43154),
            .in1(N__28846),
            .in2(_gnd_net_),
            .in3(N__30328),
            .lcout(data_in_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66739),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__2__5467_LC_11_15_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__2__5467_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__2__5467_LC_11_15_5 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_7__2__5467_LC_11_15_5  (
            .in0(N__49554),
            .in1(N__48938),
            .in2(N__41758),
            .in3(N__26364),
            .lcout(data_out_frame_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66739),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i17_LC_11_15_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i17_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i17_LC_11_15_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \quad_counter1.count_i0_i17_LC_11_15_7  (
            .in0(N__26350),
            .in1(N__37250),
            .in2(_gnd_net_),
            .in3(N__38492),
            .lcout(encoder1_position_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66739),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i19_LC_11_16_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i19_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i19_LC_11_16_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i19_LC_11_16_0  (
            .in0(N__43193),
            .in1(N__28845),
            .in2(_gnd_net_),
            .in3(N__36595),
            .lcout(data_in_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66753),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i21_LC_11_16_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i21_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i21_LC_11_16_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter1.count_i0_i21_LC_11_16_1  (
            .in0(N__28610),
            .in1(N__26644),
            .in2(_gnd_net_),
            .in3(N__38499),
            .lcout(encoder1_position_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66753),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i23_LC_11_16_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i23_LC_11_16_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i23_LC_11_16_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i23_LC_11_16_2  (
            .in0(N__38500),
            .in1(N__26638),
            .in2(_gnd_net_),
            .in3(N__32892),
            .lcout(encoder1_position_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66753),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i29_LC_11_16_3 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i29_LC_11_16_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i29_LC_11_16_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter1.count_i0_i29_LC_11_16_3  (
            .in0(N__28958),
            .in1(N__26632),
            .in2(_gnd_net_),
            .in3(N__38501),
            .lcout(encoder1_position_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66753),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_11_16_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_11_16_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_11_16_4  (
            .in0(N__39807),
            .in1(N__26626),
            .in2(_gnd_net_),
            .in3(N__26607),
            .lcout(\c0.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i30_LC_11_16_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i30_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i30_LC_11_16_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i30_LC_11_16_6  (
            .in0(N__38502),
            .in1(N__26581),
            .in2(_gnd_net_),
            .in3(N__35518),
            .lcout(encoder1_position_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66753),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_11_16_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_11_16_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_11_16_7  (
            .in0(N__26575),
            .in1(N__36286),
            .in2(_gnd_net_),
            .in3(N__39806),
            .lcout(\c0.n5_adj_4346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__3__5474_LC_11_17_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__3__5474_LC_11_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__3__5474_LC_11_17_0 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_6__3__5474_LC_11_17_0  (
            .in0(N__49517),
            .in1(N__49006),
            .in2(N__33394),
            .in3(N__27210),
            .lcout(data_out_frame_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66767),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__7__5446_LC_11_17_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__7__5446_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__7__5446_LC_11_17_1 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_9__7__5446_LC_11_17_1  (
            .in0(N__49005),
            .in1(N__49413),
            .in2(N__33253),
            .in3(N__26541),
            .lcout(data_out_frame_9_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66767),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_45_LC_11_17_3 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_45_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.o_Tx_Serial_45_LC_11_17_3 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \c0.tx.o_Tx_Serial_45_LC_11_17_3  (
            .in0(N__26493),
            .in1(N__30748),
            .in2(_gnd_net_),
            .in3(N__41491),
            .lcout(tx_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66767),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1604_LC_11_17_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1604_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1604_LC_11_17_4 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \c0.i3_4_lut_adj_1604_LC_11_17_4  (
            .in0(N__33864),
            .in1(N__39626),
            .in2(N__36817),
            .in3(N__26938),
            .lcout(),
            .ltout(\c0.n23574_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1675_LC_11_17_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1675_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1675_LC_11_17_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_1675_LC_11_17_5  (
            .in0(N__27310),
            .in1(N__26932),
            .in2(N__26914),
            .in3(N__26911),
            .lcout(\c0.n38_adj_4387 ),
            .ltout(\c0.n38_adj_4387_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20438_2_lut_3_lut_LC_11_17_6 .C_ON=1'b0;
    defparam \c0.i20438_2_lut_3_lut_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i20438_2_lut_3_lut_LC_11_17_6 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \c0.i20438_2_lut_3_lut_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__39273),
            .in2(N__26896),
            .in3(N__37147),
            .lcout(\c0.tx_transmit_N_3651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__5__5456_LC_11_18_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__5__5456_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__5__5456_LC_11_18_0 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_out_frame_8__5__5456_LC_11_18_0  (
            .in0(N__48978),
            .in1(N__49519),
            .in2(N__27091),
            .in3(N__35725),
            .lcout(data_out_frame_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66781),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__5__5432_LC_11_18_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__5__5432_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__5__5432_LC_11_18_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_11__5__5432_LC_11_18_1  (
            .in0(N__49518),
            .in1(N__48979),
            .in2(N__28615),
            .in3(N__27123),
            .lcout(data_out_frame_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66781),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__2__5483_LC_11_18_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__2__5483_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__2__5483_LC_11_18_2 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_out_frame_5__2__5483_LC_11_18_2  (
            .in0(N__48976),
            .in1(N__39487),
            .in2(N__49551),
            .in3(N__26889),
            .lcout(data_out_frame_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66781),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20169_4_lut_LC_11_18_3 .C_ON=1'b0;
    defparam \c0.i20169_4_lut_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i20169_4_lut_LC_11_18_3 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \c0.i20169_4_lut_LC_11_18_3  (
            .in0(N__27991),
            .in1(N__33988),
            .in2(N__26863),
            .in3(N__26779),
            .lcout(n23864),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__6__5479_LC_11_18_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__6__5479_LC_11_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__6__5479_LC_11_18_4 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_out_frame_5__6__5479_LC_11_18_4  (
            .in0(N__48977),
            .in1(N__42307),
            .in2(N__49552),
            .in3(N__26673),
            .lcout(data_out_frame_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66781),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_11_18_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_11_18_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_11_18_5  (
            .in0(N__39749),
            .in1(N__26659),
            .in2(_gnd_net_),
            .in3(N__28911),
            .lcout(\c0.n11_adj_4218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20456_LC_11_18_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20456_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20456_LC_11_18_6 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_20456_LC_11_18_6  (
            .in0(N__36894),
            .in1(N__28929),
            .in2(N__27124),
            .in3(N__39750),
            .lcout(),
            .ltout(\c0.n24141_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n24141_bdd_4_lut_LC_11_18_7 .C_ON=1'b0;
    defparam \c0.n24141_bdd_4_lut_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.n24141_bdd_4_lut_LC_11_18_7 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n24141_bdd_4_lut_LC_11_18_7  (
            .in0(N__36895),
            .in1(N__27112),
            .in2(N__27094),
            .in3(N__27087),
            .lcout(\c0.n24144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Bit_Index_2__bdd_4_lut_20490_LC_11_19_0.C_ON=1'b0;
    defparam r_Bit_Index_2__bdd_4_lut_20490_LC_11_19_0.SEQ_MODE=4'b0000;
    defparam r_Bit_Index_2__bdd_4_lut_20490_LC_11_19_0.LUT_INIT=16'b1010111111000000;
    LogicCell40 r_Bit_Index_2__bdd_4_lut_20490_LC_11_19_0 (
            .in0(N__27066),
            .in1(N__27054),
            .in2(N__26978),
            .in3(N__27043),
            .lcout(),
            .ltout(n24189_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n24189_bdd_4_lut_LC_11_19_1.C_ON=1'b0;
    defparam n24189_bdd_4_lut_LC_11_19_1.SEQ_MODE=4'b0000;
    defparam n24189_bdd_4_lut_LC_11_19_1.LUT_INIT=16'b1111000010101100;
    LogicCell40 n24189_bdd_4_lut_LC_11_19_1 (
            .in0(N__27016),
            .in1(N__27255),
            .in2(N__26992),
            .in3(N__26970),
            .lcout(n24192),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i8_LC_11_19_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i8_LC_11_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i8_LC_11_19_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i8_LC_11_19_2  (
            .in0(N__30502),
            .in1(N__43155),
            .in2(_gnd_net_),
            .in3(N__27245),
            .lcout(data_in_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66793),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i0_LC_11_19_3 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i0_LC_11_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i0_LC_11_19_3 .LUT_INIT=16'b0010001011001100;
    LogicCell40 \c0.tx.r_Bit_Index_i0_LC_11_19_3  (
            .in0(N__30729),
            .in1(N__30443),
            .in2(_gnd_net_),
            .in3(N__29193),
            .lcout(r_Bit_Index_0_adj_4553),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66793),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i1_LC_11_19_4 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i1_LC_11_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i1_LC_11_19_4 .LUT_INIT=16'b0110101000100010;
    LogicCell40 \c0.tx.r_Bit_Index_i1_LC_11_19_4  (
            .in0(N__26971),
            .in1(N__29192),
            .in2(N__30453),
            .in3(N__30730),
            .lcout(r_Bit_Index_1_adj_4552),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66793),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1694_LC_11_19_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1694_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1694_LC_11_19_5 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \c0.i6_4_lut_adj_1694_LC_11_19_5  (
            .in0(N__43045),
            .in1(N__36994),
            .in2(N__27247),
            .in3(N__29069),
            .lcout(\c0.n16_adj_4476 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i1_LC_11_19_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i1_LC_11_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i1_LC_11_19_6 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \c0.tx.r_Tx_Data_i1_LC_11_19_6  (
            .in0(N__27256),
            .in1(N__27352),
            .in2(N__27343),
            .in3(N__29117),
            .lcout(r_Tx_Data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66793),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_LC_11_19_7 .C_ON=1'b0;
    defparam \c0.i6_4_lut_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_LC_11_19_7 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i6_4_lut_LC_11_19_7  (
            .in0(N__43044),
            .in1(N__29068),
            .in2(N__27246),
            .in3(N__30618),
            .lcout(\c0.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1888_LC_11_20_0 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1888_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1888_LC_11_20_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i8_4_lut_adj_1888_LC_11_20_0  (
            .in0(N__43411),
            .in1(N__37799),
            .in2(N__41011),
            .in3(N__34247),
            .lcout(\c0.n20_adj_4482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__3__5482_LC_11_20_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__3__5482_LC_11_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__3__5482_LC_11_20_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_5__3__5482_LC_11_20_1  (
            .in0(N__49549),
            .in1(N__48975),
            .in2(N__41815),
            .in3(N__27228),
            .lcout(data_out_frame_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66803),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_11_20_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_11_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_11_20_3  (
            .in0(N__39799),
            .in1(N__37102),
            .in2(_gnd_net_),
            .in3(N__27211),
            .lcout(\c0.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__5__5480_LC_11_20_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__5__5480_LC_11_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__5__5480_LC_11_20_4 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_out_frame_5__5__5480_LC_11_20_4  (
            .in0(N__48974),
            .in1(N__49550),
            .in2(N__27180),
            .in3(N__40213),
            .lcout(data_out_frame_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66803),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20471_LC_11_20_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20471_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20471_LC_11_20_5 .LUT_INIT=16'b1101100010101010;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_20471_LC_11_20_5  (
            .in0(N__39800),
            .in1(N__27157),
            .in2(N__29089),
            .in3(N__36887),
            .lcout(),
            .ltout(\c0.n24165_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n24165_bdd_4_lut_LC_11_20_6 .C_ON=1'b0;
    defparam \c0.n24165_bdd_4_lut_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.n24165_bdd_4_lut_LC_11_20_6 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n24165_bdd_4_lut_LC_11_20_6  (
            .in0(N__36888),
            .in1(N__34030),
            .in2(N__27142),
            .in3(N__37018),
            .lcout(\c0.n24168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i22_LC_11_21_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i22_LC_11_21_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i22_LC_11_21_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i22_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(N__34302),
            .in2(_gnd_net_),
            .in3(N__52858),
            .lcout(\c0.FRAME_MATCHER_state_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66813),
            .ce(),
            .sr(N__29173));
    defparam \quad_counter0.i3_4_lut_LC_11_22_1 .C_ON=1'b0;
    defparam \quad_counter0.i3_4_lut_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i3_4_lut_LC_11_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \quad_counter0.i3_4_lut_LC_11_22_1  (
            .in0(N__27358),
            .in1(N__27973),
            .in2(N__27868),
            .in3(N__27503),
            .lcout(count_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i9_4_lut_LC_11_22_2 .C_ON=1'b0;
    defparam \quad_counter0.i9_4_lut_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i9_4_lut_LC_11_22_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \quad_counter0.i9_4_lut_LC_11_22_2  (
            .in0(N__27645),
            .in1(N__27633),
            .in2(N__27622),
            .in3(N__27606),
            .lcout(\quad_counter0.n25_adj_4201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1072_1_lut_2_lut_LC_11_22_3 .C_ON=1'b0;
    defparam \quad_counter0.i1072_1_lut_2_lut_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1072_1_lut_2_lut_LC_11_22_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \quad_counter0.i1072_1_lut_2_lut_LC_11_22_3  (
            .in0(_gnd_net_),
            .in1(N__27972),
            .in2(_gnd_net_),
            .in3(N__27864),
            .lcout(\quad_counter0.n2227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.B_65_LC_11_22_4 .C_ON=1'b0;
    defparam \quad_counter0.B_65_LC_11_22_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.B_65_LC_11_22_4 .LUT_INIT=16'b1010101011101000;
    LogicCell40 \quad_counter0.B_65_LC_11_22_4  (
            .in0(N__27504),
            .in1(N__27583),
            .in2(N__27538),
            .in3(N__27372),
            .lcout(B_filtered),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66825),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.B_delayed_68_LC_11_22_6 .C_ON=1'b0;
    defparam \quad_counter0.B_delayed_68_LC_11_22_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.B_delayed_68_LC_11_22_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \quad_counter0.B_delayed_68_LC_11_22_6  (
            .in0(N__27505),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.B_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66825),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i12_4_lut_LC_11_23_0 .C_ON=1'b0;
    defparam \quad_counter0.i12_4_lut_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12_4_lut_LC_11_23_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \quad_counter0.i12_4_lut_LC_11_23_0  (
            .in0(N__27492),
            .in1(N__27480),
            .in2(N__27469),
            .in3(N__27453),
            .lcout(\quad_counter0.n28_adj_4198 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i10_4_lut_LC_11_23_2 .C_ON=1'b0;
    defparam \quad_counter0.i10_4_lut_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i10_4_lut_LC_11_23_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i10_4_lut_LC_11_23_2  (
            .in0(N__27441),
            .in1(N__27429),
            .in2(N__27418),
            .in3(N__27402),
            .lcout(),
            .ltout(\quad_counter0.n26_adj_4199_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i15_4_lut_LC_11_23_3 .C_ON=1'b0;
    defparam \quad_counter0.i15_4_lut_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i15_4_lut_LC_11_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i15_4_lut_LC_11_23_3  (
            .in0(N__27391),
            .in1(N__34048),
            .in2(N__27385),
            .in3(N__27382),
            .lcout(n12909),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.A_delayed_67_LC_11_23_4 .C_ON=1'b0;
    defparam \quad_counter0.A_delayed_67_LC_11_23_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.A_delayed_67_LC_11_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.A_delayed_67_LC_11_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27859),
            .lcout(\quad_counter0.A_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66837),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.A_filtered_I_0_2_lut_LC_11_23_6 .C_ON=1'b0;
    defparam \quad_counter0.A_filtered_I_0_2_lut_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.A_filtered_I_0_2_lut_LC_11_23_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \quad_counter0.A_filtered_I_0_2_lut_LC_11_23_6  (
            .in0(_gnd_net_),
            .in1(N__27971),
            .in2(_gnd_net_),
            .in3(N__27858),
            .lcout(\quad_counter0.count_direction ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i12_4_lut_adj_1161_LC_11_24_1 .C_ON=1'b0;
    defparam \quad_counter0.i12_4_lut_adj_1161_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12_4_lut_adj_1161_LC_11_24_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \quad_counter0.i12_4_lut_adj_1161_LC_11_24_1  (
            .in0(N__27957),
            .in1(N__27945),
            .in2(N__27934),
            .in3(N__27918),
            .lcout(\quad_counter0.n28_adj_4202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i9_4_lut_adj_1164_LC_11_24_2 .C_ON=1'b0;
    defparam \quad_counter0.i9_4_lut_adj_1164_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i9_4_lut_adj_1164_LC_11_24_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \quad_counter0.i9_4_lut_adj_1164_LC_11_24_2  (
            .in0(N__27906),
            .in1(N__27894),
            .in2(N__27883),
            .in3(N__27713),
            .lcout(\quad_counter0.n25_adj_4205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.A_63_LC_11_24_3 .C_ON=1'b0;
    defparam \quad_counter0.A_63_LC_11_24_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.A_63_LC_11_24_3 .LUT_INIT=16'b1111111001000000;
    LogicCell40 \quad_counter0.A_63_LC_11_24_3  (
            .in0(N__28132),
            .in1(N__27832),
            .in2(N__27799),
            .in3(N__27863),
            .lcout(A_filtered),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66848),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1764_LC_11_24_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1764_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1764_LC_11_24_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1764_LC_11_24_4  (
            .in0(N__53012),
            .in1(N__37846),
            .in2(_gnd_net_),
            .in3(N__53195),
            .lcout(\c0.n21362 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_11_24_6.C_ON=1'b0;
    defparam i1_3_lut_LC_11_24_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_11_24_6.LUT_INIT=16'b1111111101100110;
    LogicCell40 i1_3_lut_LC_11_24_6 (
            .in0(N__27831),
            .in1(N__27795),
            .in2(_gnd_net_),
            .in3(N__28131),
            .lcout(n14421),
            .ltout(n14421_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_delay_counter__i0_LC_11_24_7 .C_ON=1'b0;
    defparam \quad_counter0.a_delay_counter__i0_LC_11_24_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i0_LC_11_24_7 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \quad_counter0.a_delay_counter__i0_LC_11_24_7  (
            .in0(N__27746),
            .in1(N__27724),
            .in2(N__27718),
            .in3(N__27715),
            .lcout(a_delay_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66848),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i11_4_lut_adj_1163_LC_11_25_4 .C_ON=1'b0;
    defparam \quad_counter0.i11_4_lut_adj_1163_LC_11_25_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i11_4_lut_adj_1163_LC_11_25_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i11_4_lut_adj_1163_LC_11_25_4  (
            .in0(N__27696),
            .in1(N__27684),
            .in2(N__27673),
            .in3(N__27657),
            .lcout(),
            .ltout(\quad_counter0.n27_adj_4204_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i15_4_lut_adj_1165_LC_11_25_5 .C_ON=1'b0;
    defparam \quad_counter0.i15_4_lut_adj_1165_LC_11_25_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i15_4_lut_adj_1165_LC_11_25_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i15_4_lut_adj_1165_LC_11_25_5  (
            .in0(N__28147),
            .in1(N__28072),
            .in2(N__28141),
            .in3(N__28138),
            .lcout(n9821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i10_4_lut_adj_1162_LC_11_25_7 .C_ON=1'b0;
    defparam \quad_counter0.i10_4_lut_adj_1162_LC_11_25_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i10_4_lut_adj_1162_LC_11_25_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i10_4_lut_adj_1162_LC_11_25_7  (
            .in0(N__28122),
            .in1(N__28110),
            .in2(N__28099),
            .in3(N__28083),
            .lcout(\quad_counter0.n26_adj_4203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__1__5300_LC_12_6_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__1__5300_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__1__5300_LC_12_6_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame_28__1__5300_LC_12_6_4  (
            .in0(N__28066),
            .in1(N__30981),
            .in2(N__28042),
            .in3(N__29215),
            .lcout(\c0.data_out_frame_28_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66638),
            .ce(N__40952),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1801_LC_12_7_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1801_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1801_LC_12_7_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1801_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__31458),
            .in2(_gnd_net_),
            .in3(N__32212),
            .lcout(\c0.n21062 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1582_LC_12_7_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1582_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1582_LC_12_7_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1582_LC_12_7_1  (
            .in0(N__31770),
            .in1(N__29563),
            .in2(N__32389),
            .in3(N__35614),
            .lcout(\c0.n20376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_12_8_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_12_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_12_8_0  (
            .in0(N__28006),
            .in1(N__27997),
            .in2(_gnd_net_),
            .in3(N__39833),
            .lcout(\c0.n26_adj_4519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1864_LC_12_8_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1864_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1864_LC_12_8_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1864_LC_12_8_1  (
            .in0(N__31631),
            .in1(N__29805),
            .in2(N__31420),
            .in3(N__31132),
            .lcout(\c0.n12542 ),
            .ltout(\c0.n12542_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_3_lut_4_lut_LC_12_8_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_3_lut_4_lut_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_3_lut_4_lut_LC_12_8_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_3_lut_4_lut_LC_12_8_2  (
            .in0(N__31683),
            .in1(N__29270),
            .in2(N__27976),
            .in3(N__31632),
            .lcout(),
            .ltout(\c0.n14_adj_4340_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1495_LC_12_8_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1495_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1495_LC_12_8_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_1495_LC_12_8_3  (
            .in0(N__31089),
            .in1(N__29209),
            .in2(N__28192),
            .in3(N__31569),
            .lcout(data_out_frame_29__2__N_1749),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1863_LC_12_8_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1863_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1863_LC_12_8_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1863_LC_12_8_5  (
            .in0(N__29602),
            .in1(N__29804),
            .in2(N__31419),
            .in3(N__31131),
            .lcout(\c0.n20320 ),
            .ltout(\c0.n20320_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1880_LC_12_8_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1880_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1880_LC_12_8_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1880_LC_12_8_6  (
            .in0(N__34399),
            .in1(N__31682),
            .in2(N__28183),
            .in3(N__31415),
            .lcout(\c0.n21219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1845_LC_12_8_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1845_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1845_LC_12_8_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1845_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(N__29354),
            .in2(_gnd_net_),
            .in3(N__29416),
            .lcout(\c0.n21128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1707_LC_12_9_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1707_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1707_LC_12_9_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1707_LC_12_9_0  (
            .in0(N__35122),
            .in1(N__29695),
            .in2(N__28356),
            .in3(N__53386),
            .lcout(\c0.n22180 ),
            .ltout(\c0.n22180_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_4_lut_LC_12_9_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_4_lut_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_4_lut_LC_12_9_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i1_2_lut_4_lut_4_lut_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__28352),
            .in2(N__28180),
            .in3(N__28169),
            .lcout(\c0.n10498 ),
            .ltout(\c0.n10498_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1835_LC_12_9_2 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1835_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1835_LC_12_9_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_1835_LC_12_9_2  (
            .in0(N__28498),
            .in1(N__28153),
            .in2(N__28177),
            .in3(N__32931),
            .lcout(\c0.n21058 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1591_LC_12_9_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1591_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1591_LC_12_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1591_LC_12_9_3  (
            .in0(N__31285),
            .in1(N__31630),
            .in2(N__31348),
            .in3(N__31130),
            .lcout(\c0.n22024 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1840_LC_12_9_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1840_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1840_LC_12_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1840_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__31209),
            .in2(_gnd_net_),
            .in3(N__34344),
            .lcout(\c0.n20253 ),
            .ltout(\c0.n20253_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1834_LC_12_9_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1834_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1834_LC_12_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_1834_LC_12_9_5  (
            .in0(N__28363),
            .in1(N__31839),
            .in2(N__28174),
            .in3(N__28170),
            .lcout(\c0.n15_adj_4513 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1811_LC_12_9_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1811_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1811_LC_12_9_6 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \c0.i1_2_lut_adj_1811_LC_12_9_6  (
            .in0(N__32505),
            .in1(N__29600),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n21998 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1411_LC_12_9_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1411_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1411_LC_12_9_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_1411_LC_12_9_7  (
            .in0(N__53387),
            .in1(_gnd_net_),
            .in2(N__29705),
            .in3(_gnd_net_),
            .lcout(\c0.n22066 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1610_LC_12_10_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1610_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1610_LC_12_10_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1610_LC_12_10_0  (
            .in0(N__28344),
            .in1(N__32035),
            .in2(N__32799),
            .in3(N__31272),
            .lcout(\c0.n10496 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1484_LC_12_10_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1484_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1484_LC_12_10_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1484_LC_12_10_1  (
            .in0(N__31273),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28345),
            .lcout(),
            .ltout(\c0.n21071_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__0__5293_LC_12_10_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__0__5293_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__0__5293_LC_12_10_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame_29__0__5293_LC_12_10_2  (
            .in0(N__28225),
            .in1(N__28255),
            .in2(N__28273),
            .in3(N__28270),
            .lcout(\c0.data_out_frame_29_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66665),
            .ce(N__40944),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1799_LC_12_10_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1799_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1799_LC_12_10_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1799_LC_12_10_3  (
            .in0(N__31438),
            .in1(N__29608),
            .in2(N__32449),
            .in3(N__31152),
            .lcout(\c0.n17_adj_4501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i26_3_lut_LC_12_10_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i26_3_lut_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i26_3_lut_LC_12_10_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_0_i26_3_lut_LC_12_10_4  (
            .in0(N__28249),
            .in1(N__29479),
            .in2(_gnd_net_),
            .in3(N__39834),
            .lcout(\c0.n26_adj_4423 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1798_LC_12_10_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1798_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1798_LC_12_10_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1798_LC_12_10_5  (
            .in0(N__32617),
            .in1(N__32210),
            .in2(N__31349),
            .in3(N__29767),
            .lcout(\c0.n16_adj_4500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1615_LC_12_11_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1615_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1615_LC_12_11_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1615_LC_12_11_0  (
            .in0(N__28392),
            .in1(N__35386),
            .in2(N__28218),
            .in3(N__28489),
            .lcout(),
            .ltout(\c0.n6_adj_4313_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1420_LC_12_11_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1420_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1420_LC_12_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1420_LC_12_11_1  (
            .in0(N__35310),
            .in1(N__34870),
            .in2(N__28375),
            .in3(N__38965),
            .lcout(\c0.n21156 ),
            .ltout(\c0.n21156_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1713_LC_12_11_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1713_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1713_LC_12_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1713_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__29854),
            .in2(N__28372),
            .in3(N__34793),
            .lcout(\c0.n21231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1613_LC_12_11_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1613_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1613_LC_12_11_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_adj_1613_LC_12_11_4  (
            .in0(N__28393),
            .in1(N__28488),
            .in2(N__36078),
            .in3(N__35385),
            .lcout(\c0.n10_adj_4330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1464_LC_12_11_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1464_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1464_LC_12_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1464_LC_12_11_5  (
            .in0(N__32857),
            .in1(N__32823),
            .in2(N__35283),
            .in3(N__28391),
            .lcout(\c0.n21175 ),
            .ltout(\c0.n21175_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1712_LC_12_11_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1712_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1712_LC_12_11_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1712_LC_12_11_6  (
            .in0(N__29829),
            .in1(N__34794),
            .in2(N__28369),
            .in3(N__31151),
            .lcout(\c0.n21150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1423_LC_12_11_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1423_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1423_LC_12_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1423_LC_12_11_7  (
            .in0(N__35309),
            .in1(N__39035),
            .in2(_gnd_net_),
            .in3(N__28624),
            .lcout(\c0.n22991 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1652_LC_12_12_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1652_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1652_LC_12_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1652_LC_12_12_0  (
            .in0(N__29978),
            .in1(N__34622),
            .in2(N__31892),
            .in3(N__35609),
            .lcout(\c0.n20276 ),
            .ltout(\c0.n20276_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1808_LC_12_12_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1808_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1808_LC_12_12_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1808_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28366),
            .in3(N__31257),
            .lcout(\c0.n21116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1674_LC_12_12_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1674_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1674_LC_12_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1674_LC_12_12_2  (
            .in0(N__29980),
            .in1(N__34623),
            .in2(_gnd_net_),
            .in3(N__35610),
            .lcout(),
            .ltout(\c0.n21110_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1886_LC_12_12_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1886_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1886_LC_12_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1886_LC_12_12_3  (
            .in0(N__35120),
            .in1(N__32371),
            .in2(N__28501),
            .in3(N__31886),
            .lcout(\c0.n14_adj_4514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1428_LC_12_12_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1428_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1428_LC_12_12_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1428_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__32273),
            .in2(_gnd_net_),
            .in3(N__28474),
            .lcout(\c0.n22277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i4_LC_12_12_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i4_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i4_LC_12_12_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter1.count_i0_i4_LC_12_12_5  (
            .in0(N__35121),
            .in1(N__38396),
            .in2(_gnd_net_),
            .in3(N__28438),
            .lcout(encoder1_position_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66685),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1394_LC_12_12_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1394_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1394_LC_12_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1394_LC_12_12_6  (
            .in0(N__29977),
            .in1(N__36454),
            .in2(_gnd_net_),
            .in3(N__38063),
            .lcout(\c0.n21065 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1728_LC_12_12_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1728_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1728_LC_12_12_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1728_LC_12_12_7  (
            .in0(N__34621),
            .in1(N__29979),
            .in2(N__32975),
            .in3(N__32856),
            .lcout(\c0.n21166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1449_LC_12_13_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1449_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1449_LC_12_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1449_LC_12_13_2  (
            .in0(N__29664),
            .in1(N__31252),
            .in2(N__32901),
            .in3(N__29998),
            .lcout(\c0.n17_adj_4323 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1839_LC_12_13_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1839_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1839_LC_12_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1839_LC_12_13_3  (
            .in0(N__41872),
            .in1(N__39056),
            .in2(_gnd_net_),
            .in3(N__39495),
            .lcout(\c0.n22102 ),
            .ltout(\c0.n22102_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1451_LC_12_13_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1451_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1451_LC_12_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1451_LC_12_13_4  (
            .in0(N__28422),
            .in1(N__38515),
            .in2(N__28405),
            .in3(N__28402),
            .lcout(),
            .ltout(\c0.n15_adj_4325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1452_LC_12_13_5 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1452_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1452_LC_12_13_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1452_LC_12_13_5  (
            .in0(N__41293),
            .in1(N__31757),
            .in2(N__28396),
            .in3(N__35461),
            .lcout(\c0.n21041 ),
            .ltout(\c0.n21041_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1453_LC_12_13_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1453_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1453_LC_12_13_6 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \c0.i1_2_lut_adj_1453_LC_12_13_6  (
            .in0(N__35369),
            .in1(_gnd_net_),
            .in2(N__28378),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n22361_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1422_LC_12_13_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1422_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1422_LC_12_13_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1422_LC_12_13_7  (
            .in0(N__28633),
            .in1(N__41682),
            .in2(N__28627),
            .in3(N__35932),
            .lcout(\c0.n10_adj_4314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__6__5455_LC_12_14_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__6__5455_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__6__5455_LC_12_14_0 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_8__6__5455_LC_12_14_0  (
            .in0(N__49335),
            .in1(N__49001),
            .in2(N__35899),
            .in3(N__28566),
            .lcout(data_out_frame_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66713),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__1__5460_LC_12_14_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__1__5460_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__1__5460_LC_12_14_1 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_8__1__5460_LC_12_14_1  (
            .in0(N__48999),
            .in1(N__49336),
            .in2(N__38728),
            .in3(N__33474),
            .lcout(data_out_frame_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66713),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1689_LC_12_14_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1689_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1689_LC_12_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1689_LC_12_14_3  (
            .in0(N__28611),
            .in1(N__36558),
            .in2(_gnd_net_),
            .in3(N__38648),
            .lcout(\c0.n22408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i3_LC_12_14_4 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i3_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i3_LC_12_14_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i3_LC_12_14_4  (
            .in0(N__42202),
            .in1(N__33103),
            .in2(_gnd_net_),
            .in3(N__41673),
            .lcout(encoder0_position_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66713),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n24153_bdd_4_lut_LC_12_14_5 .C_ON=1'b0;
    defparam \c0.n24153_bdd_4_lut_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.n24153_bdd_4_lut_LC_12_14_5 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n24153_bdd_4_lut_LC_12_14_5  (
            .in0(N__29898),
            .in1(N__28582),
            .in2(N__28567),
            .in3(N__36908),
            .lcout(\c0.n24156 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__6__5423_LC_12_14_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__6__5423_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__6__5423_LC_12_14_6 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_12__6__5423_LC_12_14_6  (
            .in0(N__49334),
            .in1(N__49000),
            .in2(N__29665),
            .in3(N__28539),
            .lcout(data_out_frame_12_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66713),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1445_LC_12_14_7 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1445_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1445_LC_12_14_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1445_LC_12_14_7  (
            .in0(N__36504),
            .in1(N__29937),
            .in2(N__41683),
            .in3(N__38724),
            .lcout(\c0.n19_adj_4319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__3__5434_LC_12_15_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__3__5434_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__3__5434_LC_12_15_0 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_out_frame_11__3__5434_LC_12_15_0  (
            .in0(N__48945),
            .in1(N__49403),
            .in2(N__28521),
            .in3(N__30029),
            .lcout(data_out_frame_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66727),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i4_LC_12_15_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i4_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i4_LC_12_15_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i4_LC_12_15_1  (
            .in0(N__43192),
            .in1(N__28811),
            .in2(_gnd_net_),
            .in3(N__36382),
            .lcout(data_in_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66727),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i24_LC_12_15_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i24_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i24_LC_12_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i24_LC_12_15_2  (
            .in0(N__38503),
            .in1(N__28690),
            .in2(_gnd_net_),
            .in3(N__29947),
            .lcout(encoder1_position_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66727),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1469_LC_12_15_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1469_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1469_LC_12_15_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1469_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__37060),
            .in2(_gnd_net_),
            .in3(N__35895),
            .lcout(\c0.n22224 ),
            .ltout(\c0.n22224_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1471_LC_12_15_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1471_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1471_LC_12_15_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1471_LC_12_15_4  (
            .in0(N__29042),
            .in1(N__28639),
            .in2(N__28666),
            .in3(N__36028),
            .lcout(\c0.n13349 ),
            .ltout(\c0.n13349_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1482_LC_12_15_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1482_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1482_LC_12_15_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1482_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28663),
            .in3(N__28781),
            .lcout(\c0.n6_adj_4334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1693_LC_12_15_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1693_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1693_LC_12_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1693_LC_12_15_6  (
            .in0(N__44619),
            .in1(N__41871),
            .in2(_gnd_net_),
            .in3(N__41750),
            .lcout(\c0.n22412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i14_LC_12_16_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i14_LC_12_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i14_LC_12_16_0 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_in_0___i14_LC_12_16_0  (
            .in0(N__43219),
            .in1(_gnd_net_),
            .in2(N__28897),
            .in3(N__36426),
            .lcout(data_in_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66740),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20406_4_lut_LC_12_16_1 .C_ON=1'b0;
    defparam \c0.i20406_4_lut_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i20406_4_lut_LC_12_16_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.i20406_4_lut_LC_12_16_1  (
            .in0(N__33460),
            .in1(N__36889),
            .in2(N__34696),
            .in3(N__33968),
            .lcout(n24104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1470_LC_12_16_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1470_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1470_LC_12_16_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1470_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__35772),
            .in2(_gnd_net_),
            .in3(N__38246),
            .lcout(\c0.n22405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__1__5444_LC_12_16_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__1__5444_LC_12_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__1__5444_LC_12_16_5 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_frame_10__1__5444_LC_12_16_5  (
            .in0(N__49391),
            .in1(N__36924),
            .in2(N__33017),
            .in3(N__48891),
            .lcout(data_out_frame_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66740),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__7__5438_LC_12_16_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__7__5438_LC_12_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__7__5438_LC_12_16_6 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_out_frame_10__7__5438_LC_12_16_6  (
            .in0(N__48889),
            .in1(N__49393),
            .in2(N__28741),
            .in3(N__28782),
            .lcout(data_out_frame_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66740),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__7__5454_LC_12_16_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__7__5454_LC_12_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__7__5454_LC_12_16_7 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_8__7__5454_LC_12_16_7  (
            .in0(N__49392),
            .in1(N__48890),
            .in2(N__36265),
            .in3(N__28722),
            .lcout(data_out_frame_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66740),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1547_LC_12_17_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1547_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1547_LC_12_17_0 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i7_4_lut_adj_1547_LC_12_17_0  (
            .in0(N__36427),
            .in1(N__30278),
            .in2(N__36961),
            .in3(N__30580),
            .lcout(\c0.n19_adj_4367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i15_LC_12_17_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i15_LC_12_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i15_LC_12_17_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i15_LC_12_17_1  (
            .in0(N__30279),
            .in1(N__36960),
            .in2(_gnd_net_),
            .in3(N__43260),
            .lcout(data_in_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66754),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i16_LC_12_17_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i16_LC_12_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i16_LC_12_17_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i16_LC_12_17_2  (
            .in0(N__43258),
            .in1(N__36625),
            .in2(_gnd_net_),
            .in3(N__30498),
            .lcout(data_in_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66754),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__7__5430_LC_12_17_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__7__5430_LC_12_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__7__5430_LC_12_17_3 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_out_frame_11__7__5430_LC_12_17_3  (
            .in0(N__48933),
            .in1(N__32893),
            .in2(N__49451),
            .in3(N__28704),
            .lcout(data_out_frame_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66754),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i20_LC_12_17_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i20_LC_12_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i20_LC_12_17_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i20_LC_12_17_4  (
            .in0(N__43259),
            .in1(N__34192),
            .in2(_gnd_net_),
            .in3(N__29074),
            .lcout(data_in_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66754),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1771_LC_12_17_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1771_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1771_LC_12_17_5 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i6_4_lut_adj_1771_LC_12_17_5  (
            .in0(N__30557),
            .in1(N__28888),
            .in2(N__41960),
            .in3(N__41994),
            .lcout(\c0.n15_adj_4496 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i6_LC_12_17_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i6_LC_12_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i6_LC_12_17_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i6_LC_12_17_6  (
            .in0(N__28889),
            .in1(N__43261),
            .in2(_gnd_net_),
            .in3(N__30300),
            .lcout(data_in_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66754),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__3__5426_LC_12_17_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__3__5426_LC_12_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__3__5426_LC_12_17_7 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_out_frame_12__3__5426_LC_12_17_7  (
            .in0(N__48934),
            .in1(N__32979),
            .in2(N__49452),
            .in3(N__28912),
            .lcout(data_out_frame_12_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66754),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1756_LC_12_18_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1756_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1756_LC_12_18_0 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i1_4_lut_adj_1756_LC_12_18_0  (
            .in0(N__41998),
            .in1(N__28844),
            .in2(N__30256),
            .in3(N__28864),
            .lcout(),
            .ltout(\c0.n7_adj_4492_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1761_LC_12_18_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1761_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1761_LC_12_18_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i5_4_lut_adj_1761_LC_12_18_1  (
            .in0(N__40242),
            .in1(N__28857),
            .in2(N__28900),
            .in3(N__28870),
            .lcout(\c0.n63_adj_4301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_LC_12_18_3 .C_ON=1'b0;
    defparam \c0.i3_2_lut_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_LC_12_18_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i3_2_lut_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__28896),
            .in2(_gnd_net_),
            .in3(N__30366),
            .lcout(\c0.n9_adj_4493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i7_LC_12_18_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i7_LC_12_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i7_LC_12_18_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i7_LC_12_18_4  (
            .in0(N__28858),
            .in1(N__30283),
            .in2(_gnd_net_),
            .in3(N__43262),
            .lcout(data_in_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66768),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1706_LC_12_18_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1706_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1706_LC_12_18_5 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i3_4_lut_adj_1706_LC_12_18_5  (
            .in0(N__30550),
            .in1(N__41967),
            .in2(N__28822),
            .in3(N__30591),
            .lcout(\c0.n23600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1769_LC_12_18_6 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1769_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1769_LC_12_18_6 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.i5_3_lut_adj_1769_LC_12_18_6  (
            .in0(N__28856),
            .in1(N__40241),
            .in2(_gnd_net_),
            .in3(N__30252),
            .lcout(),
            .ltout(\c0.n14_adj_4495_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1772_LC_12_18_7 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1772_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1772_LC_12_18_7 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i8_4_lut_adj_1772_LC_12_18_7  (
            .in0(N__28843),
            .in1(N__28818),
            .in2(N__28795),
            .in3(N__28792),
            .lcout(\c0.n21767 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1773_LC_12_19_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1773_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1773_LC_12_19_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i2_2_lut_adj_1773_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(N__35253),
            .in2(_gnd_net_),
            .in3(N__34193),
            .lcout(),
            .ltout(\c0.n10_adj_4231_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1241_LC_12_19_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1241_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1241_LC_12_19_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i7_4_lut_adj_1241_LC_12_19_1  (
            .in0(N__34165),
            .in1(N__36993),
            .in2(N__29164),
            .in3(N__29161),
            .lcout(\c0.n13003 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_3_lut_4_lut_LC_12_19_3 .C_ON=1'b0;
    defparam \c0.tx.i2_3_lut_4_lut_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_3_lut_4_lut_LC_12_19_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \c0.tx.i2_3_lut_4_lut_LC_12_19_3  (
            .in0(N__41445),
            .in1(N__39268),
            .in2(N__33771),
            .in3(N__30711),
            .lcout(n9539),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__0__5445_LC_12_19_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__0__5445_LC_12_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__0__5445_LC_12_19_4 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_10__0__5445_LC_12_19_4  (
            .in0(N__49512),
            .in1(N__48944),
            .in2(N__29962),
            .in3(N__29088),
            .lcout(data_out_frame_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66782),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i28_LC_12_19_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i28_LC_12_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i28_LC_12_19_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i28_LC_12_19_5  (
            .in0(N__64872),
            .in1(N__43267),
            .in2(_gnd_net_),
            .in3(N__29070),
            .lcout(data_in_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66782),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i9_LC_12_19_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i9_LC_12_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i9_LC_12_19_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_in_0___i9_LC_12_19_6  (
            .in0(N__43266),
            .in1(_gnd_net_),
            .in2(N__30558),
            .in3(N__36220),
            .lcout(data_in_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66782),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__2__5435_LC_12_19_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__2__5435_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__2__5435_LC_12_19_7 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_11__2__5435_LC_12_19_7  (
            .in0(N__48943),
            .in1(N__49513),
            .in2(N__29050),
            .in3(N__29010),
            .lcout(data_out_frame_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66782),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20481_LC_12_20_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20481_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_20481_LC_12_20_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_20481_LC_12_20_0  (
            .in0(N__30133),
            .in1(N__36883),
            .in2(N__29011),
            .in3(N__39804),
            .lcout(\c0.n24177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__0__5485_LC_12_20_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__0__5485_LC_12_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__0__5485_LC_12_20_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_5__0__5485_LC_12_20_1  (
            .in0(N__49476),
            .in1(N__48896),
            .in2(N__44623),
            .in3(N__28983),
            .lcout(data_out_frame_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66794),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__5__5440_LC_12_20_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__5__5440_LC_12_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__5__5440_LC_12_20_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.data_out_frame_10__5__5440_LC_12_20_3  (
            .in0(N__49475),
            .in1(N__28966),
            .in2(N__28930),
            .in3(N__48897),
            .lcout(data_out_frame_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66794),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_1181_LC_12_20_4 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_1181_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_1181_LC_12_20_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.tx.i1_2_lut_adj_1181_LC_12_20_4  (
            .in0(N__33768),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30643),
            .lcout(),
            .ltout(\c0.tx.n16631_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_4_lut_adj_1187_LC_12_20_5 .C_ON=1'b0;
    defparam \c0.tx.i2_4_lut_adj_1187_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_4_lut_adj_1187_LC_12_20_5 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \c0.tx.i2_4_lut_adj_1187_LC_12_20_5  (
            .in0(N__30707),
            .in1(N__41443),
            .in2(N__29203),
            .in3(N__33706),
            .lcout(\c0.tx.n14296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_4_lut_LC_12_20_6 .C_ON=1'b0;
    defparam \c0.tx.i2_4_lut_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_4_lut_LC_12_20_6 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \c0.tx.i2_4_lut_LC_12_20_6  (
            .in0(N__33767),
            .in1(N__30706),
            .in2(N__41467),
            .in3(N__30642),
            .lcout(n14442),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i2_LC_12_20_7 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i2_LC_12_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i2_LC_12_20_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.tx.r_SM_Main_i2_LC_12_20_7  (
            .in0(N__30644),
            .in1(N__33769),
            .in2(N__30721),
            .in3(N__41444),
            .lcout(r_SM_Main_2_adj_4549),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66794),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i3_LC_12_21_0 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i3_LC_12_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i3_LC_12_21_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i3_LC_12_21_0  (
            .in0(N__30844),
            .in1(N__41456),
            .in2(_gnd_net_),
            .in3(N__30826),
            .lcout(\c0.tx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66804),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1770_LC_12_21_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1770_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1770_LC_12_21_2 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1770_LC_12_21_2  (
            .in0(N__34301),
            .in1(N__52981),
            .in2(_gnd_net_),
            .in3(N__53194),
            .lcout(\c0.n21370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1597_LC_12_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1597_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1597_LC_12_21_4 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i1_2_lut_adj_1597_LC_12_21_4  (
            .in0(_gnd_net_),
            .in1(N__46176),
            .in2(_gnd_net_),
            .in3(N__42985),
            .lcout(\c0.n38_adj_4390 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i1_LC_12_21_6 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i1_LC_12_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i1_LC_12_21_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i1_LC_12_21_6  (
            .in0(N__30898),
            .in1(N__41455),
            .in2(_gnd_net_),
            .in3(N__30880),
            .lcout(\c0.tx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66804),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i2_LC_12_21_7 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i2_LC_12_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i2_LC_12_21_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i2_LC_12_21_7  (
            .in0(N__41454),
            .in1(N__30871),
            .in2(_gnd_net_),
            .in3(N__30853),
            .lcout(\c0.tx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66804),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1776_LC_12_22_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1776_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1776_LC_12_22_0 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1776_LC_12_22_0  (
            .in0(N__37334),
            .in1(N__53181),
            .in2(_gnd_net_),
            .in3(N__53011),
            .lcout(\c0.n21376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1598_LC_12_22_7 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1598_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1598_LC_12_22_7 .LUT_INIT=16'b1111111100110001;
    LogicCell40 \c0.i1_4_lut_adj_1598_LC_12_22_7  (
            .in0(N__31009),
            .in1(N__42834),
            .in2(N__46177),
            .in3(N__40471),
            .lcout(\c0.n4_adj_4391 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i8_LC_12_23_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i8_LC_12_23_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i8_LC_12_23_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i8_LC_12_23_0  (
            .in0(_gnd_net_),
            .in1(N__34246),
            .in2(_gnd_net_),
            .in3(N__52870),
            .lcout(\c0.FRAME_MATCHER_state_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66826),
            .ce(),
            .sr(N__34222));
    defparam \c0.FRAME_MATCHER_state_i17_LC_12_24_2 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i17_LC_12_24_2 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i17_LC_12_24_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i17_LC_12_24_2  (
            .in0(_gnd_net_),
            .in1(N__37847),
            .in2(_gnd_net_),
            .in3(N__52873),
            .lcout(\c0.FRAME_MATCHER_state_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66838),
            .ce(),
            .sr(N__29233));
    defparam \c0.FRAME_MATCHER_state_i18_LC_12_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i18_LC_12_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i18_LC_12_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i18_LC_12_25_0  (
            .in0(_gnd_net_),
            .in1(N__37903),
            .in2(_gnd_net_),
            .in3(N__52874),
            .lcout(\c0.FRAME_MATCHER_state_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66849),
            .ce(),
            .sr(N__37570));
    defparam \c0.i1_2_lut_3_lut_adj_1762_LC_12_26_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1762_LC_12_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1762_LC_12_26_7 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1762_LC_12_26_7  (
            .in0(N__37876),
            .in1(N__53175),
            .in2(_gnd_net_),
            .in3(N__53027),
            .lcout(\c0.n21360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1759_LC_12_27_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1759_LC_12_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1759_LC_12_27_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1759_LC_12_27_4  (
            .in0(N__34564),
            .in1(N__53197),
            .in2(_gnd_net_),
            .in3(N__53028),
            .lcout(\c0.n21356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1846_LC_13_6_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1846_LC_13_6_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1846_LC_13_6_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1846_LC_13_6_0  (
            .in0(N__31993),
            .in1(N__31434),
            .in2(N__29227),
            .in3(N__31570),
            .lcout(\c0.n12_adj_4516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1874_LC_13_7_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1874_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1874_LC_13_7_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1874_LC_13_7_0  (
            .in0(N__34454),
            .in1(N__29578),
            .in2(_gnd_net_),
            .in3(N__31070),
            .lcout(\c0.n9_adj_4339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1885_LC_13_7_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1885_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1885_LC_13_7_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1885_LC_13_7_3  (
            .in0(N__31404),
            .in1(N__29411),
            .in2(_gnd_net_),
            .in3(N__34452),
            .lcout(\c0.n22018 ),
            .ltout(\c0.n22018_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1398_LC_13_7_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1398_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1398_LC_13_7_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1398_LC_13_7_4  (
            .in0(N__32204),
            .in1(N__29577),
            .in2(N__29380),
            .in3(N__30967),
            .lcout(\c0.n21946 ),
            .ltout(\c0.n21946_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1627_LC_13_7_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1627_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1627_LC_13_7_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1627_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__29358),
            .in2(N__29362),
            .in3(N__29412),
            .lcout(\c0.n6_adj_4402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_3_lut_4_lut_LC_13_7_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_3_lut_4_lut_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_3_lut_4_lut_LC_13_7_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_3_lut_4_lut_LC_13_7_7  (
            .in0(N__31688),
            .in1(N__34453),
            .in2(N__31351),
            .in3(N__31295),
            .lcout(\c0.n22188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1599_LC_13_8_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1599_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1599_LC_13_8_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1599_LC_13_8_0  (
            .in0(N__31634),
            .in1(N__31341),
            .in2(N__31418),
            .in3(N__31297),
            .lcout(),
            .ltout(\c0.n12491_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__6__5295_LC_13_8_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__6__5295_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__6__5295_LC_13_8_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_28__6__5295_LC_13_8_1  (
            .in0(N__29466),
            .in1(N__29359),
            .in2(N__29320),
            .in3(N__34362),
            .lcout(\c0.data_out_frame_28_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66644),
            .ce(N__40950),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i26_3_lut_LC_13_8_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i26_3_lut_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i26_3_lut_LC_13_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_6_i26_3_lut_LC_13_8_2  (
            .in0(N__31777),
            .in1(N__29317),
            .in2(_gnd_net_),
            .in3(N__39836),
            .lcout(\c0.n26_adj_4351 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1608_LC_13_8_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1608_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1608_LC_13_8_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_adj_1608_LC_13_8_3  (
            .in0(N__31296),
            .in1(N__31337),
            .in2(N__31219),
            .in3(N__31633),
            .lcout(),
            .ltout(\c0.n7_adj_4307_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1401_LC_13_8_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1401_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1401_LC_13_8_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1401_LC_13_8_4  (
            .in0(N__31088),
            .in1(N__29271),
            .in2(N__29296),
            .in3(N__29529),
            .lcout(data_out_frame_29__3__N_1662),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__4__5289_LC_13_8_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__4__5289_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__4__5289_LC_13_8_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_29__4__5289_LC_13_8_5  (
            .in0(N__29530),
            .in1(N__29491),
            .in2(N__31102),
            .in3(N__29272),
            .lcout(\c0.data_out_frame_29_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66644),
            .ce(N__40950),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1832_LC_13_8_6 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1832_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1832_LC_13_8_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_3_lut_adj_1832_LC_13_8_6  (
            .in0(N__31405),
            .in1(N__31217),
            .in2(_gnd_net_),
            .in3(N__31071),
            .lcout(\c0.n22151 ),
            .ltout(\c0.n22151_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__5__5288_LC_13_8_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__5__5288_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__5__5288_LC_13_8_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.data_out_frame_29__5__5288_LC_13_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29485),
            .in3(N__29742),
            .lcout(\c0.data_out_frame_29_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66644),
            .ce(N__40950),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1618_LC_13_9_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1618_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1618_LC_13_9_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1618_LC_13_9_0  (
            .in0(N__32380),
            .in1(N__31988),
            .in2(_gnd_net_),
            .in3(N__32932),
            .lcout(),
            .ltout(\c0.n6_adj_4397_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__0__5301_LC_13_9_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__0__5301_LC_13_9_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__0__5301_LC_13_9_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame_28__0__5301_LC_13_9_1  (
            .in0(N__29728),
            .in1(N__32114),
            .in2(N__29482),
            .in3(N__29806),
            .lcout(\c0.data_out_frame_28_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66651),
            .ce(N__40954),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1825_LC_13_9_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1825_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1825_LC_13_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1825_LC_13_9_2  (
            .in0(N__32113),
            .in1(N__32245),
            .in2(N__31838),
            .in3(N__29727),
            .lcout(\c0.n21876 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__5__5296_LC_13_9_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__5__5296_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__5__5296_LC_13_9_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.data_out_frame_28__5__5296_LC_13_9_4  (
            .in0(N__32211),
            .in1(_gnd_net_),
            .in2(N__29473),
            .in3(N__31462),
            .lcout(\c0.data_out_frame_28_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66651),
            .ce(N__40954),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i26_3_lut_LC_13_9_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i26_3_lut_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i26_3_lut_LC_13_9_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_5_i26_3_lut_LC_13_9_5  (
            .in0(N__39837),
            .in1(N__29455),
            .in2(_gnd_net_),
            .in3(N__29449),
            .lcout(\c0.n26_adj_4347 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1714_LC_13_10_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1714_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1714_LC_13_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1714_LC_13_10_0  (
            .in0(N__29853),
            .in1(N__31208),
            .in2(_gnd_net_),
            .in3(N__29766),
            .lcout(\c0.n21210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1819_LC_13_10_1 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1819_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1819_LC_13_10_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_3_lut_adj_1819_LC_13_10_1  (
            .in0(N__31656),
            .in1(N__29424),
            .in2(_gnd_net_),
            .in3(N__32248),
            .lcout(),
            .ltout(\c0.n6_adj_4509_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1820_LC_13_10_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1820_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1820_LC_13_10_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1820_LC_13_10_2  (
            .in0(N__34928),
            .in1(N__29575),
            .in2(N__29611),
            .in3(N__34817),
            .lcout(\c0.n22393 ),
            .ltout(\c0.n22393_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1822_LC_13_10_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1822_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1822_LC_13_10_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1822_LC_13_10_3  (
            .in0(N__29601),
            .in1(N__31218),
            .in2(N__29584),
            .in3(N__32014),
            .lcout(),
            .ltout(\c0.n14_adj_4510_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1823_LC_13_10_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1823_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1823_LC_13_10_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1823_LC_13_10_4  (
            .in0(N__38295),
            .in1(N__31922),
            .in2(N__29581),
            .in3(N__29509),
            .lcout(\c0.n22346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1875_LC_13_10_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1875_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1875_LC_13_10_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1875_LC_13_10_5  (
            .in0(N__29576),
            .in1(N__34445),
            .in2(_gnd_net_),
            .in3(N__29520),
            .lcout(\c0.n10_adj_4511 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1818_LC_13_10_7 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1818_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1818_LC_13_10_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_3_lut_adj_1818_LC_13_10_7  (
            .in0(N__32733),
            .in1(N__53392),
            .in2(_gnd_net_),
            .in3(N__29824),
            .lcout(\c0.n22177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1865_LC_13_11_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1865_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1865_LC_13_11_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1865_LC_13_11_0  (
            .in0(N__29851),
            .in1(N__38966),
            .in2(N__32738),
            .in3(N__29780),
            .lcout(\c0.n20274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1424_LC_13_11_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1424_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1424_LC_13_11_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_1424_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__29850),
            .in2(_gnd_net_),
            .in3(N__29764),
            .lcout(\c0.n21192 ),
            .ltout(\c0.n21192_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1463_LC_13_11_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1463_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1463_LC_13_11_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_1463_LC_13_11_2  (
            .in0(N__30082),
            .in1(N__29503),
            .in2(N__29497),
            .in3(N__38590),
            .lcout(\c0.n20931 ),
            .ltout(\c0.n20931_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1867_LC_13_11_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1867_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1867_LC_13_11_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1867_LC_13_11_3  (
            .in0(N__38967),
            .in1(N__32726),
            .in2(N__29494),
            .in3(N__29825),
            .lcout(\c0.n21283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1421_LC_13_11_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1421_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1421_LC_13_11_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_1421_LC_13_11_4  (
            .in0(N__29852),
            .in1(_gnd_net_),
            .in2(N__29830),
            .in3(_gnd_net_),
            .lcout(\c0.n12554 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1868_LC_13_11_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1868_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1868_LC_13_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1868_LC_13_11_5  (
            .in0(N__29781),
            .in1(N__32725),
            .in2(N__38971),
            .in3(N__29765),
            .lcout(\c0.n21189 ),
            .ltout(\c0.n21189_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1802_LC_13_11_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1802_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1802_LC_13_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1802_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__31377),
            .in2(N__29746),
            .in3(N__29743),
            .lcout(\c0.n20151 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1878_LC_13_11_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1878_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1878_LC_13_11_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1878_LC_13_11_7  (
            .in0(N__35213),
            .in1(N__32824),
            .in2(N__32302),
            .in3(N__29721),
            .lcout(\c0.n10513 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1697_LC_13_12_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1697_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1697_LC_13_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1697_LC_13_12_0  (
            .in0(N__38294),
            .in1(N__35116),
            .in2(N__32739),
            .in3(N__29706),
            .lcout(\c0.n10467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1742_LC_13_12_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1742_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1742_LC_13_12_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1742_LC_13_12_1  (
            .in0(N__29659),
            .in1(_gnd_net_),
            .in2(N__36460),
            .in3(N__35316),
            .lcout(\c0.n13480 ),
            .ltout(\c0.n13480_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1737_LC_13_12_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1737_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1737_LC_13_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1737_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__31877),
            .in2(N__29671),
            .in3(N__31956),
            .lcout(\c0.n21122 ),
            .ltout(\c0.n21122_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1589_LC_13_12_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1589_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1589_LC_13_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1589_LC_13_12_3  (
            .in0(N__32367),
            .in1(N__31882),
            .in2(N__29668),
            .in3(N__32420),
            .lcout(\c0.data_out_frame_29__7__N_1144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20421_2_lut_3_lut_4_lut_LC_13_12_4 .C_ON=1'b0;
    defparam \c0.i20421_2_lut_3_lut_4_lut_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i20421_2_lut_3_lut_4_lut_LC_13_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20421_2_lut_3_lut_4_lut_LC_13_12_4  (
            .in0(N__31881),
            .in1(N__36458),
            .in2(N__35320),
            .in3(N__29660),
            .lcout(\c0.n24119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1426_LC_13_12_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1426_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1426_LC_13_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1426_LC_13_12_5  (
            .in0(N__30164),
            .in1(N__39292),
            .in2(_gnd_net_),
            .in3(N__39430),
            .lcout(\c0.n20767 ),
            .ltout(\c0.n20767_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1427_LC_13_12_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1427_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1427_LC_13_12_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1427_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29965),
            .in3(N__34627),
            .lcout(\c0.n21848 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1882_LC_13_12_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1882_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1882_LC_13_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1882_LC_13_12_7  (
            .in0(N__31957),
            .in1(N__32493),
            .in2(_gnd_net_),
            .in3(N__32421),
            .lcout(\c0.n21112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1409_LC_13_13_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1409_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1409_LC_13_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1409_LC_13_13_0  (
            .in0(N__36165),
            .in1(N__33244),
            .in2(N__29957),
            .in3(N__38563),
            .lcout(\c0.n21943 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i10_LC_13_13_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i10_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i10_LC_13_13_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i10_LC_13_13_2  (
            .in0(N__29914),
            .in1(N__38459),
            .in2(_gnd_net_),
            .in3(N__35209),
            .lcout(encoder1_position_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66686),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__6__5447_LC_13_13_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__6__5447_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__6__5447_LC_13_13_3 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_9__6__5447_LC_13_13_3  (
            .in0(N__49332),
            .in1(N__49026),
            .in2(N__29902),
            .in3(N__36166),
            .lcout(data_out_frame_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66686),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__6__5415_LC_13_13_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__6__5415_LC_13_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__6__5415_LC_13_13_4 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_13__6__5415_LC_13_13_4  (
            .in0(N__49024),
            .in1(N__49333),
            .in2(N__34984),
            .in3(N__29883),
            .lcout(data_out_frame_13_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66686),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__4__5457_LC_13_13_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__4__5457_LC_13_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__4__5457_LC_13_13_5 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_8__4__5457_LC_13_13_5  (
            .in0(N__49331),
            .in1(N__49025),
            .in2(N__30232),
            .in3(N__38874),
            .lcout(data_out_frame_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66686),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i11_LC_13_13_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i11_LC_13_13_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i11_LC_13_13_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i11_LC_13_13_6  (
            .in0(N__29866),
            .in1(N__38460),
            .in2(_gnd_net_),
            .in3(N__32965),
            .lcout(encoder1_position_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66686),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_13_13_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_13_13_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_13_13_7  (
            .in0(N__39818),
            .in1(N__35002),
            .in2(_gnd_net_),
            .in3(N__35170),
            .lcout(\c0.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1462_LC_13_14_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1462_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1462_LC_13_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1462_LC_13_14_0  (
            .in0(N__53388),
            .in1(N__35284),
            .in2(N__41605),
            .in3(N__39060),
            .lcout(\c0.n14_adj_4329 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i7_LC_13_14_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i7_LC_13_14_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i7_LC_13_14_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter1.count_i0_i7_LC_13_14_1  (
            .in0(N__34907),
            .in1(N__30073),
            .in2(_gnd_net_),
            .in3(N__38465),
            .lcout(encoder1_position_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66700),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i13_LC_13_14_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i13_LC_13_14_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i13_LC_13_14_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i13_LC_13_14_2  (
            .in0(N__38461),
            .in1(N__30061),
            .in2(_gnd_net_),
            .in3(N__38046),
            .lcout(encoder1_position_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66700),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1690_LC_13_14_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1690_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1690_LC_13_14_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1690_LC_13_14_3  (
            .in0(N__38247),
            .in1(N__35762),
            .in2(N__30030),
            .in3(N__48533),
            .lcout(\c0.n21855 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i19_LC_13_14_4 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i19_LC_13_14_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i19_LC_13_14_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \quad_counter1.count_i0_i19_LC_13_14_4  (
            .in0(N__30049),
            .in1(_gnd_net_),
            .in2(N__38496),
            .in3(N__30025),
            .lcout(encoder1_position_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66700),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_LC_13_14_5 .C_ON=1'b0;
    defparam \c0.i11_3_lut_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_LC_13_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i11_3_lut_LC_13_14_5  (
            .in0(N__30004),
            .in1(N__35668),
            .in2(_gnd_net_),
            .in3(N__30238),
            .lcout(\c0.n23557 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i2_LC_13_14_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i2_LC_13_14_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i2_LC_13_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i2_LC_13_14_6  (
            .in0(N__42222),
            .in1(N__33112),
            .in2(_gnd_net_),
            .in3(N__53448),
            .lcout(encoder0_position_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66700),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i30_LC_13_14_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i30_LC_13_14_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i30_LC_13_14_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i30_LC_13_14_7  (
            .in0(N__48553),
            .in1(N__33325),
            .in2(_gnd_net_),
            .in3(N__42223),
            .lcout(encoder0_position_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66700),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i25_LC_13_15_0 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i25_LC_13_15_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i25_LC_13_15_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i25_LC_13_15_0  (
            .in0(N__38466),
            .in1(N__29992),
            .in2(_gnd_net_),
            .in3(N__33010),
            .lcout(encoder1_position_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66714),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i7_LC_13_15_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i7_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i7_LC_13_15_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \quad_counter0.count_i0_i7_LC_13_15_1  (
            .in0(N__33199),
            .in1(_gnd_net_),
            .in2(N__42231),
            .in3(N__33249),
            .lcout(encoder0_position_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66714),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1441_LC_13_15_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1441_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1441_LC_13_15_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1441_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(N__33230),
            .in2(_gnd_net_),
            .in3(N__41811),
            .lcout(),
            .ltout(\c0.n21914_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1446_LC_13_15_3 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1446_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1446_LC_13_15_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1446_LC_13_15_3  (
            .in0(N__53436),
            .in1(N__38167),
            .in2(N__30241),
            .in3(N__37061),
            .lcout(\c0.n21_adj_4320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i19_LC_13_15_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i19_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i19_LC_13_15_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i19_LC_13_15_5  (
            .in0(N__42180),
            .in1(N__33286),
            .in2(_gnd_net_),
            .in3(N__38652),
            .lcout(encoder0_position_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66714),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20185_3_lut_LC_13_15_6 .C_ON=1'b0;
    defparam \c0.i20185_3_lut_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i20185_3_lut_LC_13_15_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i20185_3_lut_LC_13_15_6  (
            .in0(N__39817),
            .in1(N__30192),
            .in2(_gnd_net_),
            .in3(N__30231),
            .lcout(\c0.n23880 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__4__5449_LC_13_15_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__4__5449_LC_13_15_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__4__5449_LC_13_15_7 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \c0.data_out_frame_9__4__5449_LC_13_15_7  (
            .in0(N__39040),
            .in1(N__48946),
            .in2(N__30196),
            .in3(N__49402),
            .lcout(data_out_frame_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66714),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i27_LC_13_16_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i27_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i27_LC_13_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i27_LC_13_16_1  (
            .in0(N__38506),
            .in1(N__30184),
            .in2(_gnd_net_),
            .in3(N__30163),
            .lcout(encoder1_position_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66728),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__2__5443_LC_13_16_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__2__5443_LC_13_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__2__5443_LC_13_16_2 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_10__2__5443_LC_13_16_2  (
            .in0(N__49472),
            .in1(N__48887),
            .in2(N__35659),
            .in3(N__30129),
            .lcout(data_out_frame_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66728),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__4__5481_LC_13_16_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__4__5481_LC_13_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__4__5481_LC_13_16_3 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_5__4__5481_LC_13_16_3  (
            .in0(N__48886),
            .in1(N__49474),
            .in2(N__42403),
            .in3(N__30111),
            .lcout(data_out_frame_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66728),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__4__5473_LC_13_16_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__4__5473_LC_13_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__4__5473_LC_13_16_4 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_frame_6__4__5473_LC_13_16_4  (
            .in0(N__49473),
            .in1(N__30384),
            .in2(N__38785),
            .in3(N__48888),
            .lcout(data_out_frame_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66728),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20139_4_lut_LC_13_16_5 .C_ON=1'b0;
    defparam \c0.i20139_4_lut_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20139_4_lut_LC_13_16_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i20139_4_lut_LC_13_16_5  (
            .in0(N__30340),
            .in1(N__36381),
            .in2(N__36310),
            .in3(N__36594),
            .lcout(\c0.n23834 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1691_LC_13_16_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1691_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1691_LC_13_16_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1691_LC_13_16_7  (
            .in0(N__35997),
            .in1(N__36122),
            .in2(N__33243),
            .in3(N__41810),
            .lcout(\c0.n22449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i4_LC_13_17_0 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i4_LC_13_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i4_LC_13_17_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i4_LC_13_17_0  (
            .in0(N__30809),
            .in1(N__41486),
            .in2(_gnd_net_),
            .in3(N__30793),
            .lcout(\c0.tx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66741),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1536_LC_13_17_2 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1536_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1536_LC_13_17_2 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \c0.i8_4_lut_adj_1536_LC_13_17_2  (
            .in0(N__30370),
            .in1(N__30299),
            .in2(N__36216),
            .in3(N__36646),
            .lcout(),
            .ltout(\c0.n20_adj_4362_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_adj_1596_LC_13_17_3 .C_ON=1'b0;
    defparam \c0.i11_3_lut_adj_1596_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_adj_1596_LC_13_17_3 .LUT_INIT=16'b1111110011111111;
    LogicCell40 \c0.i11_3_lut_adj_1596_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__30355),
            .in2(N__30349),
            .in3(N__30346),
            .lcout(\c0.n63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1702_LC_13_17_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1702_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1702_LC_13_17_5 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i7_4_lut_adj_1702_LC_13_17_5  (
            .in0(N__36948),
            .in1(N__30339),
            .in2(N__30301),
            .in3(N__36587),
            .lcout(),
            .ltout(\c0.n17_adj_4479_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1703_LC_13_17_6 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1703_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1703_LC_13_17_6 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i9_4_lut_adj_1703_LC_13_17_6  (
            .in0(N__30277),
            .in1(N__36645),
            .in2(N__30259),
            .in3(N__36343),
            .lcout(\c0.n13006 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1765_LC_13_18_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1765_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1765_LC_13_18_0 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \c0.i5_3_lut_adj_1765_LC_13_18_0  (
            .in0(N__41893),
            .in1(N__36624),
            .in2(_gnd_net_),
            .in3(N__30478),
            .lcout(\c0.n13023 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i5_LC_13_18_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i5_LC_13_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i5_LC_13_18_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i5_LC_13_18_1  (
            .in0(N__30513),
            .in1(N__43269),
            .in2(_gnd_net_),
            .in3(N__41968),
            .lcout(data_in_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66755),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1695_LC_13_18_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1695_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1695_LC_13_18_2 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \c0.i7_4_lut_adj_1695_LC_13_18_2  (
            .in0(N__30619),
            .in1(N__30592),
            .in2(N__35260),
            .in3(N__30579),
            .lcout(\c0.n17_adj_4477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_47_LC_13_18_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_47_LC_13_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Active_47_LC_13_18_3 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \c0.tx.r_Tx_Active_47_LC_13_18_3  (
            .in0(N__30568),
            .in1(N__37142),
            .in2(_gnd_net_),
            .in3(N__30720),
            .lcout(\c0.tx_active ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66755),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i10_LC_13_18_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i10_LC_13_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i10_LC_13_18_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i10_LC_13_18_4  (
            .in0(N__34164),
            .in1(_gnd_net_),
            .in2(N__43273),
            .in3(N__36324),
            .lcout(data_in_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66755),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i1_LC_13_18_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i1_LC_13_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i1_LC_13_18_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_in_0___i1_LC_13_18_5  (
            .in0(N__30526),
            .in1(_gnd_net_),
            .in2(N__30559),
            .in3(N__43268),
            .lcout(data_in_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66755),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1763_LC_13_18_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1763_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1763_LC_13_18_7 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.i4_4_lut_adj_1763_LC_13_18_7  (
            .in0(N__36323),
            .in1(N__30525),
            .in2(N__30514),
            .in3(N__30494),
            .lcout(\c0.n10_adj_4494 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1699_LC_13_19_0 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1699_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1699_LC_13_19_0 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i9_4_lut_adj_1699_LC_13_19_0  (
            .in0(N__34156),
            .in1(N__34197),
            .in2(N__30472),
            .in3(N__30460),
            .lcout(\c0.n117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1744_LC_13_19_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1744_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1744_LC_13_19_1 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1744_LC_13_19_1  (
            .in0(N__39264),
            .in1(N__37135),
            .in2(_gnd_net_),
            .in3(N__37171),
            .lcout(\c0.n44_adj_4336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1448020_i1_3_lut_LC_13_19_2.C_ON=1'b0;
    defparam i1448020_i1_3_lut_LC_13_19_2.SEQ_MODE=4'b0000;
    defparam i1448020_i1_3_lut_LC_13_19_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 i1448020_i1_3_lut_LC_13_19_2 (
            .in0(N__30454),
            .in1(N__30409),
            .in2(_gnd_net_),
            .in3(N__30400),
            .lcout(),
            .ltout(o_Tx_Serial_N_3783_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i26_3_lut_LC_13_19_3 .C_ON=1'b0;
    defparam \c0.tx.i26_3_lut_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i26_3_lut_LC_13_19_3 .LUT_INIT=16'b0101010100001010;
    LogicCell40 \c0.tx.i26_3_lut_LC_13_19_3  (
            .in0(N__30704),
            .in1(_gnd_net_),
            .in2(N__30751),
            .in3(N__33763),
            .lcout(\c0.tx.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i1_LC_13_19_4 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i1_LC_13_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i1_LC_13_19_4 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \c0.tx.r_SM_Main_i1_LC_13_19_4  (
            .in0(N__30650),
            .in1(N__30705),
            .in2(N__33772),
            .in3(N__41490),
            .lcout(r_SM_Main_1_adj_4550),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66769),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_1184_LC_13_19_6 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_1184_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_1184_LC_13_19_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.i1_2_lut_adj_1184_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(N__33756),
            .in2(_gnd_net_),
            .in3(N__30703),
            .lcout(\c0.tx.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i7_LC_13_19_7 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i7_LC_13_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i7_LC_13_19_7 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.tx.r_Clock_Count__i7_LC_13_19_7  (
            .in0(N__31024),
            .in1(N__31047),
            .in2(N__41496),
            .in3(N__41382),
            .lcout(r_Clock_Count_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66769),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_LC_13_20_0 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_LC_13_20_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.i1_2_lut_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__41547),
            .in2(_gnd_net_),
            .in3(N__30778),
            .lcout(),
            .ltout(\c0.tx.n6_adj_4214_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4_4_lut_adj_1180_LC_13_20_1 .C_ON=1'b0;
    defparam \c0.tx.i4_4_lut_adj_1180_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4_4_lut_adj_1180_LC_13_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx.i4_4_lut_adj_1180_LC_13_20_1  (
            .in0(N__41342),
            .in1(N__31043),
            .in2(N__30664),
            .in3(N__30958),
            .lcout(\c0.tx.n16630 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_LC_13_20_2 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_LC_13_20_2 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \c0.tx.i1_4_lut_LC_13_20_2  (
            .in0(N__41457),
            .in1(N__41343),
            .in2(N__30943),
            .in3(N__41548),
            .lcout(n8),
            .ltout(n8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i5_LC_13_20_3 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i5_LC_13_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i5_LC_13_20_3 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \c0.tx.r_Clock_Count__i5_LC_13_20_3  (
            .in0(N__30760),
            .in1(N__30781),
            .in2(N__30622),
            .in3(N__41458),
            .lcout(r_Clock_Count_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66783),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_1186_LC_13_20_4 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_1186_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_1186_LC_13_20_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx.i1_2_lut_adj_1186_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(N__30816),
            .in2(_gnd_net_),
            .in3(N__30842),
            .lcout(),
            .ltout(\c0.tx.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4_4_lut_LC_13_20_5 .C_ON=1'b0;
    defparam \c0.tx.i4_4_lut_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4_4_lut_LC_13_20_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx.i4_4_lut_LC_13_20_5  (
            .in0(N__30934),
            .in1(N__30896),
            .in2(N__30961),
            .in3(N__30869),
            .lcout(\c0.tx.n31 ),
            .ltout(\c0.tx.n31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4_4_lut_adj_1185_LC_13_20_6 .C_ON=1'b0;
    defparam \c0.tx.i4_4_lut_adj_1185_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4_4_lut_adj_1185_LC_13_20_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \c0.tx.i4_4_lut_adj_1185_LC_13_20_6  (
            .in0(N__31042),
            .in1(N__30779),
            .in2(N__30952),
            .in3(N__30949),
            .lcout(\c0.tx.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_2_lut_LC_13_21_0 .C_ON=1'b1;
    defparam \c0.tx.add_59_2_lut_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_2_lut_LC_13_21_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_2_lut_LC_13_21_0  (
            .in0(N__41374),
            .in1(N__30933),
            .in2(_gnd_net_),
            .in3(N__30901),
            .lcout(\c0.tx.n23960 ),
            .ltout(),
            .carryin(bfn_13_21_0_),
            .carryout(\c0.tx.n19540 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_3_lut_LC_13_21_1 .C_ON=1'b1;
    defparam \c0.tx.add_59_3_lut_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_3_lut_LC_13_21_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_3_lut_LC_13_21_1  (
            .in0(N__41377),
            .in1(N__30897),
            .in2(_gnd_net_),
            .in3(N__30874),
            .lcout(\c0.tx.n23961 ),
            .ltout(),
            .carryin(\c0.tx.n19540 ),
            .carryout(\c0.tx.n19541 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_4_lut_LC_13_21_2 .C_ON=1'b1;
    defparam \c0.tx.add_59_4_lut_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_4_lut_LC_13_21_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_4_lut_LC_13_21_2  (
            .in0(N__41376),
            .in1(N__30870),
            .in2(_gnd_net_),
            .in3(N__30847),
            .lcout(\c0.tx.n23958 ),
            .ltout(),
            .carryin(\c0.tx.n19541 ),
            .carryout(\c0.tx.n19542 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_5_lut_LC_13_21_3 .C_ON=1'b1;
    defparam \c0.tx.add_59_5_lut_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_5_lut_LC_13_21_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_5_lut_LC_13_21_3  (
            .in0(N__41378),
            .in1(N__30843),
            .in2(_gnd_net_),
            .in3(N__30820),
            .lcout(\c0.tx.n23963 ),
            .ltout(),
            .carryin(\c0.tx.n19542 ),
            .carryout(\c0.tx.n19543 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_6_lut_LC_13_21_4 .C_ON=1'b1;
    defparam \c0.tx.add_59_6_lut_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_6_lut_LC_13_21_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_6_lut_LC_13_21_4  (
            .in0(N__41375),
            .in1(N__30817),
            .in2(_gnd_net_),
            .in3(N__30784),
            .lcout(\c0.tx.n23953 ),
            .ltout(),
            .carryin(\c0.tx.n19543 ),
            .carryout(\c0.tx.n19544 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_7_lut_LC_13_21_5 .C_ON=1'b1;
    defparam \c0.tx.add_59_7_lut_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_7_lut_LC_13_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_7_lut_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(N__30780),
            .in2(_gnd_net_),
            .in3(N__30754),
            .lcout(n316),
            .ltout(),
            .carryin(\c0.tx.n19544 ),
            .carryout(\c0.tx.n19545 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_8_lut_LC_13_21_6 .C_ON=1'b1;
    defparam \c0.tx.add_59_8_lut_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_8_lut_LC_13_21_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_8_lut_LC_13_21_6  (
            .in0(N__41373),
            .in1(N__41546),
            .in2(_gnd_net_),
            .in3(N__31051),
            .lcout(\c0.tx.n23987 ),
            .ltout(),
            .carryin(\c0.tx.n19545 ),
            .carryout(\c0.tx.n19546 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_9_lut_LC_13_21_7 .C_ON=1'b1;
    defparam \c0.tx.add_59_9_lut_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_9_lut_LC_13_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_9_lut_LC_13_21_7  (
            .in0(_gnd_net_),
            .in1(N__31048),
            .in2(_gnd_net_),
            .in3(N__31015),
            .lcout(n314),
            .ltout(),
            .carryin(\c0.tx.n19546 ),
            .carryout(\c0.tx.n19547 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_10_lut_LC_13_22_0 .C_ON=1'b0;
    defparam \c0.tx.add_59_10_lut_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_10_lut_LC_13_22_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.tx.add_59_10_lut_LC_13_22_0  (
            .in0(N__41344),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31012),
            .lcout(n313),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1585_LC_13_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1585_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1585_LC_13_22_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_1585_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(N__68638),
            .in2(_gnd_net_),
            .in3(N__42643),
            .lcout(\c0.n12878 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i27_LC_13_23_7 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i27_LC_13_23_7 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i27_LC_13_23_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i27_LC_13_23_7  (
            .in0(_gnd_net_),
            .in1(N__34279),
            .in2(_gnd_net_),
            .in3(N__52869),
            .lcout(\c0.FRAME_MATCHER_state_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66814),
            .ce(),
            .sr(N__34264));
    defparam \c0.FRAME_MATCHER_state_i9_LC_13_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i9_LC_13_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i9_LC_13_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i9_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__37545),
            .in2(_gnd_net_),
            .in3(N__52871),
            .lcout(\c0.FRAME_MATCHER_state_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66827),
            .ce(),
            .sr(N__37582));
    defparam \c0.FRAME_MATCHER_state_i16_LC_13_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i16_LC_13_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i16_LC_13_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i16_LC_13_25_0  (
            .in0(_gnd_net_),
            .in1(N__37881),
            .in2(_gnd_net_),
            .in3(N__52872),
            .lcout(\c0.FRAME_MATCHER_state_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66839),
            .ce(),
            .sr(N__31003));
    defparam \c0.FRAME_MATCHER_state_i14_LC_13_27_5 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i14_LC_13_27_5 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i14_LC_13_27_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i14_LC_13_27_5  (
            .in0(_gnd_net_),
            .in1(N__34565),
            .in2(_gnd_net_),
            .in3(N__52889),
            .lcout(\c0.FRAME_MATCHER_state_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66858),
            .ce(),
            .sr(N__30988));
    defparam \c0.i2_2_lut_4_lut_adj_1879_LC_14_7_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_adj_1879_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_adj_1879_LC_14_7_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_2_lut_4_lut_adj_1879_LC_14_7_2  (
            .in0(N__34387),
            .in1(N__31687),
            .in2(N__31416),
            .in3(N__30982),
            .lcout(\c0.n6_adj_4305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i64_4_lut_LC_14_7_3 .C_ON=1'b0;
    defparam \c0.i64_4_lut_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.i64_4_lut_LC_14_7_3 .LUT_INIT=16'b0010111010001011;
    LogicCell40 \c0.i64_4_lut_LC_14_7_3  (
            .in0(N__31852),
            .in1(N__34386),
            .in2(N__31504),
            .in3(N__31969),
            .lcout(\c0.n21050 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1842_LC_14_7_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1842_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1842_LC_14_7_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1842_LC_14_7_4  (
            .in0(N__32518),
            .in1(N__31468),
            .in2(N__31693),
            .in3(N__31989),
            .lcout(\c0.n20658 ),
            .ltout(\c0.n20658_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1844_LC_14_7_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1844_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1844_LC_14_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1844_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(N__31457),
            .in2(N__31441),
            .in3(N__32109),
            .lcout(\c0.n22166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1709_LC_14_7_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1709_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1709_LC_14_7_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1709_LC_14_7_6  (
            .in0(N__34388),
            .in1(N__31707),
            .in2(N__31417),
            .in3(N__31635),
            .lcout(\c0.n21811 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1412_LC_14_8_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1412_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1412_LC_14_8_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1412_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__31350),
            .in2(_gnd_net_),
            .in3(N__31294),
            .lcout(\c0.n21168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1410_LC_14_8_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1410_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1410_LC_14_8_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_3_lut_adj_1410_LC_14_8_1  (
            .in0(N__31159),
            .in1(_gnd_net_),
            .in2(N__33064),
            .in3(N__31128),
            .lcout(\c0.n20298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1404_LC_14_8_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1404_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1404_LC_14_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1404_LC_14_8_2  (
            .in0(N__31213),
            .in1(N__33060),
            .in2(_gnd_net_),
            .in3(N__31158),
            .lcout(\c0.n22736 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1487_LC_14_8_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1487_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1487_LC_14_8_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_3_lut_adj_1487_LC_14_8_6  (
            .in0(N__31129),
            .in1(N__34455),
            .in2(_gnd_net_),
            .in3(N__32641),
            .lcout(\c0.n21135 ),
            .ltout(\c0.n21135_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1794_LC_14_8_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1794_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1794_LC_14_8_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_1794_LC_14_8_7  (
            .in0(N__31093),
            .in1(N__31072),
            .in2(N__31054),
            .in3(N__31565),
            .lcout(\c0.n23260 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1790_LC_14_9_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1790_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1790_LC_14_9_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1790_LC_14_9_0  (
            .in0(N__31729),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31527),
            .lcout(),
            .ltout(\c0.n6_adj_4497_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__6__5287_LC_14_9_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__6__5287_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__6__5287_LC_14_9_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame_29__6__5287_LC_14_9_1  (
            .in0(N__31537),
            .in1(N__31720),
            .in2(N__31801),
            .in3(N__31797),
            .lcout(\c0.data_out_frame_29_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66645),
            .ce(N__40946),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1588_LC_14_9_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1588_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1588_LC_14_9_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1588_LC_14_9_2  (
            .in0(N__31771),
            .in1(N__35605),
            .in2(N__32385),
            .in3(N__31536),
            .lcout(\c0.n21852 ),
            .ltout(\c0.n21852_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1827_LC_14_9_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1827_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1827_LC_14_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1827_LC_14_9_3  (
            .in0(N__32323),
            .in1(N__31741),
            .in2(N__31732),
            .in3(N__31728),
            .lcout(),
            .ltout(\c0.n10_adj_4512_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1828_LC_14_9_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1828_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1828_LC_14_9_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1828_LC_14_9_4  (
            .in0(N__31719),
            .in1(N__31708),
            .in2(N__31696),
            .in3(N__31515),
            .lcout(\c0.n20201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1488_LC_14_9_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1488_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1488_LC_14_9_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1488_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__31692),
            .in2(_gnd_net_),
            .in3(N__31623),
            .lcout(),
            .ltout(\c0.n21162_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1816_LC_14_9_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1816_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1816_LC_14_9_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1816_LC_14_9_6  (
            .in0(N__31582),
            .in1(N__31561),
            .in2(N__31540),
            .in3(N__32626),
            .lcout(\c0.n12526 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__7__5286_LC_14_9_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__7__5286_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__7__5286_LC_14_9_7 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.data_out_frame_29__7__5286_LC_14_9_7  (
            .in0(N__31528),
            .in1(_gnd_net_),
            .in2(N__31519),
            .in3(N__32561),
            .lcout(\c0.data_out_frame_29_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66645),
            .ce(N__40946),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__7__5414_LC_14_10_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__7__5414_LC_14_10_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__7__5414_LC_14_10_0 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_frame_13__7__5414_LC_14_10_0  (
            .in0(N__49322),
            .in1(N__32064),
            .in2(N__34933),
            .in3(N__48980),
            .lcout(data_out_frame_13_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66652),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1812_LC_14_10_1 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1812_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1812_LC_14_10_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_1812_LC_14_10_1  (
            .in0(N__32246),
            .in1(N__32002),
            .in2(N__32050),
            .in3(N__32013),
            .lcout(\c0.n20_adj_4505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1620_LC_14_10_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1620_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1620_LC_14_10_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1620_LC_14_10_2  (
            .in0(N__33057),
            .in1(N__32446),
            .in2(_gnd_net_),
            .in3(N__32141),
            .lcout(\c0.n22072 ),
            .ltout(\c0.n22072_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1619_LC_14_10_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1619_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1619_LC_14_10_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1619_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(N__31912),
            .in2(N__31996),
            .in3(N__32100),
            .lcout(\c0.n22073 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1647_LC_14_10_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1647_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1647_LC_14_10_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1647_LC_14_10_4  (
            .in0(N__33058),
            .in1(N__31894),
            .in2(N__32384),
            .in3(N__31968),
            .lcout(\c0.n20249 ),
            .ltout(\c0.n20249_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1726_LC_14_10_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1726_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1726_LC_14_10_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1726_LC_14_10_5  (
            .in0(N__32247),
            .in1(N__32554),
            .in2(N__31930),
            .in3(N__32512),
            .lcout(\c0.n12528 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1395_LC_14_10_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1395_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1395_LC_14_10_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1395_LC_14_10_6  (
            .in0(_gnd_net_),
            .in1(N__32373),
            .in2(_gnd_net_),
            .in3(N__31893),
            .lcout(\c0.n21842 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1850_LC_14_10_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1850_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1850_LC_14_10_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i1_2_lut_adj_1850_LC_14_10_7  (
            .in0(N__32447),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33059),
            .lcout(\c0.n20230 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1611_LC_14_11_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1611_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1611_LC_14_11_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1611_LC_14_11_0  (
            .in0(N__34978),
            .in1(N__35134),
            .in2(N__32724),
            .in3(N__34927),
            .lcout(\c0.n6_adj_4394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1869_LC_14_11_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1869_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1869_LC_14_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1869_LC_14_11_1  (
            .in0(N__35135),
            .in1(N__38296),
            .in2(_gnd_net_),
            .in3(N__32704),
            .lcout(),
            .ltout(\c0.n22163_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1813_LC_14_11_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1813_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1813_LC_14_11_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_1813_LC_14_11_2  (
            .in0(N__34979),
            .in1(N__34857),
            .in2(N__32653),
            .in3(N__34792),
            .lcout(),
            .ltout(\c0.n19_adj_4506_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1815_LC_14_11_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1815_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1815_LC_14_11_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1815_LC_14_11_3  (
            .in0(N__32572),
            .in1(N__32650),
            .in2(N__32644),
            .in3(N__32637),
            .lcout(\c0.n6_adj_4508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1814_LC_14_11_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1814_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1814_LC_14_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1814_LC_14_11_4  (
            .in0(N__32616),
            .in1(N__32593),
            .in2(N__35064),
            .in3(N__33050),
            .lcout(\c0.n21_adj_4507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1881_LC_14_11_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1881_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1881_LC_14_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1881_LC_14_11_7  (
            .in0(N__32553),
            .in1(N__32494),
            .in2(_gnd_net_),
            .in3(N__32442),
            .lcout(\c0.n21253 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1851_LC_14_12_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1851_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1851_LC_14_12_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1851_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__32372),
            .in2(_gnd_net_),
            .in3(N__32919),
            .lcout(\c0.n22078 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1877_LC_14_12_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1877_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1877_LC_14_12_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1877_LC_14_12_1  (
            .in0(N__35208),
            .in1(N__32816),
            .in2(N__32309),
            .in3(N__32233),
            .lcout(\c0.n20180 ),
            .ltout(\c0.n20180_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1890_LC_14_12_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1890_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1890_LC_14_12_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1890_LC_14_12_2  (
            .in0(N__32186),
            .in1(N__33056),
            .in2(N__32152),
            .in3(N__32135),
            .lcout(\c0.n20465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1710_LC_14_12_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1710_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1710_LC_14_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1710_LC_14_12_4  (
            .in0(N__35201),
            .in1(N__32918),
            .in2(N__33084),
            .in3(N__32852),
            .lcout(\c0.n21196 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1437_LC_14_12_5 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1437_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1437_LC_14_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1437_LC_14_12_5  (
            .in0(N__35568),
            .in1(N__39488),
            .in2(N__33018),
            .in3(N__35401),
            .lcout(\c0.n20232 ),
            .ltout(\c0.n20232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1439_LC_14_12_6 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1439_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1439_LC_14_12_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.i1_3_lut_adj_1439_LC_14_12_6  (
            .in0(N__32955),
            .in1(_gnd_net_),
            .in2(N__32935),
            .in3(N__35590),
            .lcout(\c0.n21146 ),
            .ltout(\c0.n21146_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1440_LC_14_12_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1440_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1440_LC_14_12_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1440_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32905),
            .in3(N__35200),
            .lcout(\c0.n22483 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1417_LC_14_13_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1417_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1417_LC_14_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1417_LC_14_13_0  (
            .in0(N__32902),
            .in1(N__36058),
            .in2(N__38149),
            .in3(N__32845),
            .lcout(\c0.n20744 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i27_LC_14_13_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i27_LC_14_13_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i27_LC_14_13_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i27_LC_14_13_1  (
            .in0(N__33366),
            .in1(N__42248),
            .in2(_gnd_net_),
            .in3(N__33343),
            .lcout(encoder0_position_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66674),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i1_LC_14_13_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i1_LC_14_13_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i1_LC_14_13_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \quad_counter0.count_i0_i1_LC_14_13_2  (
            .in0(N__33121),
            .in1(_gnd_net_),
            .in2(N__42252),
            .in3(N__35765),
            .lcout(encoder0_position_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66674),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__1__5420_LC_14_13_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__1__5420_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__1__5420_LC_14_13_3 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_frame_13__1__5420_LC_14_13_3  (
            .in0(N__49272),
            .in1(N__34731),
            .in2(N__32800),
            .in3(N__48895),
            .lcout(data_out_frame_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66674),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i20_LC_14_13_4 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i20_LC_14_13_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i20_LC_14_13_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \quad_counter0.count_i0_i20_LC_14_13_4  (
            .in0(N__33277),
            .in1(_gnd_net_),
            .in2(N__42253),
            .in3(N__36121),
            .lcout(encoder0_position_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66674),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i13_LC_14_13_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i13_LC_14_13_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i13_LC_14_13_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter0.count_i0_i13_LC_14_13_5  (
            .in0(N__33175),
            .in1(N__42240),
            .in2(_gnd_net_),
            .in3(N__35713),
            .lcout(encoder0_position_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66674),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i14_LC_14_13_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i14_LC_14_13_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i14_LC_14_13_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \quad_counter0.count_i0_i14_LC_14_13_6  (
            .in0(N__42241),
            .in1(_gnd_net_),
            .in2(N__35890),
            .in3(N__33310),
            .lcout(encoder0_position_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66674),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1862_LC_14_13_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1862_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1862_LC_14_13_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1862_LC_14_13_7  (
            .in0(N__38257),
            .in1(N__35877),
            .in2(N__33376),
            .in3(N__35812),
            .lcout(\c0.n20160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_1_LC_14_14_0 .C_ON=1'b1;
    defparam \quad_counter0.add_645_1_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_1_LC_14_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \quad_counter0.add_645_1_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__33606),
            .in2(N__33679),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\quad_counter0.n19580 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_2_lut_LC_14_14_1 .C_ON=1'b1;
    defparam \quad_counter0.add_645_2_lut_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_2_lut_LC_14_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_2_lut_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__37046),
            .in2(N__33145),
            .in3(N__33124),
            .lcout(n2271),
            .ltout(),
            .carryin(\quad_counter0.n19580 ),
            .carryout(\quad_counter0.n19581 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_3_lut_LC_14_14_2 .C_ON=1'b1;
    defparam \quad_counter0.add_645_3_lut_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_3_lut_LC_14_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_3_lut_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__35764),
            .in2(N__33680),
            .in3(N__33115),
            .lcout(n2270),
            .ltout(),
            .carryin(\quad_counter0.n19581 ),
            .carryout(\quad_counter0.n19582 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_4_lut_LC_14_14_3 .C_ON=1'b1;
    defparam \quad_counter0.add_645_4_lut_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_4_lut_LC_14_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_4_lut_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__53457),
            .in2(N__33676),
            .in3(N__33106),
            .lcout(n2269),
            .ltout(),
            .carryin(\quad_counter0.n19582 ),
            .carryout(\quad_counter0.n19583 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_5_lut_LC_14_14_4 .C_ON=1'b1;
    defparam \quad_counter0.add_645_5_lut_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_5_lut_LC_14_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_5_lut_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__41696),
            .in2(N__33681),
            .in3(N__33091),
            .lcout(n2268),
            .ltout(),
            .carryin(\quad_counter0.n19583 ),
            .carryout(\quad_counter0.n19584 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_6_lut_LC_14_14_5 .C_ON=1'b1;
    defparam \quad_counter0.add_645_6_lut_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_6_lut_LC_14_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_6_lut_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__39036),
            .in2(N__33677),
            .in3(N__33088),
            .lcout(n2267),
            .ltout(),
            .carryin(\quad_counter0.n19584 ),
            .carryout(\quad_counter0.n19585 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_7_lut_LC_14_14_6 .C_ON=1'b1;
    defparam \quad_counter0.add_645_7_lut_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_7_lut_LC_14_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_7_lut_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__36062),
            .in2(N__33682),
            .in3(N__33259),
            .lcout(n2266),
            .ltout(),
            .carryin(\quad_counter0.n19585 ),
            .carryout(\quad_counter0.n19586 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_8_lut_LC_14_14_7 .C_ON=1'b1;
    defparam \quad_counter0.add_645_8_lut_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_8_lut_LC_14_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_8_lut_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(N__36159),
            .in2(N__33678),
            .in3(N__33256),
            .lcout(n2265),
            .ltout(),
            .carryin(\quad_counter0.n19586 ),
            .carryout(\quad_counter0.n19587 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_9_lut_LC_14_15_0 .C_ON=1'b1;
    defparam \quad_counter0.add_645_9_lut_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_9_lut_LC_14_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_9_lut_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__33628),
            .in2(N__33245),
            .in3(N__33193),
            .lcout(n2264),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\quad_counter0.n19588 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_10_lut_LC_14_15_1 .C_ON=1'b1;
    defparam \quad_counter0.add_645_10_lut_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_10_lut_LC_14_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_10_lut_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__40305),
            .in2(N__33683),
            .in3(N__33190),
            .lcout(n2263),
            .ltout(),
            .carryin(\quad_counter0.n19588 ),
            .carryout(\quad_counter0.n19589 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_11_lut_LC_14_15_2 .C_ON=1'b1;
    defparam \quad_counter0.add_645_11_lut_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_11_lut_LC_14_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_11_lut_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__33632),
            .in2(N__38723),
            .in3(N__33187),
            .lcout(n2262),
            .ltout(),
            .carryin(\quad_counter0.n19589 ),
            .carryout(\quad_counter0.n19590 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_12_lut_LC_14_15_3 .C_ON=1'b1;
    defparam \quad_counter0.add_645_12_lut_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_12_lut_LC_14_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_12_lut_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__39975),
            .in2(N__33684),
            .in3(N__33184),
            .lcout(n2261),
            .ltout(),
            .carryin(\quad_counter0.n19590 ),
            .carryout(\quad_counter0.n19591 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_13_lut_LC_14_15_4 .C_ON=1'b1;
    defparam \quad_counter0.add_645_13_lut_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_13_lut_LC_14_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_13_lut_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__33636),
            .in2(N__39394),
            .in3(N__33181),
            .lcout(n2260),
            .ltout(),
            .carryin(\quad_counter0.n19591 ),
            .carryout(\quad_counter0.n19592 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_14_lut_LC_14_15_5 .C_ON=1'b1;
    defparam \quad_counter0.add_645_14_lut_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_14_lut_LC_14_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_14_lut_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__38869),
            .in2(N__33685),
            .in3(N__33178),
            .lcout(n2259),
            .ltout(),
            .carryin(\quad_counter0.n19592 ),
            .carryout(\quad_counter0.n19593 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_15_lut_LC_14_15_6 .C_ON=1'b1;
    defparam \quad_counter0.add_645_15_lut_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_15_lut_LC_14_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_15_lut_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(N__33640),
            .in2(N__35724),
            .in3(N__33166),
            .lcout(n2258),
            .ltout(),
            .carryin(\quad_counter0.n19593 ),
            .carryout(\quad_counter0.n19594 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_16_lut_LC_14_15_7 .C_ON=1'b1;
    defparam \quad_counter0.add_645_16_lut_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_16_lut_LC_14_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_16_lut_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__35891),
            .in2(N__33686),
            .in3(N__33301),
            .lcout(n2257),
            .ltout(),
            .carryin(\quad_counter0.n19594 ),
            .carryout(\quad_counter0.n19595 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_17_lut_LC_14_16_0 .C_ON=1'b1;
    defparam \quad_counter0.add_645_17_lut_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_17_lut_LC_14_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_17_lut_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__36252),
            .in2(N__33691),
            .in3(N__33298),
            .lcout(n2256),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\quad_counter0.n19596 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_18_lut_LC_14_16_1 .C_ON=1'b1;
    defparam \quad_counter0.add_645_18_lut_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_18_lut_LC_14_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_18_lut_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__33663),
            .in2(N__39114),
            .in3(N__33295),
            .lcout(n2255),
            .ltout(),
            .carryin(\quad_counter0.n19596 ),
            .carryout(\quad_counter0.n19597 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_19_lut_LC_14_16_2 .C_ON=1'b1;
    defparam \quad_counter0.add_645_19_lut_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_19_lut_LC_14_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_19_lut_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__33664),
            .in2(N__36556),
            .in3(N__33292),
            .lcout(n2254),
            .ltout(),
            .carryin(\quad_counter0.n19597 ),
            .carryout(\quad_counter0.n19598 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_20_lut_LC_14_16_3 .C_ON=1'b1;
    defparam \quad_counter0.add_645_20_lut_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_20_lut_LC_14_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_20_lut_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__41754),
            .in2(N__33692),
            .in3(N__33289),
            .lcout(n2253),
            .ltout(),
            .carryin(\quad_counter0.n19598 ),
            .carryout(\quad_counter0.n19599 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_21_lut_LC_14_16_4 .C_ON=1'b1;
    defparam \quad_counter0.add_645_21_lut_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_21_lut_LC_14_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_21_lut_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__33668),
            .in2(N__38662),
            .in3(N__33280),
            .lcout(n2252),
            .ltout(),
            .carryin(\quad_counter0.n19599 ),
            .carryout(\quad_counter0.n19600 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_22_lut_LC_14_16_5 .C_ON=1'b1;
    defparam \quad_counter0.add_645_22_lut_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_22_lut_LC_14_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_22_lut_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__36123),
            .in2(N__33693),
            .in3(N__33268),
            .lcout(n2251),
            .ltout(),
            .carryin(\quad_counter0.n19600 ),
            .carryout(\quad_counter0.n19601 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_23_lut_LC_14_16_6 .C_ON=1'b1;
    defparam \quad_counter0.add_645_23_lut_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_23_lut_LC_14_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_23_lut_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__33672),
            .in2(N__35993),
            .in3(N__33265),
            .lcout(n2250),
            .ltout(),
            .carryin(\quad_counter0.n19601 ),
            .carryout(\quad_counter0.n19602 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_24_lut_LC_14_16_7 .C_ON=1'b1;
    defparam \quad_counter0.add_645_24_lut_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_24_lut_LC_14_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_24_lut_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(N__42045),
            .in2(N__33694),
            .in3(N__33262),
            .lcout(n2249),
            .ltout(),
            .carryin(\quad_counter0.n19602 ),
            .carryout(\quad_counter0.n19603 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_25_lut_LC_14_17_0 .C_ON=1'b1;
    defparam \quad_counter0.add_645_25_lut_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_25_lut_LC_14_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_25_lut_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__33644),
            .in2(N__40366),
            .in3(N__33406),
            .lcout(n2248),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\quad_counter0.n19604 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_26_lut_LC_14_17_1 .C_ON=1'b1;
    defparam \quad_counter0.add_645_26_lut_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_26_lut_LC_14_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_26_lut_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__39320),
            .in2(N__33687),
            .in3(N__33403),
            .lcout(n2247),
            .ltout(),
            .carryin(\quad_counter0.n19604 ),
            .carryout(\quad_counter0.n19605 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_27_lut_LC_14_17_2 .C_ON=1'b1;
    defparam \quad_counter0.add_645_27_lut_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_27_lut_LC_14_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_27_lut_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__33648),
            .in2(N__39907),
            .in3(N__33400),
            .lcout(n2246),
            .ltout(),
            .carryin(\quad_counter0.n19605 ),
            .carryout(\quad_counter0.n19606 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_28_lut_LC_14_17_3 .C_ON=1'b1;
    defparam \quad_counter0.add_645_28_lut_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_28_lut_LC_14_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_28_lut_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__40059),
            .in2(N__33688),
            .in3(N__33397),
            .lcout(n2245),
            .ltout(),
            .carryin(\quad_counter0.n19606 ),
            .carryout(\quad_counter0.n19607 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_29_lut_LC_14_17_4 .C_ON=1'b1;
    defparam \quad_counter0.add_645_29_lut_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_29_lut_LC_14_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_29_lut_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(N__33652),
            .in2(N__33387),
            .in3(N__33334),
            .lcout(n2244),
            .ltout(),
            .carryin(\quad_counter0.n19607 ),
            .carryout(\quad_counter0.n19608 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_30_lut_LC_14_17_5 .C_ON=1'b1;
    defparam \quad_counter0.add_645_30_lut_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_30_lut_LC_14_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_30_lut_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__38784),
            .in2(N__33689),
            .in3(N__33331),
            .lcout(n2243),
            .ltout(),
            .carryin(\quad_counter0.n19608 ),
            .carryout(\quad_counter0.n19609 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_31_lut_LC_14_17_6 .C_ON=1'b1;
    defparam \quad_counter0.add_645_31_lut_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_31_lut_LC_14_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_31_lut_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(N__33656),
            .in2(N__38248),
            .in3(N__33328),
            .lcout(n2242),
            .ltout(),
            .carryin(\quad_counter0.n19609 ),
            .carryout(\quad_counter0.n19610 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_32_lut_LC_14_17_7 .C_ON=1'b1;
    defparam \quad_counter0.add_645_32_lut_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_32_lut_LC_14_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_645_32_lut_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__48551),
            .in2(N__33690),
            .in3(N__33313),
            .lcout(n2241),
            .ltout(),
            .carryin(\quad_counter0.n19610 ),
            .carryout(\quad_counter0.n19611 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_645_33_lut_LC_14_18_0 .C_ON=1'b0;
    defparam \quad_counter0.add_645_33_lut_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_645_33_lut_LC_14_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \quad_counter0.add_645_33_lut_LC_14_18_0  (
            .in0(N__41628),
            .in1(N__33605),
            .in2(_gnd_net_),
            .in3(N__33496),
            .lcout(n2240),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1390_LC_14_18_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1390_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1390_LC_14_18_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1390_LC_14_18_1  (
            .in0(N__37945),
            .in1(N__37468),
            .in2(_gnd_net_),
            .in3(N__37501),
            .lcout(),
            .ltout(\c0.n14474_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18960_4_lut_LC_14_18_2 .C_ON=1'b0;
    defparam \c0.i18960_4_lut_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i18960_4_lut_LC_14_18_2 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \c0.i18960_4_lut_LC_14_18_2  (
            .in0(N__37502),
            .in1(N__42506),
            .in2(N__33493),
            .in3(N__37409),
            .lcout(\c0.n22651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__1__5452_LC_14_18_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__1__5452_LC_14_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__1__5452_LC_14_18_3 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_9__1__5452_LC_14_18_3  (
            .in0(N__49450),
            .in1(N__48743),
            .in2(N__35776),
            .in3(N__33490),
            .lcout(data_out_frame_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66742),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n24183_bdd_4_lut_LC_14_18_4 .C_ON=1'b0;
    defparam \c0.n24183_bdd_4_lut_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.n24183_bdd_4_lut_LC_14_18_4 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n24183_bdd_4_lut_LC_14_18_4  (
            .in0(N__33489),
            .in1(N__36652),
            .in2(N__33481),
            .in3(N__36890),
            .lcout(\c0.n24186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i23_LC_14_18_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i23_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i23_LC_14_18_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i23_LC_14_18_5  (
            .in0(N__42106),
            .in1(N__33448),
            .in2(_gnd_net_),
            .in3(N__40355),
            .lcout(encoder0_position_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66742),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i31_LC_14_18_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i31_LC_14_18_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i31_LC_14_18_6 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \quad_counter0.count_i0_i31_LC_14_18_6  (
            .in0(N__42107),
            .in1(N__33442),
            .in2(N__41645),
            .in3(_gnd_net_),
            .lcout(encoder0_position_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66742),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__7__5462_LC_14_18_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__7__5462_LC_14_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__7__5462_LC_14_18_7 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_7__7__5462_LC_14_18_7  (
            .in0(N__49449),
            .in1(N__48742),
            .in2(N__40367),
            .in3(N__33432),
            .lcout(data_out_frame_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66742),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__1__5484_LC_14_19_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__1__5484_LC_14_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__1__5484_LC_14_19_0 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_out_frame_5__1__5484_LC_14_19_0  (
            .in0(N__48737),
            .in1(N__49455),
            .in2(N__33418),
            .in3(N__41870),
            .lcout(data_out_frame_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66756),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20396_3_lut_LC_14_19_1 .C_ON=1'b0;
    defparam \c0.i20396_3_lut_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i20396_3_lut_LC_14_19_1 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \c0.i20396_3_lut_LC_14_19_1  (
            .in0(N__33944),
            .in1(N__33414),
            .in2(_gnd_net_),
            .in3(N__39815),
            .lcout(\c0.n24093 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1204_LC_14_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1204_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1204_LC_14_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1204_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__44929),
            .in2(_gnd_net_),
            .in3(N__59353),
            .lcout(\c0.n22358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__1__5468_LC_14_19_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__1__5468_LC_14_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__1__5468_LC_14_19_3 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_7__1__5468_LC_14_19_3  (
            .in0(N__49453),
            .in1(N__48739),
            .in2(N__34009),
            .in3(N__36559),
            .lcout(data_out_frame_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66756),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__7__5478_LC_14_19_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__7__5478_LC_14_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__7__5478_LC_14_19_4 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_5__7__5478_LC_14_19_4  (
            .in0(N__48738),
            .in1(N__49456),
            .in2(N__42352),
            .in3(N__33804),
            .lcout(data_out_frame_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66756),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__0__5461_LC_14_19_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__0__5461_LC_14_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__0__5461_LC_14_19_5 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_8__0__5461_LC_14_19_5  (
            .in0(N__49454),
            .in1(N__48740),
            .in2(N__40312),
            .in3(N__34023),
            .lcout(data_out_frame_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66756),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_14_19_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_14_19_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_14_19_6  (
            .in0(N__39816),
            .in1(N__34005),
            .in2(_gnd_net_),
            .in3(N__37083),
            .lcout(),
            .ltout(\c0.n5_adj_4518_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20167_4_lut_LC_14_19_7 .C_ON=1'b0;
    defparam \c0.i20167_4_lut_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i20167_4_lut_LC_14_19_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \c0.i20167_4_lut_LC_14_19_7  (
            .in0(N__33945),
            .in1(N__33997),
            .in2(N__33991),
            .in3(N__36909),
            .lcout(\c0.n23862 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1682_LC_14_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1682_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1682_LC_14_20_0 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1682_LC_14_20_0  (
            .in0(N__68570),
            .in1(N__46148),
            .in2(_gnd_net_),
            .in3(N__42639),
            .lcout(\c0.n20_adj_4327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20358_3_lut_LC_14_20_2 .C_ON=1'b0;
    defparam \c0.i20358_3_lut_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i20358_3_lut_LC_14_20_2 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \c0.i20358_3_lut_LC_14_20_2  (
            .in0(N__39814),
            .in1(N__33943),
            .in2(_gnd_net_),
            .in3(N__33805),
            .lcout(\c0.n24054 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i3737_2_lut_LC_14_20_3 .C_ON=1'b0;
    defparam \c0.tx.i3737_2_lut_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i3737_2_lut_LC_14_20_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.tx.i3737_2_lut_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__33770),
            .in2(_gnd_net_),
            .in3(N__39269),
            .lcout(\c0.tx.n7086 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1389_LC_14_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1389_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1389_LC_14_20_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1389_LC_14_20_4  (
            .in0(N__37469),
            .in1(N__37424),
            .in2(_gnd_net_),
            .in3(N__37494),
            .lcout(\c0.n9668 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1900_LC_14_20_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1900_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1900_LC_14_20_5 .LUT_INIT=16'b1000000011110000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1900_LC_14_20_5  (
            .in0(N__37495),
            .in1(N__37389),
            .in2(N__37432),
            .in3(N__37470),
            .lcout(data_out_frame_29_7_N_1483_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i12_LC_14_20_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i12_LC_14_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i12_LC_14_20_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i12_LC_14_20_6  (
            .in0(N__43263),
            .in1(N__34198),
            .in2(_gnd_net_),
            .in3(N__36367),
            .lcout(data_in_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66770),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i18_LC_14_20_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i18_LC_14_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i18_LC_14_20_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i18_LC_14_20_7  (
            .in0(N__43264),
            .in1(N__34157),
            .in2(_gnd_net_),
            .in3(N__43043),
            .lcout(data_in_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66770),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1872_LC_14_21_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1872_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1872_LC_14_21_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i5_4_lut_adj_1872_LC_14_21_4  (
            .in0(N__34542),
            .in1(N__34129),
            .in2(N__41155),
            .in3(N__34036),
            .lcout(\c0.n13_adj_4388 ),
            .ltout(\c0.n13_adj_4388_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1887_LC_14_21_5 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1887_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1887_LC_14_21_5 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \c0.i1_3_lut_adj_1887_LC_14_21_5  (
            .in0(N__37819),
            .in1(_gnd_net_),
            .in2(N__34132),
            .in3(N__37620),
            .lcout(\c0.n21789 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1393_LC_14_22_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1393_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1393_LC_14_22_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_1393_LC_14_22_1  (
            .in0(N__43539),
            .in1(N__34308),
            .in2(N__37335),
            .in3(N__37753),
            .lcout(\c0.n23135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i11_4_lut_LC_14_22_2 .C_ON=1'b0;
    defparam \quad_counter0.i11_4_lut_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i11_4_lut_LC_14_22_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i11_4_lut_LC_14_22_2  (
            .in0(N__34123),
            .in1(N__34105),
            .in2(N__34087),
            .in3(N__34066),
            .lcout(\quad_counter0.n27_adj_4200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1358_LC_14_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1358_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1358_LC_14_22_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_1358_LC_14_22_3  (
            .in0(_gnd_net_),
            .in1(N__34277),
            .in2(_gnd_net_),
            .in3(N__34503),
            .lcout(\c0.n14457 ),
            .ltout(\c0.n14457_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_adj_1645_LC_14_22_4 .C_ON=1'b0;
    defparam \c0.i21_4_lut_adj_1645_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_adj_1645_LC_14_22_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i21_4_lut_adj_1645_LC_14_22_4  (
            .in0(N__34309),
            .in1(N__41053),
            .in2(N__34282),
            .in3(N__41007),
            .lcout(\c0.n49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1774_LC_14_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1774_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1774_LC_14_22_5 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1774_LC_14_22_5  (
            .in0(N__37609),
            .in1(N__53193),
            .in2(_gnd_net_),
            .in3(N__52947),
            .lcout(\c0.n21372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1522_LC_14_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1522_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1522_LC_14_22_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_1522_LC_14_22_6  (
            .in0(N__34278),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40652),
            .lcout(\c0.n21330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1526_LC_14_22_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1526_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1526_LC_14_22_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_1526_LC_14_22_7  (
            .in0(N__40653),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34504),
            .lcout(\c0.n21326 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1635_LC_14_23_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1635_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1635_LC_14_23_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i2_2_lut_adj_1635_LC_14_23_0  (
            .in0(_gnd_net_),
            .in1(N__37914),
            .in2(_gnd_net_),
            .in3(N__43455),
            .lcout(),
            .ltout(\c0.n30_adj_4411_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_LC_14_23_1 .C_ON=1'b0;
    defparam \c0.i22_4_lut_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_LC_14_23_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i22_4_lut_LC_14_23_1  (
            .in0(N__41151),
            .in1(N__34576),
            .in2(N__34252),
            .in3(N__34248),
            .lcout(\c0.n50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1751_LC_14_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1751_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1751_LC_14_23_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1751_LC_14_23_3  (
            .in0(N__52974),
            .in1(N__34249),
            .in2(_gnd_net_),
            .in3(N__53170),
            .lcout(\c0.n21344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1778_LC_14_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1778_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1778_LC_14_23_4 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1778_LC_14_23_4  (
            .in0(N__53169),
            .in1(N__42547),
            .in2(N__37803),
            .in3(N__42767),
            .lcout(\c0.n21336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1746_LC_14_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1746_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1746_LC_14_23_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1746_LC_14_23_7  (
            .in0(N__42766),
            .in1(N__42870),
            .in2(_gnd_net_),
            .in3(N__40633),
            .lcout(\c0.n4_adj_4345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i25_LC_14_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i25_LC_14_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i25_LC_14_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i25_LC_14_24_0  (
            .in0(_gnd_net_),
            .in1(N__37752),
            .in2(_gnd_net_),
            .in3(N__52860),
            .lcout(\c0.FRAME_MATCHER_state_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66815),
            .ce(),
            .sr(N__37726));
    defparam \c0.i16_4_lut_adj_1636_LC_14_25_1 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1636_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1636_LC_14_25_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i16_4_lut_adj_1636_LC_14_25_1  (
            .in0(N__34567),
            .in1(N__37750),
            .in2(N__34543),
            .in3(N__37880),
            .lcout(\c0.n44_adj_4412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1768_LC_14_25_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1768_LC_14_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1768_LC_14_25_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1768_LC_14_25_2  (
            .in0(N__53189),
            .in1(N__34540),
            .in2(_gnd_net_),
            .in3(N__53009),
            .lcout(\c0.n21368 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1891_LC_14_25_6 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1891_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1891_LC_14_25_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_1891_LC_14_25_6  (
            .in0(N__37541),
            .in1(N__37716),
            .in2(N__42936),
            .in3(N__34566),
            .lcout(\c0.n19_adj_4481 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i21_LC_14_26_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i21_LC_14_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i21_LC_14_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i21_LC_14_26_0  (
            .in0(_gnd_net_),
            .in1(N__34541),
            .in2(_gnd_net_),
            .in3(N__52885),
            .lcout(\c0.FRAME_MATCHER_state_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66840),
            .ce(),
            .sr(N__34516));
    defparam \c0.FRAME_MATCHER_state_i29_LC_14_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i29_LC_14_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i29_LC_14_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i29_LC_14_27_0  (
            .in0(_gnd_net_),
            .in1(N__34502),
            .in2(_gnd_net_),
            .in3(N__52887),
            .lcout(\c0.FRAME_MATCHER_state_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66850),
            .ce(),
            .sr(N__34486));
    defparam \c0.i6_4_lut_adj_1623_LC_15_9_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1623_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1623_LC_15_9_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_1623_LC_15_9_0  (
            .in0(N__52183),
            .in1(N__54685),
            .in2(N__61072),
            .in3(N__48241),
            .lcout(\c0.n14_adj_4400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1795_LC_15_9_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1795_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1795_LC_15_9_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1795_LC_15_9_1  (
            .in0(N__34477),
            .in1(N__34456),
            .in2(N__34398),
            .in3(N__34366),
            .lcout(),
            .ltout(\c0.n16_adj_4498_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__7__5294_LC_15_9_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__7__5294_LC_15_9_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__7__5294_LC_15_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_28__7__5294_LC_15_9_2  (
            .in0(N__34343),
            .in1(N__34318),
            .in2(N__34312),
            .in3(N__34774),
            .lcout(\c0.data_out_frame_28_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66639),
            .ce(N__40945),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1796_LC_15_9_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1796_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1796_LC_15_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1796_LC_15_9_3  (
            .in0(N__34861),
            .in1(N__34834),
            .in2(N__34827),
            .in3(N__34801),
            .lcout(\c0.n17_adj_4499 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i26_3_lut_LC_15_9_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i26_3_lut_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i26_3_lut_LC_15_9_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_7_i26_3_lut_LC_15_9_4  (
            .in0(N__39734),
            .in1(N__34768),
            .in2(_gnd_net_),
            .in3(N__34759),
            .lcout(\c0.n26_adj_4359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_15_9_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_15_9_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_15_9_5  (
            .in0(N__34735),
            .in1(N__34717),
            .in2(_gnd_net_),
            .in3(N__39733),
            .lcout(\c0.n11_adj_4520 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1543_LC_15_10_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1543_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1543_LC_15_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i6_4_lut_adj_1543_LC_15_10_0  (
            .in0(N__50350),
            .in1(N__44165),
            .in2(N__47523),
            .in3(N__51712),
            .lcout(\c0.n14_adj_4364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i30_LC_15_10_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i30_LC_15_10_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i30_LC_15_10_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i30_LC_15_10_1  (
            .in0(N__67214),
            .in1(N__43216),
            .in2(_gnd_net_),
            .in3(N__35245),
            .lcout(data_in_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66646),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__3__5458_LC_15_10_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__3__5458_LC_15_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__3__5458_LC_15_10_2 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_frame_8__3__5458_LC_15_10_2  (
            .in0(N__49255),
            .in1(N__34668),
            .in2(N__39391),
            .in3(N__48949),
            .lcout(data_out_frame_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66646),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_15_10_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_15_10_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_15_10_3  (
            .in0(N__39732),
            .in1(N__35080),
            .in2(_gnd_net_),
            .in3(N__34584),
            .lcout(\c0.n11_adj_4303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__4__5425_LC_15_10_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__4__5425_LC_15_10_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__4__5425_LC_15_10_4 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_12__4__5425_LC_15_10_4  (
            .in0(N__49254),
            .in1(N__48947),
            .in2(N__34588),
            .in3(N__34636),
            .lcout(data_out_frame_12_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66646),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__0__5429_LC_15_10_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__0__5429_LC_15_10_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__0__5429_LC_15_10_6 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_frame_12__0__5429_LC_15_10_6  (
            .in0(N__49253),
            .in1(N__35334),
            .in2(N__35395),
            .in3(N__48948),
            .lcout(data_out_frame_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66646),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1456_LC_15_11_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1456_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1456_LC_15_11_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1456_LC_15_11_0  (
            .in0(N__34925),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35308),
            .lcout(\c0.n22174 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i22_LC_15_11_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i22_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i22_LC_15_11_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i22_LC_15_11_1  (
            .in0(N__35252),
            .in1(N__43175),
            .in2(_gnd_net_),
            .in3(N__36406),
            .lcout(data_in_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66653),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__2__5427_LC_15_11_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__2__5427_LC_15_11_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__2__5427_LC_15_11_2 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_12__2__5427_LC_15_11_2  (
            .in0(N__49269),
            .in1(N__49045),
            .in2(N__35169),
            .in3(N__35221),
            .lcout(data_out_frame_12_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66653),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1657_LC_15_11_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1657_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1657_LC_15_11_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1657_LC_15_11_3  (
            .in0(N__40057),
            .in1(N__39903),
            .in2(N__39390),
            .in3(N__42351),
            .lcout(\c0.n21918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1476_LC_15_11_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1476_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1476_LC_15_11_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1476_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__40304),
            .in2(_gnd_net_),
            .in3(N__40369),
            .lcout(\c0.n22474 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__4__5417_LC_15_11_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__4__5417_LC_15_11_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__4__5417_LC_15_11_5 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_13__4__5417_LC_15_11_5  (
            .in0(N__49044),
            .in1(N__49271),
            .in2(N__35140),
            .in3(N__35079),
            .lcout(data_out_frame_13_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66653),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__2__5419_LC_15_11_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__2__5419_LC_15_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__2__5419_LC_15_11_6 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_13__2__5419_LC_15_11_6  (
            .in0(N__49270),
            .in1(N__49046),
            .in2(N__35065),
            .in3(N__34998),
            .lcout(data_out_frame_13_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66653),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1418_LC_15_11_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1418_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1418_LC_15_11_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1418_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(N__34980),
            .in2(_gnd_net_),
            .in3(N__34926),
            .lcout(\c0.n21896 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1438_LC_15_12_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1438_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1438_LC_15_12_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1438_LC_15_12_1  (
            .in0(N__39426),
            .in1(N__40261),
            .in2(N__35655),
            .in3(N__42046),
            .lcout(\c0.n20236 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1447_LC_15_12_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1447_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1447_LC_15_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1447_LC_15_12_3  (
            .in0(N__35431),
            .in1(N__35572),
            .in2(N__35545),
            .in3(N__35536),
            .lcout(),
            .ltout(\c0.n16_adj_4321_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_adj_1448_LC_15_12_4 .C_ON=1'b0;
    defparam \c0.i8_3_lut_adj_1448_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_adj_1448_LC_15_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i8_3_lut_adj_1448_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__35529),
            .in2(N__35479),
            .in3(N__38059),
            .lcout(),
            .ltout(\c0.n18_adj_4322_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1450_LC_15_12_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1450_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1450_LC_15_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1450_LC_15_12_5  (
            .in0(N__53502),
            .in1(N__38905),
            .in2(N__35476),
            .in3(N__35473),
            .lcout(\c0.n14_adj_4324 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1826_LC_15_13_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1826_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1826_LC_15_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1826_LC_15_13_0  (
            .in0(N__38677),
            .in1(N__37263),
            .in2(N__36557),
            .in3(N__35928),
            .lcout(\c0.n22376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1465_LC_15_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1465_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1465_LC_15_13_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1465_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__35701),
            .in2(_gnd_net_),
            .in3(N__35872),
            .lcout(\c0.n13619 ),
            .ltout(\c0.n13619_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1467_LC_15_13_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1467_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1467_LC_15_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1467_LC_15_13_2  (
            .in0(N__38676),
            .in1(N__38242),
            .in2(N__35425),
            .in3(N__53409),
            .lcout(\c0.n10_adj_4331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1431_LC_15_13_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1431_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1431_LC_15_13_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1431_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__36549),
            .in2(_gnd_net_),
            .in3(N__38667),
            .lcout(),
            .ltout(\c0.n13524_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1436_LC_15_13_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1436_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1436_LC_15_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1436_LC_15_13_4  (
            .in0(N__35422),
            .in1(N__38821),
            .in2(N__35404),
            .in3(N__35824),
            .lcout(\c0.n10_adj_4317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1906_LC_15_13_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1906_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1906_LC_15_13_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1906_LC_15_13_5  (
            .in0(N__38243),
            .in1(N__38783),
            .in2(N__48570),
            .in3(N__35810),
            .lcout(\c0.n20328 ),
            .ltout(\c0.n20328_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1692_LC_15_13_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1692_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1692_LC_15_13_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1692_LC_15_13_6  (
            .in0(N__35873),
            .in1(_gnd_net_),
            .in2(N__35842),
            .in3(N__35702),
            .lcout(\c0.n22367 ),
            .ltout(\c0.n22367_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1435_LC_15_13_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1435_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1435_LC_15_13_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1435_LC_15_13_7  (
            .in0(N__38599),
            .in1(N__36027),
            .in2(N__35827),
            .in3(N__36258),
            .lcout(\c0.n23569 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1443_LC_15_14_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1443_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1443_LC_15_14_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1443_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__39014),
            .in2(_gnd_net_),
            .in3(N__36056),
            .lcout(\c0.n22230 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1442_LC_15_14_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1442_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1442_LC_15_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1442_LC_15_14_1  (
            .in0(N__36154),
            .in1(N__35979),
            .in2(_gnd_net_),
            .in3(N__42396),
            .lcout(\c0.n22382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i0_LC_15_14_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i0_LC_15_14_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i0_LC_15_14_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i0_LC_15_14_2  (
            .in0(N__42249),
            .in1(N__35818),
            .in2(_gnd_net_),
            .in3(N__37047),
            .lcout(encoder0_position_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66675),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_3_lut_4_lut_LC_15_14_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_3_lut_4_lut_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_3_lut_4_lut_LC_15_14_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_3_lut_3_lut_4_lut_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__48552),
            .in2(_gnd_net_),
            .in3(N__35811),
            .lcout(),
            .ltout(\c0.n22461_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1444_LC_15_14_4 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1444_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1444_LC_15_14_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1444_LC_15_14_4  (
            .in0(N__35787),
            .in1(N__35763),
            .in2(N__35728),
            .in3(N__35703),
            .lcout(\c0.n20_adj_4318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i6_LC_15_14_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i6_LC_15_14_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i6_LC_15_14_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i6_LC_15_14_5  (
            .in0(N__36155),
            .in1(N__42251),
            .in2(_gnd_net_),
            .in3(N__36172),
            .lcout(encoder0_position_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66675),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1472_LC_15_14_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1472_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1472_LC_15_14_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1472_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__36111),
            .in2(_gnd_net_),
            .in3(N__41799),
            .lcout(\c0.n21970 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i5_LC_15_14_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i5_LC_15_14_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i5_LC_15_14_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i5_LC_15_14_7  (
            .in0(N__36057),
            .in1(N__42250),
            .in2(_gnd_net_),
            .in3(N__36088),
            .lcout(encoder0_position_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66675),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1688_LC_15_15_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1688_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1688_LC_15_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1688_LC_15_15_0  (
            .in0(N__41648),
            .in1(N__38756),
            .in2(N__48566),
            .in3(N__39091),
            .lcout(\c0.n21808 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i21_LC_15_15_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i21_LC_15_15_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i21_LC_15_15_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i21_LC_15_15_1  (
            .in0(N__35989),
            .in1(N__36010),
            .in2(_gnd_net_),
            .in3(N__42208),
            .lcout(encoder0_position_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66687),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i9_LC_15_15_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i9_LC_15_15_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i9_LC_15_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i9_LC_15_15_2  (
            .in0(N__42209),
            .in1(N__35953),
            .in2(_gnd_net_),
            .in3(N__38722),
            .lcout(encoder0_position_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66687),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i11_LC_15_15_3 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i11_LC_15_15_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i11_LC_15_15_3 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \quad_counter0.count_i0_i11_LC_15_15_3  (
            .in0(N__35947),
            .in1(N__42204),
            .in2(N__39393),
            .in3(_gnd_net_),
            .lcout(encoder0_position_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66687),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i17_LC_15_15_4 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i17_LC_15_15_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i17_LC_15_15_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \quad_counter0.count_i0_i17_LC_15_15_4  (
            .in0(N__35938),
            .in1(_gnd_net_),
            .in2(N__42239),
            .in3(N__36531),
            .lcout(encoder0_position_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1479_LC_15_15_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1479_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1479_LC_15_15_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1479_LC_15_15_5  (
            .in0(N__44608),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41649),
            .lcout(\c0.n10394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1640_LC_15_15_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1640_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1640_LC_15_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1640_LC_15_15_6  (
            .in0(N__41647),
            .in1(N__44607),
            .in2(N__36257),
            .in3(N__36530),
            .lcout(\c0.n22248 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1711_LC_15_15_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1711_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1711_LC_15_15_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1711_LC_15_15_7  (
            .in0(N__39288),
            .in1(N__36499),
            .in2(N__39392),
            .in3(N__39403),
            .lcout(\c0.n13338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i182_LC_15_16_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i182_LC_15_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i182_LC_15_16_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i182_LC_15_16_1  (
            .in0(N__59168),
            .in1(N__67201),
            .in2(_gnd_net_),
            .in3(N__63455),
            .lcout(data_in_frame_22_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66701),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1701_LC_15_16_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1701_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1701_LC_15_16_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_1701_LC_15_16_2  (
            .in0(N__36196),
            .in1(N__36299),
            .in2(N__36425),
            .in3(N__36377),
            .lcout(\c0.n16_adj_4478 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i2_LC_15_16_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i2_LC_15_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i2_LC_15_16_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i2_LC_15_16_3  (
            .in0(N__36300),
            .in1(N__43217),
            .in2(_gnd_net_),
            .in3(N__36331),
            .lcout(data_in_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66701),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__5__5472_LC_15_16_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__5__5472_LC_15_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__5__5472_LC_15_16_4 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_6__5__5472_LC_15_16_4  (
            .in0(N__49570),
            .in1(N__48833),
            .in2(N__38245),
            .in3(N__36285),
            .lcout(data_out_frame_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66701),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i15_LC_15_16_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i15_LC_15_16_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i15_LC_15_16_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i15_LC_15_16_5  (
            .in0(N__42168),
            .in1(N__36271),
            .in2(_gnd_net_),
            .in3(N__36256),
            .lcout(encoder0_position_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66701),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i17_LC_15_16_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i17_LC_15_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i17_LC_15_16_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i17_LC_15_16_6  (
            .in0(N__36197),
            .in1(N__43218),
            .in2(_gnd_net_),
            .in3(N__40243),
            .lcout(data_in_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66701),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i24_LC_15_16_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i24_LC_15_16_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i24_LC_15_16_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \quad_counter0.count_i0_i24_LC_15_16_7  (
            .in0(N__36178),
            .in1(_gnd_net_),
            .in2(N__42221),
            .in3(N__39324),
            .lcout(encoder0_position_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66701),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i31_LC_15_17_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i31_LC_15_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i31_LC_15_17_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_in_0___i31_LC_15_17_0  (
            .in0(N__43243),
            .in1(_gnd_net_),
            .in2(N__65591),
            .in3(N__36985),
            .lcout(data_in_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66715),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i226_LC_15_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i226_LC_15_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i226_LC_15_17_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i226_LC_15_17_1  (
            .in0(N__64561),
            .in1(N__63853),
            .in2(N__49962),
            .in3(N__67672),
            .lcout(\c0.data_in_frame_28_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66715),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i29_LC_15_17_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i29_LC_15_17_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i29_LC_15_17_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i29_LC_15_17_2  (
            .in0(N__42167),
            .in1(N__37000),
            .in2(_gnd_net_),
            .in3(N__38221),
            .lcout(encoder0_position_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66715),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i32_LC_15_17_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i32_LC_15_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i32_LC_15_17_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i32_LC_15_17_3  (
            .in0(N__68974),
            .in1(N__43245),
            .in2(_gnd_net_),
            .in3(N__36643),
            .lcout(data_in_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66715),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i23_LC_15_17_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i23_LC_15_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i23_LC_15_17_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i23_LC_15_17_4  (
            .in0(N__43239),
            .in1(N__36986),
            .in2(_gnd_net_),
            .in3(N__36947),
            .lcout(data_in_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66715),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_17_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_17_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_17_5  (
            .in0(N__36928),
            .in1(N__36818),
            .in2(N__37222),
            .in3(N__39726),
            .lcout(\c0.n24183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i24_LC_15_17_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i24_LC_15_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i24_LC_15_17_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i24_LC_15_17_6  (
            .in0(N__36644),
            .in1(_gnd_net_),
            .in2(N__43265),
            .in3(N__36623),
            .lcout(data_in_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66715),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i27_LC_15_17_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i27_LC_15_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i27_LC_15_17_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i27_LC_15_17_7  (
            .in0(N__36586),
            .in1(N__43244),
            .in2(_gnd_net_),
            .in3(N__68377),
            .lcout(data_in_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66715),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_LC_15_18_0 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_LC_15_18_0 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_LC_15_18_0  (
            .in0(N__56934),
            .in1(N__57027),
            .in2(_gnd_net_),
            .in3(N__56836),
            .lcout(\c0.rx.n21783 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__1__5436_LC_15_18_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__1__5436_LC_15_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__1__5436_LC_15_18_1 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_frame_11__1__5436_LC_15_18_1  (
            .in0(N__37221),
            .in1(N__48741),
            .in2(N__37264),
            .in3(N__49427),
            .lcout(data_out_frame_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66729),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_3_lut_LC_15_18_2 .C_ON=1'b0;
    defparam \c0.i20_3_lut_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i20_3_lut_LC_15_18_2 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \c0.i20_3_lut_LC_15_18_2  (
            .in0(N__49425),
            .in1(N__39138),
            .in2(_gnd_net_),
            .in3(N__40150),
            .lcout(),
            .ltout(\c0.n9_adj_4415_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1748_LC_15_18_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1748_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1748_LC_15_18_3 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \c0.i2_3_lut_adj_1748_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__40734),
            .in2(N__37207),
            .in3(N__40775),
            .lcout(n14252),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20381_3_lut_LC_15_18_5 .C_ON=1'b0;
    defparam \c0.i20381_3_lut_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20381_3_lut_LC_15_18_5 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \c0.i20381_3_lut_LC_15_18_5  (
            .in0(N__37170),
            .in1(_gnd_net_),
            .in2(N__37146),
            .in3(N__39248),
            .lcout(\c0.n23965 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1494_LC_15_18_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1494_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1494_LC_15_18_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_1494_LC_15_18_6  (
            .in0(N__37111),
            .in1(N__40149),
            .in2(N__40744),
            .in3(N__37360),
            .lcout(n22661),
            .ltout(n22661_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__3__5466_LC_15_18_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__3__5466_LC_15_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__3__5466_LC_15_18_7 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \c0.data_out_frame_7__3__5466_LC_15_18_7  (
            .in0(N__37098),
            .in1(N__49426),
            .in2(N__37105),
            .in3(N__38666),
            .lcout(data_out_frame_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66729),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1263_2_lut_3_lut_LC_15_19_0 .C_ON=1'b0;
    defparam \c0.i1263_2_lut_3_lut_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1263_2_lut_3_lut_LC_15_19_0 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \c0.i1263_2_lut_3_lut_LC_15_19_0  (
            .in0(N__40445),
            .in1(N__40595),
            .in2(_gnd_net_),
            .in3(N__42705),
            .lcout(\c0.n3239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__1__5476_LC_15_19_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__1__5476_LC_15_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__1__5476_LC_15_19_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_6__1__5476_LC_15_19_1  (
            .in0(N__49443),
            .in1(N__48736),
            .in2(N__39902),
            .in3(N__37084),
            .lcout(data_out_frame_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66743),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__0__5453_LC_15_19_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__0__5453_LC_15_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__0__5453_LC_15_19_2 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_9__0__5453_LC_15_19_2  (
            .in0(N__48735),
            .in1(N__49444),
            .in2(N__37071),
            .in3(N__37014),
            .lcout(data_out_frame_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66743),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1234_LC_15_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1234_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1234_LC_15_19_3 .LUT_INIT=16'b1110110011111111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1234_LC_15_19_3  (
            .in0(N__42704),
            .in1(N__40446),
            .in2(N__42507),
            .in3(N__40113),
            .lcout(\c0.n12967 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1698_LC_15_19_4 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1698_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1698_LC_15_19_4 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \c0.i1_3_lut_adj_1698_LC_15_19_4  (
            .in0(N__37297),
            .in1(N__37940),
            .in2(_gnd_net_),
            .in3(N__42703),
            .lcout(\c0.n12996 ),
            .ltout(\c0.n12996_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_15_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_15_19_5 .LUT_INIT=16'b1111100011111111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_LC_15_19_5  (
            .in0(N__42706),
            .in1(N__42502),
            .in2(N__37288),
            .in3(N__40114),
            .lcout(\c0.n13020 ),
            .ltout(\c0.n13020_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1677_LC_15_19_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1677_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1677_LC_15_19_6 .LUT_INIT=16'b1111011111110101;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1677_LC_15_19_6  (
            .in0(N__40447),
            .in1(N__40596),
            .in2(N__37285),
            .in3(N__42707),
            .lcout(\c0.n13021 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i0_LC_15_19_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i0_LC_15_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i0_LC_15_19_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i0_LC_15_19_7  (
            .in0(N__50107),
            .in1(N__69375),
            .in2(N__59690),
            .in3(N__59940),
            .lcout(rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66743),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_LC_15_20_0 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_LC_15_20_0 .LUT_INIT=16'b1011001100110011;
    LogicCell40 \c0.i1_3_lut_4_lut_LC_15_20_0  (
            .in0(N__37473),
            .in1(N__37428),
            .in2(N__37519),
            .in3(N__40402),
            .lcout(\c0.data_out_frame_29_7_N_1483_1 ),
            .ltout(\c0.data_out_frame_29_7_N_1483_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1678_LC_15_20_1 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1678_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1678_LC_15_20_1 .LUT_INIT=16'b1010111100001111;
    LogicCell40 \c0.i1_3_lut_adj_1678_LC_15_20_1  (
            .in0(N__37430),
            .in1(_gnd_net_),
            .in2(N__37282),
            .in3(N__37279),
            .lcout(\c0.n4_adj_4419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i157_4_lut_LC_15_20_2 .C_ON=1'b0;
    defparam \c0.i157_4_lut_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i157_4_lut_LC_15_20_2 .LUT_INIT=16'b1111110101010101;
    LogicCell40 \c0.i157_4_lut_LC_15_20_2  (
            .in0(N__37472),
            .in1(N__42498),
            .in2(N__37390),
            .in3(N__37514),
            .lcout(\c0.n6650 ),
            .ltout(\c0.n6650_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1331_LC_15_20_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1331_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1331_LC_15_20_3 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i1_4_lut_adj_1331_LC_15_20_3  (
            .in0(N__37429),
            .in1(N__37270),
            .in2(N__37273),
            .in3(N__37356),
            .lcout(\c0.n31_adj_4271 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1783_LC_15_20_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1783_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1783_LC_15_20_4 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_adj_1783_LC_15_20_4  (
            .in0(N__37471),
            .in1(N__40401),
            .in2(N__37944),
            .in3(N__37513),
            .lcout(\c0.n6_adj_4270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1696_LC_15_20_5 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1696_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1696_LC_15_20_5 .LUT_INIT=16'b1000100011111111;
    LogicCell40 \c0.i1_3_lut_adj_1696_LC_15_20_5  (
            .in0(N__37515),
            .in1(N__37388),
            .in2(_gnd_net_),
            .in3(N__37474),
            .lcout(),
            .ltout(\c0.n16958_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1491_LC_15_20_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1491_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1491_LC_15_20_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \c0.i2_3_lut_adj_1491_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__37345),
            .in2(N__37435),
            .in3(N__37431),
            .lcout(),
            .ltout(\c0.n22695_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i2_LC_15_20_7 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i2_LC_15_20_7 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i2_LC_15_20_7 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \c0.FRAME_MATCHER_state_i2_LC_15_20_7  (
            .in0(N__42568),
            .in1(N__42589),
            .in2(N__37393),
            .in3(N__40090),
            .lcout(\c0.FRAME_MATCHER_state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66757),
            .ce(),
            .sr(N__40934));
    defparam \c0.i14419_2_lut_4_lut_LC_15_21_1 .C_ON=1'b0;
    defparam \c0.i14419_2_lut_4_lut_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14419_2_lut_4_lut_LC_15_21_1 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.i14419_2_lut_4_lut_LC_15_21_1  (
            .in0(N__37818),
            .in1(N__37621),
            .in2(N__37372),
            .in3(N__42708),
            .lcout(\c0.n9207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1658_LC_15_21_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1658_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1658_LC_15_21_3 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1658_LC_15_21_3  (
            .in0(N__40575),
            .in1(N__40527),
            .in2(_gnd_net_),
            .in3(N__42709),
            .lcout(\c0.n12990 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1490_LC_15_21_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1490_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1490_LC_15_21_4 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \c0.i1_4_lut_adj_1490_LC_15_21_4  (
            .in0(N__42954),
            .in1(N__40419),
            .in2(N__42433),
            .in3(N__43340),
            .lcout(\c0.n14_adj_4337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1671_LC_15_21_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1671_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1671_LC_15_21_5 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1671_LC_15_21_5  (
            .in0(N__40745),
            .in1(N__40702),
            .in2(_gnd_net_),
            .in3(N__42710),
            .lcout(),
            .ltout(\c0.n7_adj_4352_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1533_LC_15_21_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1533_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1533_LC_15_21_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.i4_4_lut_adj_1533_LC_15_21_6  (
            .in0(N__54093),
            .in1(N__43341),
            .in2(N__37339),
            .in3(N__43291),
            .lcout(\c0.n6_adj_4353 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_adj_1637_LC_15_22_0 .C_ON=1'b0;
    defparam \c0.i20_4_lut_adj_1637_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_adj_1637_LC_15_22_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i20_4_lut_adj_1637_LC_15_22_0  (
            .in0(N__38109),
            .in1(N__42937),
            .in2(N__52663),
            .in3(N__37336),
            .lcout(),
            .ltout(\c0.n48_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i26_4_lut_LC_15_22_1 .C_ON=1'b0;
    defparam \c0.i26_4_lut_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i26_4_lut_LC_15_22_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i26_4_lut_LC_15_22_1  (
            .in0(N__37525),
            .in1(N__37762),
            .in2(N__37663),
            .in3(N__37660),
            .lcout(\c0.n54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1639_LC_15_22_4 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1639_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1639_LC_15_22_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i17_4_lut_adj_1639_LC_15_22_4  (
            .in0(N__37604),
            .in1(N__37653),
            .in2(N__41104),
            .in3(N__43540),
            .lcout(\c0.n45_adj_4413 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1434_LC_15_22_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1434_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1434_LC_15_22_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_1434_LC_15_22_5  (
            .in0(N__43503),
            .in1(N__52659),
            .in2(N__37654),
            .in3(N__37603),
            .lcout(\c0.n14_adj_4316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i24_LC_15_22_6 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i24_LC_15_22_6 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i24_LC_15_22_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i24_LC_15_22_6  (
            .in0(N__37605),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52815),
            .lcout(\c0.FRAME_MATCHER_state_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66784),
            .ce(),
            .sr(N__37588));
    defparam \c0.i14273_2_lut_LC_15_23_0 .C_ON=1'b0;
    defparam \c0.i14273_2_lut_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14273_2_lut_LC_15_23_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i14273_2_lut_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__40599),
            .in2(_gnd_net_),
            .in3(N__42768),
            .lcout(\c0.data_out_frame_29_7_N_1483_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1781_LC_15_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1781_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1781_LC_15_23_1 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1781_LC_15_23_1  (
            .in0(N__42769),
            .in1(N__37686),
            .in2(N__53168),
            .in3(N__42546),
            .lcout(\c0.n21342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1752_LC_15_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1752_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1752_LC_15_23_2 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1752_LC_15_23_2  (
            .in0(N__52970),
            .in1(_gnd_net_),
            .in2(N__37555),
            .in3(N__53116),
            .lcout(\c0.n21346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1766_LC_15_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1766_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1766_LC_15_23_3 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1766_LC_15_23_3  (
            .in0(N__53115),
            .in1(_gnd_net_),
            .in2(N__37918),
            .in3(N__52971),
            .lcout(\c0.n21364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_LC_15_23_5 .C_ON=1'b0;
    defparam \c0.i18_4_lut_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_LC_15_23_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i18_4_lut_LC_15_23_5  (
            .in0(N__43504),
            .in1(N__37852),
            .in2(N__42508),
            .in3(N__37551),
            .lcout(\c0.n46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1704_LC_15_23_6 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1704_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1704_LC_15_23_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i9_4_lut_adj_1704_LC_15_23_6  (
            .in0(N__37685),
            .in1(N__38108),
            .in2(N__43456),
            .in3(N__41100),
            .lcout(),
            .ltout(\c0.n21_adj_4480_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_adj_1716_LC_15_23_7 .C_ON=1'b0;
    defparam \c0.i11_3_lut_adj_1716_LC_15_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_adj_1716_LC_15_23_7 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \c0.i11_3_lut_adj_1716_LC_15_23_7  (
            .in0(_gnd_net_),
            .in1(N__37969),
            .in2(N__37957),
            .in3(N__37954),
            .lcout(\c0.n14789 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1871_LC_15_24_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1871_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1871_LC_15_24_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_1871_LC_15_24_1  (
            .in0(N__37913),
            .in1(N__41041),
            .in2(N__37885),
            .in3(N__37848),
            .lcout(\c0.n21682 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_1638_LC_15_24_2 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_1638_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_1638_LC_15_24_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i19_4_lut_adj_1638_LC_15_24_2  (
            .in0(N__37714),
            .in1(N__37687),
            .in2(N__43410),
            .in3(N__37804),
            .lcout(\c0.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1775_LC_15_24_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1775_LC_15_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1775_LC_15_24_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1775_LC_15_24_3  (
            .in0(N__37751),
            .in1(N__53136),
            .in2(_gnd_net_),
            .in3(N__52973),
            .lcout(\c0.n21374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1753_LC_15_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1753_LC_15_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1753_LC_15_24_5 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1753_LC_15_24_5  (
            .in0(N__53137),
            .in1(N__37715),
            .in2(_gnd_net_),
            .in3(N__52972),
            .lcout(\c0.n21348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i10_LC_15_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i10_LC_15_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i10_LC_15_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i10_LC_15_25_0  (
            .in0(_gnd_net_),
            .in1(N__37717),
            .in2(_gnd_net_),
            .in3(N__52859),
            .lcout(\c0.FRAME_MATCHER_state_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66816),
            .ce(),
            .sr(N__37693));
    defparam \c0.FRAME_MATCHER_state_i7_LC_15_26_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i7_LC_15_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i7_LC_15_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i7_LC_15_26_0  (
            .in0(_gnd_net_),
            .in1(N__37684),
            .in2(_gnd_net_),
            .in3(N__52884),
            .lcout(\c0.FRAME_MATCHER_state_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66828),
            .ce(),
            .sr(N__38119));
    defparam \c0.i1_2_lut_3_lut_adj_1755_LC_15_27_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1755_LC_15_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1755_LC_15_27_5 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1755_LC_15_27_5  (
            .in0(N__38110),
            .in1(N__53010),
            .in2(_gnd_net_),
            .in3(N__53176),
            .lcout(\c0.n21350 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i11_LC_15_29_4 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i11_LC_15_29_4 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i11_LC_15_29_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i11_LC_15_29_4  (
            .in0(_gnd_net_),
            .in1(N__38107),
            .in2(_gnd_net_),
            .in3(N__52888),
            .lcout(\c0.FRAME_MATCHER_state_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66859),
            .ce(),
            .sr(N__38083));
    defparam \c0.i14074_2_lut_3_lut_LC_16_8_0 .C_ON=1'b0;
    defparam \c0.i14074_2_lut_3_lut_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14074_2_lut_3_lut_LC_16_8_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i14074_2_lut_3_lut_LC_16_8_0  (
            .in0(N__56699),
            .in1(N__56573),
            .in2(_gnd_net_),
            .in3(N__56434),
            .lcout(\c0.n17596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__5__5424_LC_16_8_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__5__5424_LC_16_8_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__5__5424_LC_16_8_4 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_12__5__5424_LC_16_8_4  (
            .in0(N__49144),
            .in1(N__49048),
            .in2(N__38071),
            .in3(N__38007),
            .lcout(data_out_frame_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66634),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1648_LC_16_9_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1648_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1648_LC_16_9_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1648_LC_16_9_0  (
            .in0(N__56589),
            .in1(N__56435),
            .in2(_gnd_net_),
            .in3(N__46030),
            .lcout(\c0.n4_adj_4373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1626_LC_16_10_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1626_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1626_LC_16_10_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1626_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__47908),
            .in2(_gnd_net_),
            .in3(N__47956),
            .lcout(\c0.n20875 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1545_LC_16_10_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1545_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1545_LC_16_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i5_4_lut_adj_1545_LC_16_10_1  (
            .in0(N__51777),
            .in1(N__43870),
            .in2(N__48171),
            .in3(N__43919),
            .lcout(\c0.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1544_LC_16_10_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1544_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1544_LC_16_10_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_1544_LC_16_10_2  (
            .in0(N__50345),
            .in1(N__51778),
            .in2(N__47522),
            .in3(N__51711),
            .lcout(\c0.n14_adj_4365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1546_LC_16_10_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1546_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1546_LC_16_10_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i5_4_lut_adj_1546_LC_16_10_3  (
            .in0(N__43871),
            .in1(N__44167),
            .in2(N__48172),
            .in3(N__43920),
            .lcout(),
            .ltout(\c0.n13_adj_4366_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14078_4_lut_LC_16_10_4 .C_ON=1'b0;
    defparam \c0.i14078_4_lut_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14078_4_lut_LC_16_10_4 .LUT_INIT=16'b0111011101110000;
    LogicCell40 \c0.i14078_4_lut_LC_16_10_4  (
            .in0(N__37993),
            .in1(N__37984),
            .in2(N__37978),
            .in3(N__37975),
            .lcout(\c0.n17600 ),
            .ltout(\c0.n17600_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1624_LC_16_10_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1624_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1624_LC_16_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_1624_LC_16_10_5  (
            .in0(N__47266),
            .in1(N__38137),
            .in2(N__38131),
            .in3(N__54832),
            .lcout(\c0.n23648 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i6_LC_16_11_4 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i6_LC_16_11_4 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i6_LC_16_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i6_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__41083),
            .in2(_gnd_net_),
            .in3(N__52886),
            .lcout(\c0.FRAME_MATCHER_state_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66643),
            .ce(),
            .sr(N__41065));
    defparam \c0.i8_4_lut_adj_1629_LC_16_11_5 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1629_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1629_LC_16_11_5 .LUT_INIT=16'b1101111111111101;
    LogicCell40 \c0.i8_4_lut_adj_1629_LC_16_11_5  (
            .in0(N__54767),
            .in1(N__41215),
            .in2(N__44257),
            .in3(N__43990),
            .lcout(\c0.n18_adj_4403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1306_LC_16_11_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1306_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1306_LC_16_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1306_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(N__52391),
            .in2(_gnd_net_),
            .in3(N__54766),
            .lcout(\c0.n21825 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1307_LC_16_12_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1307_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1307_LC_16_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1307_LC_16_12_0  (
            .in0(N__38127),
            .in1(N__47930),
            .in2(N__48317),
            .in3(N__48255),
            .lcout(\c0.n13677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i85_LC_16_12_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i85_LC_16_12_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i85_LC_16_12_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i85_LC_16_12_1  (
            .in0(N__62493),
            .in1(N__69211),
            .in2(N__63217),
            .in3(N__38128),
            .lcout(\c0.data_in_frame_10_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66650),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i67_LC_16_12_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i67_LC_16_12_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i67_LC_16_12_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i67_LC_16_12_2  (
            .in0(N__65970),
            .in1(N__62494),
            .in2(N__47937),
            .in3(N__68416),
            .lcout(\c0.data_in_frame_8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66650),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i68_LC_16_12_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i68_LC_16_12_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i68_LC_16_12_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i68_LC_16_12_3  (
            .in0(N__62491),
            .in1(N__65972),
            .in2(N__48321),
            .in3(N__64851),
            .lcout(\c0.data_in_frame_8_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66650),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1665_LC_16_12_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1665_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1665_LC_16_12_4 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1665_LC_16_12_4  (
            .in0(N__56601),
            .in1(N__56456),
            .in2(N__56742),
            .in3(N__68097),
            .lcout(n21760),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i69_LC_16_12_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i69_LC_16_12_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i69_LC_16_12_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i69_LC_16_12_5  (
            .in0(N__62492),
            .in1(N__65973),
            .in2(N__63216),
            .in3(N__47450),
            .lcout(\c0.data_in_frame_8_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66650),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i78_LC_16_12_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i78_LC_16_12_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i78_LC_16_12_6 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i78_LC_16_12_6  (
            .in0(N__67215),
            .in1(N__62495),
            .in2(N__69876),
            .in3(N__47823),
            .lcout(\c0.data_in_frame_9_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66650),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i66_LC_16_12_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i66_LC_16_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i66_LC_16_12_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i66_LC_16_12_7  (
            .in0(N__62490),
            .in1(N__65971),
            .in2(N__52407),
            .in3(N__63865),
            .lcout(\c0.data_in_frame_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66650),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1475_LC_16_13_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1475_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1475_LC_16_13_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1475_LC_16_13_0  (
            .in0(N__40058),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39898),
            .lcout(\c0.n21908 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i20_LC_16_13_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i20_LC_16_13_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i20_LC_16_13_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i20_LC_16_13_1  (
            .in0(N__38504),
            .in1(N__38311),
            .in2(_gnd_net_),
            .in3(N__38914),
            .lcout(encoder1_position_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66658),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1419_LC_16_13_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1419_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1419_LC_16_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1419_LC_16_13_2  (
            .in0(N__41601),
            .in1(N__41869),
            .in2(N__38887),
            .in3(N__39101),
            .lcout(\c0.n13839 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1468_LC_16_13_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1468_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1468_LC_16_13_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1468_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(N__48562),
            .in2(_gnd_net_),
            .in3(N__38772),
            .lcout(\c0.n22015 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.encoder0_position_29__I_0_2_lut_LC_16_13_5 .C_ON=1'b0;
    defparam \c0.encoder0_position_29__I_0_2_lut_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.encoder0_position_29__I_0_2_lut_LC_16_13_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.encoder0_position_29__I_0_2_lut_LC_16_13_5  (
            .in0(N__38773),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38244),
            .lcout(\c0.data_out_frame_29__7__N_856 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1416_LC_16_13_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1416_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1416_LC_16_13_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1416_LC_16_13_6  (
            .in0(N__38163),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38610),
            .lcout(\c0.n6_adj_4311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1481_LC_16_13_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1481_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1481_LC_16_13_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1481_LC_16_13_7  (
            .in0(N__38986),
            .in1(N__38556),
            .in2(N__38611),
            .in3(N__38809),
            .lcout(\c0.n22427 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1843_LC_16_14_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1843_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1843_LC_16_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1843_LC_16_14_0  (
            .in0(N__39476),
            .in1(N__41862),
            .in2(N__38668),
            .in3(N__41800),
            .lcout(\c0.n21885 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_1177_LC_16_14_1 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_1177_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_1177_LC_16_14_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i1_2_lut_adj_1177_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(N__59884),
            .in2(_gnd_net_),
            .in3(N__57109),
            .lcout(n18678),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1473_LC_16_14_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1473_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1473_LC_16_14_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1473_LC_16_14_2  (
            .in0(N__42034),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42395),
            .lcout(\c0.n22200 ),
            .ltout(\c0.n22200_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1848_LC_16_14_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1848_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1848_LC_16_14_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1848_LC_16_14_3  (
            .in0(N__40208),
            .in1(N__39477),
            .in2(N__38593),
            .in3(N__38579),
            .lcout(\c0.n13705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1908_LC_16_14_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1908_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1908_LC_16_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1908_LC_16_14_4  (
            .in0(N__48450),
            .in1(N__47454),
            .in2(_gnd_net_),
            .in3(N__47254),
            .lcout(\c0.n13190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i12_LC_16_15_0 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i12_LC_16_15_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i12_LC_16_15_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i12_LC_16_15_0  (
            .in0(N__42235),
            .in1(N__38545),
            .in2(_gnd_net_),
            .in3(N__38859),
            .lcout(encoder0_position_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66671),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i4_LC_16_15_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i4_LC_16_15_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i4_LC_16_15_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i4_LC_16_15_1  (
            .in0(N__39016),
            .in1(N__42237),
            .in2(_gnd_net_),
            .in3(N__38536),
            .lcout(encoder0_position_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66671),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i10_LC_16_15_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i10_LC_16_15_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i10_LC_16_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i10_LC_16_15_2  (
            .in0(N__42234),
            .in1(N__38524),
            .in2(_gnd_net_),
            .in3(N__39974),
            .lcout(encoder0_position_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66671),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i16_LC_16_15_3 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i16_LC_16_15_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i16_LC_16_15_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i16_LC_16_15_3  (
            .in0(N__39090),
            .in1(N__42236),
            .in2(_gnd_net_),
            .in3(N__39127),
            .lcout(encoder0_position_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66671),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1474_LC_16_15_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1474_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1474_LC_16_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1474_LC_16_15_4  (
            .in0(N__41722),
            .in1(N__39089),
            .in2(_gnd_net_),
            .in3(N__39475),
            .lcout(\c0.n22128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1460_LC_16_15_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1460_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1460_LC_16_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1460_LC_16_15_5  (
            .in0(N__38916),
            .in1(N__53465),
            .in2(_gnd_net_),
            .in3(N__48558),
            .lcout(),
            .ltout(\c0.n22227_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1461_LC_16_15_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1461_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1461_LC_16_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1461_LC_16_15_6  (
            .in0(N__39064),
            .in1(N__39015),
            .in2(N__38989),
            .in3(N__38985),
            .lcout(\c0.n10444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1700_LC_16_15_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1700_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1700_LC_16_15_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1700_LC_16_15_7  (
            .in0(N__38915),
            .in1(N__48557),
            .in2(N__44618),
            .in3(N__53464),
            .lcout(\c0.n6_adj_4312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1478_LC_16_16_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1478_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1478_LC_16_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1478_LC_16_16_0  (
            .in0(N__38714),
            .in1(N__38847),
            .in2(_gnd_net_),
            .in3(N__39340),
            .lcout(\c0.n22477 ),
            .ltout(\c0.n22477_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1480_LC_16_16_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1480_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1480_LC_16_16_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1480_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38812),
            .in3(N__40257),
            .lcout(\c0.n6_adj_4333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i28_LC_16_16_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i28_LC_16_16_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i28_LC_16_16_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter0.count_i0_i28_LC_16_16_2  (
            .in0(N__38800),
            .in1(N__42233),
            .in2(_gnd_net_),
            .in3(N__38771),
            .lcout(encoder0_position_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66682),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1432_LC_16_16_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1432_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1432_LC_16_16_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1432_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(N__38715),
            .in2(_gnd_net_),
            .in3(N__40368),
            .lcout(),
            .ltout(\c0.n6_adj_4315_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1433_LC_16_16_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1433_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1433_LC_16_16_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1433_LC_16_16_4  (
            .in0(N__39318),
            .in1(N__40209),
            .in2(N__39433),
            .in3(N__42338),
            .lcout(\c0.n20171 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1687_LC_16_16_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1687_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1687_LC_16_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1687_LC_16_16_5  (
            .in0(N__42337),
            .in1(N__40040),
            .in2(_gnd_net_),
            .in3(N__39893),
            .lcout(\c0.data_out_frame_29__7__N_847 ),
            .ltout(\c0.data_out_frame_29__7__N_847_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1477_LC_16_16_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1477_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1477_LC_16_16_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1477_LC_16_16_6  (
            .in0(N__39317),
            .in1(N__39966),
            .in2(N__39397),
            .in3(N__39360),
            .lcout(\c0.n10_adj_4332 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1425_LC_16_16_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1425_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1425_LC_16_16_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1425_LC_16_16_7  (
            .in0(N__39967),
            .in1(N__39319),
            .in2(N__42306),
            .in3(N__39894),
            .lcout(\c0.n21931 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_transmit_5282_LC_16_17_0 .C_ON=1'b0;
    defparam \c0.tx_transmit_5282_LC_16_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx_transmit_5282_LC_16_17_0 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \c0.tx_transmit_5282_LC_16_17_0  (
            .in0(N__40158),
            .in1(N__39166),
            .in2(N__40750),
            .in3(N__49203),
            .lcout(\c0.r_SM_Main_2_N_3755_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66697),
            .ce(),
            .sr(N__40777));
    defparam \c0.i2_3_lut_adj_1649_LC_16_17_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1649_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1649_LC_16_17_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.i2_3_lut_adj_1649_LC_16_17_2  (
            .in0(N__40776),
            .in1(N__40081),
            .in2(_gnd_net_),
            .in3(N__40455),
            .lcout(\c0.n14322 ),
            .ltout(\c0.n14322_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11334_2_lut_3_lut_LC_16_17_3 .C_ON=1'b0;
    defparam \c0.i11334_2_lut_3_lut_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11334_2_lut_3_lut_LC_16_17_3 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \c0.i11334_2_lut_3_lut_LC_16_17_3  (
            .in0(N__40600),
            .in1(_gnd_net_),
            .in2(N__39205),
            .in3(N__42799),
            .lcout(\c0.n14871 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20360_4_lut_LC_16_17_5 .C_ON=1'b0;
    defparam \c0.i20360_4_lut_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20360_4_lut_LC_16_17_5 .LUT_INIT=16'b1000000010100010;
    LogicCell40 \c0.i20360_4_lut_LC_16_17_5  (
            .in0(N__40456),
            .in1(N__51367),
            .in2(N__39190),
            .in3(N__39139),
            .lcout(\c0.n23975 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1631_LC_16_17_6 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1631_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1631_LC_16_17_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i9_4_lut_adj_1631_LC_16_17_6  (
            .in0(N__47563),
            .in1(N__39160),
            .in2(N__52246),
            .in3(N__39148),
            .lcout(\c0.n17602 ),
            .ltout(\c0.n17602_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_3_lut_4_lut_LC_16_17_7 .C_ON=1'b0;
    defparam \c0.i14_3_lut_4_lut_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i14_3_lut_4_lut_LC_16_17_7 .LUT_INIT=16'b1100111100100010;
    LogicCell40 \c0.i14_3_lut_4_lut_LC_16_17_7  (
            .in0(N__49202),
            .in1(N__51366),
            .in2(N__40084),
            .in3(N__40157),
            .lcout(\c0.n8_adj_4417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__6__5463_LC_16_18_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__6__5463_LC_16_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__6__5463_LC_16_18_0 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_7__6__5463_LC_16_18_0  (
            .in0(N__49320),
            .in1(N__48734),
            .in2(N__42041),
            .in3(N__39847),
            .lcout(data_out_frame_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66710),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i26_LC_16_18_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i26_LC_16_18_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i26_LC_16_18_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i26_LC_16_18_1  (
            .in0(N__40039),
            .in1(N__42151),
            .in2(_gnd_net_),
            .in3(N__40075),
            .lcout(encoder0_position_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66710),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i8_LC_16_18_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i8_LC_16_18_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i8_LC_16_18_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \quad_counter0.count_i0_i8_LC_16_18_2  (
            .in0(N__39994),
            .in1(_gnd_net_),
            .in2(N__42203),
            .in3(N__40284),
            .lcout(encoder0_position_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__2__5459_LC_16_18_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__2__5459_LC_16_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__2__5459_LC_16_18_3 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_8__2__5459_LC_16_18_3  (
            .in0(N__48733),
            .in1(N__49321),
            .in2(N__39979),
            .in3(N__39933),
            .lcout(data_out_frame_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66710),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i25_LC_16_18_4 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i25_LC_16_18_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i25_LC_16_18_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i25_LC_16_18_4  (
            .in0(N__42150),
            .in1(N__39919),
            .in2(_gnd_net_),
            .in3(N__39889),
            .lcout(encoder0_position_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_16_18_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_16_18_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_16_18_5  (
            .in0(N__39846),
            .in1(N__48484),
            .in2(_gnd_net_),
            .in3(N__39832),
            .lcout(\c0.n5_adj_4350 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i2_LC_16_18_6 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i2_LC_16_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i2_LC_16_18_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i2_LC_16_18_6  (
            .in0(N__39486),
            .in1(N__52069),
            .in2(_gnd_net_),
            .in3(N__44661),
            .lcout(control_mode_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1686_LC_16_18_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1686_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1686_LC_16_18_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1686_LC_16_18_7  (
            .in0(N__42375),
            .in1(N__40359),
            .in2(N__40294),
            .in3(N__42286),
            .lcout(\c0.n22032 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i144_LC_16_19_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i144_LC_16_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i144_LC_16_19_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i144_LC_16_19_1  (
            .in0(N__69840),
            .in1(N__68096),
            .in2(N__57444),
            .in3(N__68972),
            .lcout(\c0.data_in_frame_17_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66725),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4649_2_lut_LC_16_19_3 .C_ON=1'b0;
    defparam \c0.i4649_2_lut_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4649_2_lut_LC_16_19_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.i4649_2_lut_LC_16_19_3  (
            .in0(N__48697),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49201),
            .lcout(\c0.n8107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i25_LC_16_19_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i25_LC_16_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i25_LC_16_19_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i25_LC_16_19_4  (
            .in0(N__69374),
            .in1(N__43215),
            .in2(_gnd_net_),
            .in3(N__40232),
            .lcout(data_in_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66725),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i197_LC_16_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i197_LC_16_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i197_LC_16_19_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i197_LC_16_19_5  (
            .in0(N__67622),
            .in1(N__65899),
            .in2(N__58938),
            .in3(N__63173),
            .lcout(\c0.data_in_frame_24_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66725),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i5_LC_16_19_6 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i5_LC_16_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i5_LC_16_19_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i5_LC_16_19_6  (
            .in0(N__40198),
            .in1(N__47644),
            .in2(_gnd_net_),
            .in3(N__44659),
            .lcout(control_mode_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66725),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_1532_LC_16_20_0 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_1532_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_1532_LC_16_20_0 .LUT_INIT=16'b1010001000000000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_1532_LC_16_20_0  (
            .in0(N__42744),
            .in1(N__42978),
            .in2(N__46174),
            .in3(N__40418),
            .lcout(\c0.n1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1684_LC_16_20_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1684_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1684_LC_16_20_1 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1684_LC_16_20_1  (
            .in0(N__40671),
            .in1(N__40624),
            .in2(N__40512),
            .in3(N__42610),
            .lcout(),
            .ltout(\c0.n23215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1492_LC_16_20_2 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1492_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1492_LC_16_20_2 .LUT_INIT=16'b0010111100100010;
    LogicCell40 \c0.i2_4_lut_adj_1492_LC_16_20_2  (
            .in0(N__42880),
            .in1(N__42835),
            .in2(N__40174),
            .in3(N__40159),
            .lcout(\c0.n6_adj_4338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18884_2_lut_LC_16_20_3 .C_ON=1'b0;
    defparam \c0.i18884_2_lut_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i18884_2_lut_LC_16_20_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.i18884_2_lut_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(N__48788),
            .in2(_gnd_net_),
            .in3(N__50780),
            .lcout(\c0.n22575 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_7_i3_2_lut_4_lut_LC_16_20_4 .C_ON=1'b0;
    defparam \c0.select_365_Select_7_i3_2_lut_4_lut_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_7_i3_2_lut_4_lut_LC_16_20_4 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \c0.select_365_Select_7_i3_2_lut_4_lut_LC_16_20_4  (
            .in0(N__50499),
            .in1(N__45178),
            .in2(N__50849),
            .in3(N__51371),
            .lcout(\c0.n3_adj_4465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1643_LC_16_20_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1643_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1643_LC_16_20_5 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1643_LC_16_20_5  (
            .in0(N__40576),
            .in1(N__42743),
            .in2(_gnd_net_),
            .in3(N__50498),
            .lcout(\c0.data_out_frame_0__7__N_2568 ),
            .ltout(\c0.data_out_frame_0__7__N_2568_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1893_LC_16_20_6 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1893_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1893_LC_16_20_6 .LUT_INIT=16'b1111000011110111;
    LogicCell40 \c0.i2_4_lut_adj_1893_LC_16_20_6  (
            .in0(N__40623),
            .in1(N__40505),
            .in2(N__40492),
            .in3(N__40670),
            .lcout(\c0.n1220 ),
            .ltout(\c0.n1220_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_11_i3_2_lut_4_lut_LC_16_20_7 .C_ON=1'b0;
    defparam \c0.select_365_Select_11_i3_2_lut_4_lut_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_11_i3_2_lut_4_lut_LC_16_20_7 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \c0.select_365_Select_11_i3_2_lut_4_lut_LC_16_20_7  (
            .in0(N__51372),
            .in1(N__45331),
            .in2(N__40489),
            .in3(N__50500),
            .lcout(\c0.n3_adj_4458 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14213_4_lut_LC_16_21_1 .C_ON=1'b0;
    defparam \c0.i14213_4_lut_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14213_4_lut_LC_16_21_1 .LUT_INIT=16'b0000111100001000;
    LogicCell40 \c0.i14213_4_lut_LC_16_21_1  (
            .in0(N__40486),
            .in1(N__45081),
            .in2(N__46175),
            .in3(N__44821),
            .lcout(\c0.n5024 ),
            .ltout(\c0.n5024_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1592_LC_16_21_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1592_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1592_LC_16_21_2 .LUT_INIT=16'b1111111100000011;
    LogicCell40 \c0.i1_3_lut_adj_1592_LC_16_21_2  (
            .in0(_gnd_net_),
            .in1(N__42584),
            .in2(N__40474),
            .in3(N__43279),
            .lcout(\c0.n21773 ),
            .ltout(\c0.n21773_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1458_LC_16_21_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1458_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1458_LC_16_21_3 .LUT_INIT=16'b1101010111000100;
    LogicCell40 \c0.i1_4_lut_adj_1458_LC_16_21_3  (
            .in0(N__42833),
            .in1(N__40453),
            .in2(N__40459),
            .in3(N__42884),
            .lcout(),
            .ltout(\c0.n4_adj_4328_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i1_LC_16_21_4 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i1_LC_16_21_4 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i1_LC_16_21_4 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \c0.FRAME_MATCHER_state_i1_LC_16_21_4  (
            .in0(N__40454),
            .in1(N__42955),
            .in2(N__40423),
            .in3(N__40420),
            .lcout(\c0.FRAME_MATCHER_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66752),
            .ce(),
            .sr(N__40927));
    defparam \c0.FRAME_MATCHER_state_i0_LC_16_21_5 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i0_LC_16_21_5 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i0_LC_16_21_5 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \c0.FRAME_MATCHER_state_i0_LC_16_21_5  (
            .in0(N__51322),
            .in1(N__40393),
            .in2(N__40381),
            .in3(N__50537),
            .lcout(\c0.FRAME_MATCHER_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66752),
            .ce(),
            .sr(N__40927));
    defparam \c0.i18974_4_lut_LC_16_22_1 .C_ON=1'b0;
    defparam \c0.i18974_4_lut_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i18974_4_lut_LC_16_22_1 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \c0.i18974_4_lut_LC_16_22_1  (
            .in0(N__42793),
            .in1(N__40807),
            .in2(N__40798),
            .in3(N__40783),
            .lcout(\c0.n22665 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1656_LC_16_22_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1656_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1656_LC_16_22_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1656_LC_16_22_2  (
            .in0(N__40628),
            .in1(N__40535),
            .in2(N__40597),
            .in3(N__42789),
            .lcout(\c0.n63_adj_4293 ),
            .ltout(\c0.n63_adj_4293_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1670_LC_16_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1670_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1670_LC_16_22_3 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1670_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(N__40749),
            .in2(N__40705),
            .in3(N__40701),
            .lcout(\c0.n21734 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1528_LC_16_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1528_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1528_LC_16_22_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i1_2_lut_adj_1528_LC_16_22_4  (
            .in0(_gnd_net_),
            .in1(N__42611),
            .in2(_gnd_net_),
            .in3(N__42791),
            .lcout(),
            .ltout(\c0.n84_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1525_LC_16_22_5 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1525_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1525_LC_16_22_5 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \c0.i2_4_lut_adj_1525_LC_16_22_5  (
            .in0(N__43008),
            .in1(N__40687),
            .in2(N__40675),
            .in3(N__40672),
            .lcout(\c0.n7_adj_4344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1663_LC_16_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1663_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1663_LC_16_22_6 .LUT_INIT=16'b1110111111101110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1663_LC_16_22_6  (
            .in0(N__40629),
            .in1(N__40539),
            .in2(N__40598),
            .in3(N__42790),
            .lcout(\c0.n12992 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1660_LC_16_22_7 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1660_LC_16_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1660_LC_16_22_7 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_adj_1660_LC_16_22_7  (
            .in0(N__42792),
            .in1(N__40585),
            .in2(N__40540),
            .in3(N__40513),
            .lcout(\c0.n12991 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1644_LC_16_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1644_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1644_LC_16_23_0 .LUT_INIT=16'b1100110000001000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1644_LC_16_23_0  (
            .in0(N__42795),
            .in1(N__41146),
            .in2(N__42616),
            .in3(N__53128),
            .lcout(\c0.n8_adj_4396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i30_LC_16_23_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i30_LC_16_23_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i30_LC_16_23_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i30_LC_16_23_1  (
            .in0(N__41147),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52843),
            .lcout(\c0.FRAME_MATCHER_state_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66779),
            .ce(),
            .sr(N__41122));
    defparam \c0.i1_2_lut_4_lut_adj_1779_LC_16_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1779_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1779_LC_16_23_2 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1779_LC_16_23_2  (
            .in0(N__42796),
            .in1(N__41003),
            .in2(N__42545),
            .in3(N__53129),
            .lcout(\c0.n21338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1646_LC_16_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1646_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1646_LC_16_23_3 .LUT_INIT=16'b1011000010100000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1646_LC_16_23_3  (
            .in0(N__53130),
            .in1(N__42615),
            .in2(N__41052),
            .in3(N__42797),
            .lcout(\c0.n8_adj_4398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1683_LC_16_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1683_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1683_LC_16_23_5 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1683_LC_16_23_5  (
            .in0(N__42825),
            .in1(N__43007),
            .in2(N__42886),
            .in3(N__42794),
            .lcout(\c0.n21737 ),
            .ltout(\c0.n21737_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1780_LC_16_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1780_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1780_LC_16_23_6 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1780_LC_16_23_6  (
            .in0(N__42538),
            .in1(N__42798),
            .in2(N__41107),
            .in3(N__41099),
            .lcout(\c0.n21340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i19_LC_16_24_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i19_LC_16_24_3 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i19_LC_16_24_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i19_LC_16_24_3  (
            .in0(_gnd_net_),
            .in1(N__41048),
            .in2(_gnd_net_),
            .in3(N__52845),
            .lcout(\c0.FRAME_MATCHER_state_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66791),
            .ce(),
            .sr(N__41020));
    defparam \c0.FRAME_MATCHER_state_i12_LC_16_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i12_LC_16_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i12_LC_16_25_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i12_LC_16_25_0  (
            .in0(N__52847),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42928),
            .lcout(\c0.FRAME_MATCHER_state_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66801),
            .ce(),
            .sr(N__42898));
    defparam \c0.FRAME_MATCHER_state_i5_LC_16_26_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i5_LC_16_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i5_LC_16_26_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i5_LC_16_26_0  (
            .in0(N__52848),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40996),
            .lcout(\c0.FRAME_MATCHER_state_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66811),
            .ce(),
            .sr(N__40966));
    defparam \c0.i1_2_lut_3_lut_adj_1760_LC_16_27_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1760_LC_16_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1760_LC_16_27_0 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1760_LC_16_27_0  (
            .in0(N__43393),
            .in1(N__53177),
            .in2(_gnd_net_),
            .in3(N__53022),
            .lcout(\c0.n21358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i132_LC_17_8_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i132_LC_17_8_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i132_LC_17_8_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i132_LC_17_8_0  (
            .in0(N__66013),
            .in1(N__68167),
            .in2(N__58130),
            .in3(N__64883),
            .lcout(\c0.data_in_frame_16_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66636),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20141_4_lut_LC_17_8_1 .C_ON=1'b0;
    defparam \c0.i20141_4_lut_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i20141_4_lut_LC_17_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i20141_4_lut_LC_17_8_1  (
            .in0(N__43921),
            .in1(N__50388),
            .in2(N__48168),
            .in3(N__43878),
            .lcout(\c0.n23836 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i4_LC_17_8_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i4_LC_17_8_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i4_LC_17_8_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i4_LC_17_8_2  (
            .in0(N__66014),
            .in1(N__60759),
            .in2(N__48153),
            .in3(N__64884),
            .lcout(\c0.data_in_frame_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66636),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1633_LC_17_8_3 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1633_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1633_LC_17_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i14_4_lut_adj_1633_LC_17_8_3  (
            .in0(N__43818),
            .in1(N__48046),
            .in2(N__52068),
            .in3(N__44698),
            .lcout(),
            .ltout(\c0.n38_adj_4407_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_LC_17_8_4 .C_ON=1'b0;
    defparam \c0.i19_4_lut_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_LC_17_8_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.i19_4_lut_LC_17_8_4  (
            .in0(N__41239),
            .in1(N__54420),
            .in2(N__41170),
            .in3(N__44166),
            .lcout(),
            .ltout(\c0.n43_adj_4410_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_4_lut_LC_17_8_5 .C_ON=1'b0;
    defparam \c0.i23_4_lut_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i23_4_lut_LC_17_8_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \c0.i23_4_lut_LC_17_8_5  (
            .in0(N__41197),
            .in1(N__41167),
            .in2(N__41161),
            .in3(N__43549),
            .lcout(FRAME_MATCHER_state_31_N_2976_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i65_LC_17_9_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i65_LC_17_9_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i65_LC_17_9_0 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i65_LC_17_9_0  (
            .in0(N__69555),
            .in1(N__62379),
            .in2(N__65991),
            .in3(N__51938),
            .lcout(\c0.data_in_frame_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66640),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1855_LC_17_9_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1855_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1855_LC_17_9_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1855_LC_17_9_1  (
            .in0(N__47906),
            .in1(N__51800),
            .in2(N__51942),
            .in3(N__51979),
            .lcout(\c0.n22443 ),
            .ltout(\c0.n22443_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1219_LC_17_9_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1219_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1219_LC_17_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1219_LC_17_9_2  (
            .in0(N__52546),
            .in1(N__51819),
            .in2(N__41158),
            .in3(N__47844),
            .lcout(\c0.n13287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1301_LC_17_9_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1301_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1301_LC_17_9_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1301_LC_17_9_3  (
            .in0(_gnd_net_),
            .in1(N__54747),
            .in2(_gnd_net_),
            .in3(N__54663),
            .lcout(\c0.n22283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1541_LC_17_9_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1541_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1541_LC_17_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1541_LC_17_9_4  (
            .in0(_gnd_net_),
            .in1(N__41178),
            .in2(_gnd_net_),
            .in3(N__44099),
            .lcout(\c0.n21986 ),
            .ltout(\c0.n21986_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1715_LC_17_9_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1715_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1715_LC_17_9_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1715_LC_17_9_5  (
            .in0(N__47623),
            .in1(N__48028),
            .in2(N__41182),
            .in3(N__47993),
            .lcout(\c0.n13180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3725_2_lut_LC_17_9_6 .C_ON=1'b0;
    defparam \c0.i3725_2_lut_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3725_2_lut_LC_17_9_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3725_2_lut_LC_17_9_6  (
            .in0(_gnd_net_),
            .in1(N__41278),
            .in2(_gnd_net_),
            .in3(N__53328),
            .lcout(\c0.n6404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i49_LC_17_9_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i49_LC_17_9_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i49_LC_17_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i49_LC_17_9_7  (
            .in0(N__41179),
            .in1(N__69556),
            .in2(_gnd_net_),
            .in3(N__49707),
            .lcout(data_in_frame_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66640),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i43_LC_17_10_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i43_LC_17_10_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i43_LC_17_10_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i43_LC_17_10_0  (
            .in0(N__62187),
            .in1(N__60766),
            .in2(N__43630),
            .in3(N__68354),
            .lcout(\c0.data_in_frame_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66647),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i29_LC_17_10_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i29_LC_17_10_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i29_LC_17_10_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i29_LC_17_10_1  (
            .in0(N__60761),
            .in1(N__63226),
            .in2(N__43609),
            .in3(N__67460),
            .lcout(\c0.data_in_frame_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66647),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1538_LC_17_10_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1538_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1538_LC_17_10_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1538_LC_17_10_2  (
            .in0(N__43591),
            .in1(N__43690),
            .in2(N__47788),
            .in3(N__43605),
            .lcout(\c0.n13237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i30_LC_17_10_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i30_LC_17_10_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i30_LC_17_10_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i30_LC_17_10_3  (
            .in0(N__60762),
            .in1(N__67458),
            .in2(N__67209),
            .in3(N__47997),
            .lcout(\c0.data_in_frame_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66647),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i11_LC_17_10_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i11_LC_17_10_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i11_LC_17_10_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i11_LC_17_10_4  (
            .in0(N__69844),
            .in1(N__60764),
            .in2(N__52058),
            .in3(N__68353),
            .lcout(data_in_frame_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66647),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i31_LC_17_10_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i31_LC_17_10_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i31_LC_17_10_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i31_LC_17_10_5  (
            .in0(N__60763),
            .in1(N__67459),
            .in2(N__44104),
            .in3(N__65582),
            .lcout(\c0.data_in_frame_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66647),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i12_LC_17_10_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i12_LC_17_10_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i12_LC_17_10_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i12_LC_17_10_6  (
            .in0(N__69845),
            .in1(N__60765),
            .in2(N__48047),
            .in3(N__64894),
            .lcout(data_in_frame_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66647),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i14_LC_17_10_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i14_LC_17_10_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i14_LC_17_10_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i14_LC_17_10_7  (
            .in0(N__60760),
            .in1(N__69846),
            .in2(N__67208),
            .in3(N__47631),
            .lcout(data_in_frame_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66647),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1668_LC_17_11_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1668_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1668_LC_17_11_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1668_LC_17_11_0  (
            .in0(N__47624),
            .in1(N__44297),
            .in2(N__43684),
            .in3(N__43810),
            .lcout(),
            .ltout(\c0.n6_adj_4393_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1601_LC_17_11_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1601_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1601_LC_17_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1601_LC_17_11_1  (
            .in0(N__41254),
            .in1(N__41208),
            .in2(N__41188),
            .in3(N__44079),
            .lcout(\c0.n13086 ),
            .ltout(\c0.n13086_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_LC_17_11_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_LC_17_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__47446),
            .in2(N__41185),
            .in3(N__47901),
            .lcout(\c0.n6_adj_4220 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1593_LC_17_11_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1593_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1593_LC_17_11_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1593_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(N__43724),
            .in2(_gnd_net_),
            .in3(N__43868),
            .lcout(\c0.n21893 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i18_LC_17_11_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i18_LC_17_11_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i18_LC_17_11_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i18_LC_17_11_4  (
            .in0(N__69231),
            .in1(N__63716),
            .in2(N__43729),
            .in3(N__60843),
            .lcout(\c0.data_in_frame_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66654),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i34_LC_17_11_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i34_LC_17_11_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i34_LC_17_11_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i34_LC_17_11_5  (
            .in0(N__60842),
            .in1(N__44080),
            .in2(N__64551),
            .in3(N__63864),
            .lcout(\c0.data_in_frame_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66654),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i1_LC_17_11_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i1_LC_17_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i1_LC_17_11_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i1_LC_17_11_6  (
            .in0(N__43869),
            .in1(N__69563),
            .in2(N__66012),
            .in3(N__60844),
            .lcout(\c0.data_in_frame_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66654),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1831_LC_17_11_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1831_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1831_LC_17_11_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1831_LC_17_11_7  (
            .in0(N__51801),
            .in1(N__51978),
            .in2(N__47907),
            .in3(N__47239),
            .lcout(\c0.n22280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i51_LC_17_12_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i51_LC_17_12_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i51_LC_17_12_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i51_LC_17_12_0  (
            .in0(N__68355),
            .in1(N__49691),
            .in2(_gnd_net_),
            .in3(N__43771),
            .lcout(data_in_frame_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66660),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i16_LC_17_12_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i16_LC_17_12_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i16_LC_17_12_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i16_LC_17_12_1  (
            .in0(N__69847),
            .in1(N__68958),
            .in2(N__44309),
            .in3(N__60835),
            .lcout(data_in_frame_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66660),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i15_LC_17_12_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i15_LC_17_12_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i15_LC_17_12_2 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i15_LC_17_12_2  (
            .in0(N__60834),
            .in1(N__65674),
            .in2(N__69794),
            .in3(N__43817),
            .lcout(data_in_frame_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66660),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1634_LC_17_12_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1634_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1634_LC_17_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_1634_LC_17_12_4  (
            .in0(N__47633),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43728),
            .lcout(\c0.n25_adj_4408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1625_LC_17_12_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1625_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1625_LC_17_12_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_1625_LC_17_12_5  (
            .in0(N__47802),
            .in1(N__50413),
            .in2(N__41227),
            .in3(N__47246),
            .lcout(\c0.n16_adj_4401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1602_LC_17_12_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1602_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1602_LC_17_12_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1602_LC_17_12_6  (
            .in0(N__41209),
            .in1(N__43735),
            .in2(N__41581),
            .in3(N__44298),
            .lcout(\c0.n13043 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i56_LC_17_12_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i56_LC_17_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i56_LC_17_12_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i56_LC_17_12_7  (
            .in0(N__49692),
            .in1(N__68957),
            .in2(_gnd_net_),
            .in3(N__44255),
            .lcout(data_in_frame_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66660),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_LC_17_13_0 .C_ON=1'b0;
    defparam \c0.i20_4_lut_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_LC_17_13_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.i20_4_lut_LC_17_13_0  (
            .in0(N__44263),
            .in1(N__48088),
            .in2(N__51649),
            .in3(N__44449),
            .lcout(\c0.n44_adj_4409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1587_LC_17_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1587_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1587_LC_17_13_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1587_LC_17_13_1  (
            .in0(N__44136),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43899),
            .lcout(\c0.n21791 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i37_LC_17_13_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i37_LC_17_13_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i37_LC_17_13_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i37_LC_17_13_2  (
            .in0(N__60849),
            .in1(N__64550),
            .in2(N__43756),
            .in3(N__63206),
            .lcout(\c0.data_in_frame_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i19_LC_17_13_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i19_LC_17_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i19_LC_17_13_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i19_LC_17_13_3  (
            .in0(N__69226),
            .in1(N__60850),
            .in2(N__44344),
            .in3(N__68426),
            .lcout(\c0.data_in_frame_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1575_LC_17_13_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1575_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1575_LC_17_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1575_LC_17_13_4  (
            .in0(N__43833),
            .in1(N__44197),
            .in2(N__44185),
            .in3(N__43752),
            .lcout(\c0.n21934 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i20_LC_17_13_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i20_LC_17_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i20_LC_17_13_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i20_LC_17_13_5  (
            .in0(N__69227),
            .in1(N__60851),
            .in2(N__44048),
            .in3(N__64824),
            .lcout(\c0.data_in_frame_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i2_LC_17_13_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i2_LC_17_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i2_LC_17_13_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i2_LC_17_13_6  (
            .in0(N__60848),
            .in1(N__43918),
            .in2(N__66015),
            .in3(N__63850),
            .lcout(\c0.data_in_frame_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i23_LC_17_13_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i23_LC_17_13_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i23_LC_17_13_7 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0__i23_LC_17_13_7  (
            .in0(N__50381),
            .in1(N__60852),
            .in2(N__69244),
            .in3(N__65673),
            .lcout(\c0.data_in_frame_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i167_LC_17_14_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i167_LC_17_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i167_LC_17_14_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i167_LC_17_14_0  (
            .in0(N__65672),
            .in1(N__68018),
            .in2(N__41277),
            .in3(N__64523),
            .lcout(\c0.data_in_frame_20_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1650_LC_17_14_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1650_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1650_LC_17_14_1 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1650_LC_17_14_1  (
            .in0(N__56605),
            .in1(N__56465),
            .in2(N__56748),
            .in3(N__60642),
            .lcout(n21744),
            .ltout(n21744_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i52_LC_17_14_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i52_LC_17_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i52_LC_17_14_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \c0.data_in_frame_0__i52_LC_17_14_2  (
            .in0(_gnd_net_),
            .in1(N__64826),
            .in2(N__41257),
            .in3(N__41253),
            .lcout(data_in_frame_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i168_LC_17_14_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i168_LC_17_14_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i168_LC_17_14_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i168_LC_17_14_3  (
            .in0(N__68017),
            .in1(N__64519),
            .in2(N__68973),
            .in3(N__53321),
            .lcout(\c0.data_in_frame_20_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i170_LC_17_14_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i170_LC_17_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i170_LC_17_14_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i170_LC_17_14_4  (
            .in0(N__62185),
            .in1(N__68019),
            .in2(N__53279),
            .in3(N__63855),
            .lcout(\c0.data_in_frame_21_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i42_LC_17_14_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i42_LC_17_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i42_LC_17_14_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i42_LC_17_14_5  (
            .in0(N__63854),
            .in1(N__60644),
            .in2(N__44383),
            .in3(N__62186),
            .lcout(\c0.data_in_frame_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i40_LC_17_14_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i40_LC_17_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i40_LC_17_14_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i40_LC_17_14_6  (
            .in0(N__60643),
            .in1(N__68940),
            .in2(N__64552),
            .in3(N__44401),
            .lcout(\c0.data_in_frame_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i63_LC_17_14_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i63_LC_17_14_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i63_LC_17_14_7 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \c0.data_in_frame_0__i63_LC_17_14_7  (
            .in0(N__54746),
            .in1(N__60645),
            .in2(N__68671),
            .in3(N__65671),
            .lcout(\c0.data_in_frame_7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66676),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i18_LC_17_15_0 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i18_LC_17_15_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i18_LC_17_15_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i18_LC_17_15_0  (
            .in0(N__42238),
            .in1(N__41305),
            .in2(_gnd_net_),
            .in3(N__41746),
            .lcout(encoder0_position_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66688),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1430_LC_17_15_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1430_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1430_LC_17_15_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1430_LC_17_15_2  (
            .in0(N__44606),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41744),
            .lcout(\c0.n21816 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_LC_17_15_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_LC_17_15_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_LC_17_15_4  (
            .in0(N__46048),
            .in1(N__47320),
            .in2(N__45077),
            .in3(N__44728),
            .lcout(\c0.n21740 ),
            .ltout(\c0.n21740_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i5_LC_17_15_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i5_LC_17_15_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i5_LC_17_15_5 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i5_LC_17_15_5  (
            .in0(N__65932),
            .in1(N__63170),
            .in2(N__41281),
            .in3(N__50321),
            .lcout(\c0.data_in_frame_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66688),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_12_i3_2_lut_4_lut_LC_17_15_6 .C_ON=1'b0;
    defparam \c0.select_365_Select_12_i3_2_lut_4_lut_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_12_i3_2_lut_4_lut_LC_17_15_6 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_12_i3_2_lut_4_lut_LC_17_15_6  (
            .in0(N__51470),
            .in1(N__51096),
            .in2(N__45384),
            .in3(N__50660),
            .lcout(\c0.n3_adj_4456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1459_LC_17_15_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1459_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1459_LC_17_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1459_LC_17_15_7  (
            .in0(N__41745),
            .in1(N__41700),
            .in2(_gnd_net_),
            .in3(N__41650),
            .lcout(\c0.n21813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_4_i3_2_lut_4_lut_LC_17_16_0 .C_ON=1'b0;
    defparam \c0.select_365_Select_4_i3_2_lut_4_lut_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_4_i3_2_lut_4_lut_LC_17_16_0 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_4_i3_2_lut_4_lut_LC_17_16_0  (
            .in0(N__51463),
            .in1(N__51011),
            .in2(N__45085),
            .in3(N__50664),
            .lcout(\c0.n3_adj_4470 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i54_LC_17_16_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i54_LC_17_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i54_LC_17_16_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i54_LC_17_16_1  (
            .in0(N__67161),
            .in1(N__49693),
            .in2(_gnd_net_),
            .in3(N__41577),
            .lcout(data_in_frame_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66702),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_14_i3_2_lut_4_lut_LC_17_16_2 .C_ON=1'b0;
    defparam \c0.select_365_Select_14_i3_2_lut_4_lut_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_14_i3_2_lut_4_lut_LC_17_16_2 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_14_i3_2_lut_4_lut_LC_17_16_2  (
            .in0(N__51464),
            .in1(N__51012),
            .in2(N__45439),
            .in3(N__50665),
            .lcout(\c0.n3_adj_4453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_8_i3_2_lut_4_lut_LC_17_16_3 .C_ON=1'b0;
    defparam \c0.select_365_Select_8_i3_2_lut_4_lut_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_8_i3_2_lut_4_lut_LC_17_16_3 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \c0.select_365_Select_8_i3_2_lut_4_lut_LC_17_16_3  (
            .in0(N__50666),
            .in1(N__45229),
            .in2(N__51089),
            .in3(N__51465),
            .lcout(\c0.n3_adj_4463 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i6_LC_17_16_5 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i6_LC_17_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i6_LC_17_16_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i6_LC_17_16_5  (
            .in0(N__41534),
            .in1(N__41492),
            .in2(_gnd_net_),
            .in3(N__41563),
            .lcout(\c0.tx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66702),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i8_LC_17_16_6 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i8_LC_17_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i8_LC_17_16_6 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.tx.r_Clock_Count__i8_LC_17_16_6  (
            .in0(N__41512),
            .in1(N__41327),
            .in2(N__41497),
            .in3(N__41386),
            .lcout(r_Clock_Count_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66702),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i21_LC_17_17_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i21_LC_17_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i21_LC_17_17_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i21_LC_17_17_0  (
            .in0(N__41889),
            .in1(N__43157),
            .in2(_gnd_net_),
            .in3(N__41992),
            .lcout(data_in_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66716),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i210_LC_17_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i210_LC_17_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i210_LC_17_17_1 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i210_LC_17_17_1  (
            .in0(N__63815),
            .in1(N__58766),
            .in2(N__69245),
            .in3(N__67610),
            .lcout(\c0.data_in_frame_26_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66716),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i22_LC_17_17_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i22_LC_17_17_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i22_LC_17_17_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter0.count_i0_i22_LC_17_17_2  (
            .in0(N__42265),
            .in1(N__42232),
            .in2(_gnd_net_),
            .in3(N__42030),
            .lcout(encoder0_position_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66716),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i13_LC_17_17_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i13_LC_17_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i13_LC_17_17_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i13_LC_17_17_3  (
            .in0(N__41993),
            .in1(N__43169),
            .in2(_gnd_net_),
            .in3(N__41950),
            .lcout(data_in_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66716),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14264_2_lut_3_lut_LC_17_17_4 .C_ON=1'b0;
    defparam \c0.i14264_2_lut_3_lut_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14264_2_lut_3_lut_LC_17_17_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.i14264_2_lut_3_lut_LC_17_17_4  (
            .in0(N__41923),
            .in1(N__43156),
            .in2(_gnd_net_),
            .in3(N__50929),
            .lcout(\c0.n17790 ),
            .ltout(\c0.n17790_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1895_LC_17_17_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1895_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1895_LC_17_17_5 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_adj_1895_LC_17_17_5  (
            .in0(N__45069),
            .in1(N__46054),
            .in2(N__41899),
            .in3(N__47323),
            .lcout(\c0.n21775 ),
            .ltout(\c0.n21775_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i218_LC_17_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i218_LC_17_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i218_LC_17_17_6 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0__i218_LC_17_17_6  (
            .in0(N__50191),
            .in1(N__67407),
            .in2(N__41896),
            .in3(N__63816),
            .lcout(\c0.data_in_frame_27_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66716),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i29_LC_17_17_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i29_LC_17_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i29_LC_17_17_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i29_LC_17_17_7  (
            .in0(N__63188),
            .in1(N__43170),
            .in2(_gnd_net_),
            .in3(N__41888),
            .lcout(data_in_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66716),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1562_LC_17_18_0 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1562_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1562_LC_17_18_0 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \c0.i2_4_lut_adj_1562_LC_17_18_0  (
            .in0(N__42638),
            .in1(N__56599),
            .in2(N__56749),
            .in3(N__56466),
            .lcout(\c0.n19783 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i1_LC_17_18_1 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i1_LC_17_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i1_LC_17_18_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i1_LC_17_18_1  (
            .in0(N__41843),
            .in1(N__47700),
            .in2(_gnd_net_),
            .in3(N__44654),
            .lcout(control_mode_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66730),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i3_LC_17_18_3 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i3_LC_17_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i3_LC_17_18_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i3_LC_17_18_3  (
            .in0(N__41784),
            .in1(N__48058),
            .in2(_gnd_net_),
            .in3(N__44655),
            .lcout(control_mode_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66730),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i183_LC_17_18_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i183_LC_17_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i183_LC_17_18_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i183_LC_17_18_5  (
            .in0(N__65698),
            .in1(N__62729),
            .in2(_gnd_net_),
            .in3(N__59200),
            .lcout(data_in_frame_22_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66730),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i4_LC_17_18_6 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i4_LC_17_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i4_LC_17_18_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.control_mode_i0_i4_LC_17_18_6  (
            .in0(N__54421),
            .in1(_gnd_net_),
            .in2(N__44662),
            .in3(N__42385),
            .lcout(control_mode_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66730),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i7_LC_17_19_1 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i7_LC_17_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i7_LC_17_19_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \c0.control_mode_i0_i7_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(N__42336),
            .in2(N__44320),
            .in3(N__44653),
            .lcout(control_mode_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66744),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i237_LC_17_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i237_LC_17_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i237_LC_17_19_2 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i237_LC_17_19_2  (
            .in0(N__63123),
            .in1(N__44559),
            .in2(N__62205),
            .in3(N__67621),
            .lcout(\c0.data_in_frame_29_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66744),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_17_i3_2_lut_4_lut_LC_17_19_3 .C_ON=1'b0;
    defparam \c0.select_365_Select_17_i3_2_lut_4_lut_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_17_i3_2_lut_4_lut_LC_17_19_3 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \c0.select_365_Select_17_i3_2_lut_4_lut_LC_17_19_3  (
            .in0(N__50650),
            .in1(N__51398),
            .in2(N__45502),
            .in3(N__50826),
            .lcout(\c0.n3_adj_4448 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1388_LC_17_19_5 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1388_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1388_LC_17_19_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i17_4_lut_adj_1388_LC_17_19_5  (
            .in0(N__50059),
            .in1(N__44863),
            .in2(N__53956),
            .in3(N__44734),
            .lcout(n23726),
            .ltout(n23726_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i6_LC_17_19_6 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i6_LC_17_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i6_LC_17_19_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.control_mode_i0_i6_LC_17_19_6  (
            .in0(N__43822),
            .in1(_gnd_net_),
            .in2(N__42310),
            .in3(N__42293),
            .lcout(control_mode_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66744),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i235_LC_17_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i235_LC_17_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i235_LC_17_19_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i235_LC_17_19_7  (
            .in0(N__67620),
            .in1(N__68395),
            .in2(N__44899),
            .in3(N__62197),
            .lcout(\c0.data_in_frame_29_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66744),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_19_i3_2_lut_4_lut_LC_17_20_1 .C_ON=1'b0;
    defparam \c0.select_365_Select_19_i3_2_lut_4_lut_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_19_i3_2_lut_4_lut_LC_17_20_1 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \c0.select_365_Select_19_i3_2_lut_4_lut_LC_17_20_1  (
            .in0(N__50778),
            .in1(N__51388),
            .in2(N__45535),
            .in3(N__50594),
            .lcout(\c0.n3_adj_4444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i206_LC_17_20_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i206_LC_17_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i206_LC_17_20_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i206_LC_17_20_2  (
            .in0(N__69864),
            .in1(N__67202),
            .in2(N__53598),
            .in3(N__67623),
            .lcout(\c0.data_in_frame_25_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66758),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1581_LC_17_20_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1581_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1581_LC_17_20_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_1581_LC_17_20_3  (
            .in0(N__44817),
            .in1(N__46039),
            .in2(_gnd_net_),
            .in3(N__45073),
            .lcout(\c0.n12876 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_4_lut_LC_17_20_4 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_4_lut_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_4_lut_LC_17_20_4 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.i4_2_lut_3_lut_4_lut_LC_17_20_4  (
            .in0(N__43342),
            .in1(N__43363),
            .in2(N__48953),
            .in3(N__50777),
            .lcout(\c0.n21022 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_18_i3_2_lut_4_lut_LC_17_20_5 .C_ON=1'b0;
    defparam \c0.select_365_Select_18_i3_2_lut_4_lut_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_18_i3_2_lut_4_lut_LC_17_20_5 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \c0.select_365_Select_18_i3_2_lut_4_lut_LC_17_20_5  (
            .in0(N__50779),
            .in1(N__51389),
            .in2(N__45583),
            .in3(N__50595),
            .lcout(\c0.n3_adj_4446 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i233_LC_17_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i233_LC_17_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i233_LC_17_20_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i233_LC_17_20_6  (
            .in0(N__62189),
            .in1(N__69487),
            .in2(N__44791),
            .in3(N__67624),
            .lcout(\c0.data_in_frame_29_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66758),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1531_LC_17_21_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1531_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1531_LC_17_21_0 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \c0.i1_4_lut_adj_1531_LC_17_21_0  (
            .in0(N__42786),
            .in1(N__42585),
            .in2(N__42567),
            .in3(N__42409),
            .lcout(\c0.n5_adj_4342 ),
            .ltout(\c0.n5_adj_4342_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i3_LC_17_21_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i3_LC_17_21_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i3_LC_17_21_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \c0.FRAME_MATCHER_state_i3_LC_17_21_1  (
            .in0(N__42494),
            .in1(_gnd_net_),
            .in2(N__42550),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66771),
            .ce(),
            .sr(N__42445));
    defparam \c0.i3_3_lut_4_lut_adj_1749_LC_17_21_2 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_1749_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_1749_LC_17_21_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_1749_LC_17_21_2  (
            .in0(N__43362),
            .in1(N__43345),
            .in2(N__48981),
            .in3(N__50802),
            .lcout(\c0.n21686 ),
            .ltout(\c0.n21686_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_4_lut_LC_17_21_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_4_lut_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_4_lut_LC_17_21_3 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \c0.i1_4_lut_4_lut_LC_17_21_3  (
            .in0(N__42493),
            .in1(N__53188),
            .in2(N__42448),
            .in3(N__42787),
            .lcout(\c0.n21334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1530_LC_17_21_4 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1530_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1530_LC_17_21_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \c0.i1_3_lut_adj_1530_LC_17_21_4  (
            .in0(N__42785),
            .in1(N__42429),
            .in2(_gnd_net_),
            .in3(N__43344),
            .lcout(\c0.n1_adj_4349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i48_4_lut_LC_17_21_6 .C_ON=1'b0;
    defparam \c0.i48_4_lut_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i48_4_lut_LC_17_21_6 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.i48_4_lut_LC_17_21_6  (
            .in0(N__43361),
            .in1(N__43343),
            .in2(N__43306),
            .in3(N__43290),
            .lcout(\c0.n45_adj_4389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i26_LC_17_22_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i26_LC_17_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i26_LC_17_22_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i26_LC_17_22_3  (
            .in0(N__43031),
            .in1(N__43171),
            .in2(_gnd_net_),
            .in3(N__63769),
            .lcout(data_in_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66785),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1534_LC_17_22_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1534_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1534_LC_17_22_4 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_4_lut_adj_1534_LC_17_22_4  (
            .in0(N__42649),
            .in1(N__43009),
            .in2(N__43502),
            .in3(N__53026),
            .lcout(\c0.n21332 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14222_2_lut_LC_17_22_6 .C_ON=1'b0;
    defparam \c0.i14222_2_lut_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i14222_2_lut_LC_17_22_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i14222_2_lut_LC_17_22_6  (
            .in0(_gnd_net_),
            .in1(N__46158),
            .in2(_gnd_net_),
            .in3(N__42971),
            .lcout(\c0.n937 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i178_LC_17_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i178_LC_17_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i178_LC_17_22_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i178_LC_17_22_7  (
            .in0(N__44925),
            .in1(N__63768),
            .in2(_gnd_net_),
            .in3(N__59210),
            .lcout(data_in_frame_22_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66785),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1757_LC_17_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1757_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1757_LC_17_23_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1757_LC_17_23_1  (
            .in0(N__42935),
            .in1(N__53131),
            .in2(_gnd_net_),
            .in3(N__53019),
            .lcout(\c0.n21352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i179_LC_17_23_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i179_LC_17_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i179_LC_17_23_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i179_LC_17_23_2  (
            .in0(N__68352),
            .in1(N__59310),
            .in2(_gnd_net_),
            .in3(N__59211),
            .lcout(data_in_frame_22_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66795),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1747_LC_17_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1747_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1747_LC_17_23_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1747_LC_17_23_3  (
            .in0(N__42885),
            .in1(N__42826),
            .in2(_gnd_net_),
            .in3(N__42788),
            .lcout(\c0.n7_adj_4356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1758_LC_17_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1758_LC_17_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1758_LC_17_23_4 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1758_LC_17_23_4  (
            .in0(N__53020),
            .in1(_gnd_net_),
            .in2(N__53174),
            .in3(N__43451),
            .lcout(\c0.n21354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1777_LC_17_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1777_LC_17_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1777_LC_17_23_5 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1777_LC_17_23_5  (
            .in0(N__43531),
            .in1(N__53135),
            .in2(_gnd_net_),
            .in3(N__53021),
            .lcout(\c0.n21378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i240_LC_17_23_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i240_LC_17_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i240_LC_17_23_6 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i240_LC_17_23_6  (
            .in0(N__68880),
            .in1(N__50034),
            .in2(N__62204),
            .in3(N__67685),
            .lcout(\c0.data_in_frame_29_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66795),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i28_LC_17_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i28_LC_17_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i28_LC_17_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i28_LC_17_24_0  (
            .in0(_gnd_net_),
            .in1(N__43532),
            .in2(_gnd_net_),
            .in3(N__52744),
            .lcout(\c0.FRAME_MATCHER_state_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66805),
            .ce(),
            .sr(N__43510));
    defparam \c0.FRAME_MATCHER_state_i31_LC_17_25_4 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i31_LC_17_25_4 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i31_LC_17_25_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i31_LC_17_25_4  (
            .in0(_gnd_net_),
            .in1(N__43487),
            .in2(_gnd_net_),
            .in3(N__52844),
            .lcout(\c0.FRAME_MATCHER_state_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66817),
            .ce(),
            .sr(N__43465));
    defparam \c0.FRAME_MATCHER_state_i13_LC_17_26_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i13_LC_17_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i13_LC_17_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i13_LC_17_26_0  (
            .in0(_gnd_net_),
            .in1(N__43444),
            .in2(_gnd_net_),
            .in3(N__52846),
            .lcout(\c0.FRAME_MATCHER_state_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66829),
            .ce(),
            .sr(N__43420));
    defparam \c0.FRAME_MATCHER_state_i15_LC_17_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i15_LC_17_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i15_LC_17_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i15_LC_17_27_0  (
            .in0(_gnd_net_),
            .in1(N__43394),
            .in2(_gnd_net_),
            .in3(N__52745),
            .lcout(\c0.FRAME_MATCHER_state_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66841),
            .ce(),
            .sr(N__43372));
    defparam \c0.select_365_Select_0_i3_2_lut_4_lut_LC_18_3_1 .C_ON=1'b0;
    defparam \c0.select_365_Select_0_i3_2_lut_4_lut_LC_18_3_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_0_i3_2_lut_4_lut_LC_18_3_1 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_0_i3_2_lut_4_lut_LC_18_3_1  (
            .in0(N__51451),
            .in1(N__51190),
            .in2(N__56719),
            .in3(N__50680),
            .lcout(\c0.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_5_i3_2_lut_4_lut_LC_18_6_7 .C_ON=1'b0;
    defparam \c0.select_365_Select_5_i3_2_lut_4_lut_LC_18_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_5_i3_2_lut_4_lut_LC_18_6_7 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_5_i3_2_lut_4_lut_LC_18_6_7  (
            .in0(N__51471),
            .in1(N__51122),
            .in2(N__47391),
            .in3(N__50678),
            .lcout(\c0.n3_adj_4468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1680_LC_18_8_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1680_LC_18_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1680_LC_18_8_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1680_LC_18_8_0  (
            .in0(N__47725),
            .in1(N__43571),
            .in2(N__44703),
            .in3(N__51683),
            .lcout(\c0.n18_adj_4370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1550_LC_18_8_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1550_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1550_LC_18_8_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1550_LC_18_8_1  (
            .in0(N__43572),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47509),
            .lcout(\c0.n21957 ),
            .ltout(\c0.n21957_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1586_LC_18_8_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1586_LC_18_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1586_LC_18_8_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1586_LC_18_8_2  (
            .in0(N__43557),
            .in1(N__43579),
            .in2(N__43582),
            .in3(N__52054),
            .lcout(\c0.n13099 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1557_LC_18_8_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1557_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1557_LC_18_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1557_LC_18_8_3  (
            .in0(N__51684),
            .in1(N__44695),
            .in2(_gnd_net_),
            .in3(N__47726),
            .lcout(\c0.n22287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i28_LC_18_8_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i28_LC_18_8_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i28_LC_18_8_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i28_LC_18_8_4  (
            .in0(N__60867),
            .in1(N__67364),
            .in2(N__64893),
            .in3(N__43573),
            .lcout(\c0.data_in_frame_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66641),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i27_LC_18_8_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i27_LC_18_8_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i27_LC_18_8_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i27_LC_18_8_5  (
            .in0(N__67363),
            .in1(N__60869),
            .in2(N__47736),
            .in3(N__68410),
            .lcout(\c0.data_in_frame_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66641),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i45_LC_18_8_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i45_LC_18_8_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i45_LC_18_8_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i45_LC_18_8_6  (
            .in0(N__60868),
            .in1(N__63204),
            .in2(N__43561),
            .in3(N__62188),
            .lcout(\c0.data_in_frame_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66641),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i9_LC_18_8_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i9_LC_18_8_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i9_LC_18_8_7 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i9_LC_18_8_7  (
            .in0(N__44702),
            .in1(N__69567),
            .in2(N__69777),
            .in3(N__60870),
            .lcout(data_in_frame_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66641),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20143_4_lut_LC_18_9_0 .C_ON=1'b0;
    defparam \c0.i20143_4_lut_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i20143_4_lut_LC_18_9_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i20143_4_lut_LC_18_9_0  (
            .in0(N__47540),
            .in1(N__44050),
            .in2(N__44505),
            .in3(N__47501),
            .lcout(\c0.n23838 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1603_LC_18_9_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1603_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1603_LC_18_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1603_LC_18_9_2  (
            .in0(N__51685),
            .in1(N__44696),
            .in2(_gnd_net_),
            .in3(N__43644),
            .lcout(\c0.n21902 ),
            .ltout(\c0.n21902_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1609_LC_18_9_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1609_LC_18_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1609_LC_18_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1609_LC_18_9_3  (
            .in0(N__44697),
            .in1(N__51776),
            .in2(N__43651),
            .in3(N__47539),
            .lcout(\c0.n21992 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i24_LC_18_9_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i24_LC_18_9_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i24_LC_18_9_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i24_LC_18_9_4  (
            .in0(N__69168),
            .in1(N__68956),
            .in2(N__47547),
            .in3(N__60896),
            .lcout(\c0.data_in_frame_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66648),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i25_LC_18_9_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i25_LC_18_9_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i25_LC_18_9_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i25_LC_18_9_5  (
            .in0(N__60894),
            .in1(N__69548),
            .in2(N__43648),
            .in3(N__67379),
            .lcout(\c0.data_in_frame_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66648),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1540_LC_18_9_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1540_LC_18_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1540_LC_18_9_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1540_LC_18_9_6  (
            .in0(N__43636),
            .in1(N__47762),
            .in2(N__43629),
            .in3(N__47500),
            .lcout(\c0.n10_adj_4363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i7_LC_18_9_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i7_LC_18_9_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i7_LC_18_9_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i7_LC_18_9_7  (
            .in0(N__60895),
            .in1(N__51686),
            .in2(N__65647),
            .in3(N__65969),
            .lcout(\c0.data_in_frame_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66648),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i26_LC_18_10_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i26_LC_18_10_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i26_LC_18_10_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i26_LC_18_10_0  (
            .in0(N__67362),
            .in1(N__60846),
            .in2(N__47767),
            .in3(N__63863),
            .lcout(\c0.data_in_frame_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66655),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1679_LC_18_10_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1679_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1679_LC_18_10_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1679_LC_18_10_1  (
            .in0(N__54400),
            .in1(N__52034),
            .in2(N__47693),
            .in3(N__48026),
            .lcout(),
            .ltout(\c0.n21879_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1566_LC_18_10_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1566_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1566_LC_18_10_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1566_LC_18_10_2  (
            .in0(N__61092),
            .in1(N__47758),
            .in2(N__43612),
            .in3(N__44355),
            .lcout(\c0.n29_adj_4374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1554_LC_18_10_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1554_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1554_LC_18_10_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1554_LC_18_10_3  (
            .in0(_gnd_net_),
            .in1(N__47992),
            .in2(_gnd_net_),
            .in3(N__43604),
            .lcout(\c0.n22051 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i8_LC_18_10_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i8_LC_18_10_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i8_LC_18_10_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i8_LC_18_10_4  (
            .in0(N__47493),
            .in1(N__68955),
            .in2(N__66029),
            .in3(N__60847),
            .lcout(\c0.data_in_frame_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66655),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i38_LC_18_10_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i38_LC_18_10_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i38_LC_18_10_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i38_LC_18_10_5  (
            .in0(N__60845),
            .in1(N__64532),
            .in2(N__67210),
            .in3(N__61093),
            .lcout(\c0.data_in_frame_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66655),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1612_LC_18_10_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1612_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1612_LC_18_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1612_LC_18_10_6  (
            .in0(_gnd_net_),
            .in1(N__51775),
            .in2(N__47508),
            .in3(N__51687),
            .lcout(\c0.n22194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1556_LC_18_10_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1556_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1556_LC_18_10_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1556_LC_18_10_7  (
            .in0(N__47684),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48027),
            .lcout(\c0.n22290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1590_LC_18_11_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1590_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1590_LC_18_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1590_LC_18_11_0  (
            .in0(_gnd_net_),
            .in1(N__49597),
            .in2(_gnd_net_),
            .in3(N__43970),
            .lcout(\c0.n22258 ),
            .ltout(\c0.n22258_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1569_LC_18_11_1 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1569_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1569_LC_18_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1569_LC_18_11_1  (
            .in0(N__44221),
            .in1(N__47615),
            .in2(N__43675),
            .in3(N__51990),
            .lcout(),
            .ltout(\c0.n27_adj_4377_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1570_LC_18_11_2 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1570_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1570_LC_18_11_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_1570_LC_18_11_2  (
            .in0(N__43672),
            .in1(N__43927),
            .in2(N__43666),
            .in3(N__43696),
            .lcout(\c0.n14072 ),
            .ltout(\c0.n14072_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1549_LC_18_11_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1549_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1549_LC_18_11_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1549_LC_18_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43663),
            .in3(N__54363),
            .lcout(\c0.n13852 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1672_LC_18_11_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1672_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1672_LC_18_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1672_LC_18_11_4  (
            .in0(N__47616),
            .in1(N__43951),
            .in2(N__48208),
            .in3(N__43660),
            .lcout(),
            .ltout(\c0.n6_adj_4385_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1583_LC_18_11_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1583_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1583_LC_18_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1583_LC_18_11_5  (
            .in0(N__43971),
            .in1(N__44419),
            .in2(N__43654),
            .in3(N__43809),
            .lcout(\c0.n14113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1605_LC_18_11_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1605_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1605_LC_18_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1605_LC_18_11_6  (
            .in0(_gnd_net_),
            .in1(N__48139),
            .in2(_gnd_net_),
            .in3(N__50339),
            .lcout(\c0.n21803 ),
            .ltout(\c0.n21803_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1559_LC_18_11_7 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1559_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1559_LC_18_11_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1559_LC_18_11_7  (
            .in0(N__43945),
            .in1(N__43936),
            .in2(N__43930),
            .in3(N__44014),
            .lcout(\c0.n30_adj_4371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1551_LC_18_12_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1551_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1551_LC_18_12_0 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \c0.i2_3_lut_adj_1551_LC_18_12_0  (
            .in0(N__44336),
            .in1(N__43900),
            .in2(N__43879),
            .in3(_gnd_net_),
            .lcout(\c0.n13376 ),
            .ltout(\c0.n13376_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1560_LC_18_12_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1560_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1560_LC_18_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1560_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(N__43806),
            .in2(N__43837),
            .in3(N__44292),
            .lcout(\c0.n22320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1669_LC_18_12_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1669_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1669_LC_18_12_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1669_LC_18_12_2  (
            .in0(N__43808),
            .in1(N__43834),
            .in2(N__44308),
            .in3(N__44444),
            .lcout(\c0.n6_adj_4386 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1594_LC_18_12_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1594_LC_18_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1594_LC_18_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1594_LC_18_12_3  (
            .in0(N__47632),
            .in1(N__44293),
            .in2(_gnd_net_),
            .in3(N__43807),
            .lcout(),
            .ltout(\c0.n13386_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1621_LC_18_12_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1621_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1621_LC_18_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1621_LC_18_12_4  (
            .in0(N__54367),
            .in1(N__43770),
            .in2(N__43759),
            .in3(N__44065),
            .lcout(\c0.n13033 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1607_LC_18_12_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1607_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1607_LC_18_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1607_LC_18_12_5  (
            .in0(N__43751),
            .in1(N__49634),
            .in2(N__44049),
            .in3(N__44012),
            .lcout(\c0.n22261 ),
            .ltout(\c0.n22261_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1561_LC_18_12_6 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1561_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1561_LC_18_12_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_1561_LC_18_12_6  (
            .in0(N__44064),
            .in1(N__43723),
            .in2(N__43705),
            .in3(N__43702),
            .lcout(\c0.n28_adj_4372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1558_LC_18_12_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1558_LC_18_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1558_LC_18_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1558_LC_18_12_7  (
            .in0(N__44443),
            .in1(N__44103),
            .in2(_gnd_net_),
            .in3(N__44078),
            .lcout(\c0.n22218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1553_LC_18_13_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1553_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1553_LC_18_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1553_LC_18_13_0  (
            .in0(N__44203),
            .in1(N__44398),
            .in2(N__44541),
            .in3(N__44191),
            .lcout(\c0.n21928 ),
            .ltout(\c0.n21928_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1542_LC_18_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1542_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1542_LC_18_13_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1542_LC_18_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44053),
            .in3(N__44469),
            .lcout(\c0.n13861 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1595_LC_18_13_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1595_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1595_LC_18_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1595_LC_18_13_2  (
            .in0(N__44038),
            .in1(N__44013),
            .in2(N__44542),
            .in3(N__48089),
            .lcout(\c0.n21882 ),
            .ltout(\c0.n21882_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1539_LC_18_13_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1539_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1539_LC_18_13_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1539_LC_18_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43993),
            .in3(N__61103),
            .lcout(\c0.data_out_frame_0__7__N_2744 ),
            .ltout(\c0.data_out_frame_0__7__N_2744_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_LC_18_13_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_LC_18_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_LC_18_13_4  (
            .in0(N__44362),
            .in1(N__48090),
            .in2(N__43978),
            .in3(N__44399),
            .lcout(),
            .ltout(\c0.n6_adj_4272_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1334_LC_18_13_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1334_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1334_LC_18_13_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1334_LC_18_13_5  (
            .in0(N__44379),
            .in1(N__44251),
            .in2(N__43975),
            .in3(N__54815),
            .lcout(\c0.n22069 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i32_LC_18_13_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i32_LC_18_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i32_LC_18_13_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i32_LC_18_13_6  (
            .in0(N__60823),
            .in1(N__67361),
            .in2(N__43972),
            .in3(N__68975),
            .lcout(\c0.data_in_frame_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66677),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1537_LC_18_13_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1537_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1537_LC_18_13_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1537_LC_18_13_7  (
            .in0(N__44400),
            .in1(N__44378),
            .in2(N__48094),
            .in3(N__44361),
            .lcout(\c0.n4_adj_4255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_1632_LC_18_14_0 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_1632_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_1632_LC_18_14_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \c0.i15_4_lut_adj_1632_LC_18_14_0  (
            .in0(N__50307),
            .in1(N__47701),
            .in2(N__44343),
            .in3(N__44310),
            .lcout(\c0.n39_adj_4406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1330_LC_18_14_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1330_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1330_LC_18_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1330_LC_18_14_1  (
            .in0(N__44256),
            .in1(N__61124),
            .in2(_gnd_net_),
            .in3(N__44227),
            .lcout(\c0.n14037 ),
            .ltout(\c0.n14037_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1787_LC_18_14_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1787_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1787_LC_18_14_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1787_LC_18_14_2  (
            .in0(N__44220),
            .in1(_gnd_net_),
            .in2(N__44206),
            .in3(N__44468),
            .lcout(\c0.n22108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1681_LC_18_14_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1681_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1681_LC_18_14_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1681_LC_18_14_3  (
            .in0(N__44491),
            .in1(N__48154),
            .in2(N__44146),
            .in3(N__50368),
            .lcout(\c0.n6_adj_4369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1552_LC_18_14_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1552_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1552_LC_18_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1552_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(N__44135),
            .in2(N__48169),
            .in3(N__44492),
            .lcout(\c0.n5_adj_4368 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__5__I_0_2_lut_LC_18_14_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__5__I_0_2_lut_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.data_in_frame_0__5__I_0_2_lut_LC_18_14_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_in_frame_0__5__I_0_2_lut_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(N__51774),
            .in2(_gnd_net_),
            .in3(N__50306),
            .lcout(\c0.data_out_frame_29__7__N_1474 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i55_LC_18_14_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i55_LC_18_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i55_LC_18_14_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i55_LC_18_14_6  (
            .in0(N__65649),
            .in1(N__49674),
            .in2(_gnd_net_),
            .in3(N__44181),
            .lcout(data_in_frame_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66689),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i3_LC_18_14_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i3_LC_18_14_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i3_LC_18_14_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i3_LC_18_14_7  (
            .in0(N__60715),
            .in1(N__65865),
            .in2(N__68411),
            .in3(N__44145),
            .lcout(\c0.data_in_frame_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66689),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i21_LC_18_15_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i21_LC_18_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i21_LC_18_15_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i21_LC_18_15_0  (
            .in0(N__69212),
            .in1(N__60756),
            .in2(N__44506),
            .in3(N__63171),
            .lcout(\c0.data_in_frame_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66703),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_9_i3_2_lut_4_lut_LC_18_15_1 .C_ON=1'b0;
    defparam \c0.select_365_Select_9_i3_2_lut_4_lut_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_9_i3_2_lut_4_lut_LC_18_15_1 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \c0.select_365_Select_9_i3_2_lut_4_lut_LC_18_15_1  (
            .in0(N__51444),
            .in1(N__50659),
            .in2(N__45280),
            .in3(N__50962),
            .lcout(\c0.n3_adj_4462 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i41_LC_18_15_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i41_LC_18_15_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i41_LC_18_15_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i41_LC_18_15_2  (
            .in0(N__69559),
            .in1(N__60757),
            .in2(N__44473),
            .in3(N__62198),
            .lcout(\c0.data_in_frame_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66703),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1202_LC_18_15_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1202_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1202_LC_18_15_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1202_LC_18_15_3  (
            .in0(N__62590),
            .in1(N__65155),
            .in2(N__62822),
            .in3(N__63388),
            .lcout(\c0.n22057 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i48_LC_18_15_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i48_LC_18_15_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i48_LC_18_15_4 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i48_LC_18_15_4  (
            .in0(N__68944),
            .in1(N__60758),
            .in2(N__62206),
            .in3(N__47883),
            .lcout(\c0.data_in_frame_5_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66703),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_6_i3_2_lut_4_lut_LC_18_15_5 .C_ON=1'b0;
    defparam \c0.select_365_Select_6_i3_2_lut_4_lut_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_6_i3_2_lut_4_lut_LC_18_15_5 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \c0.select_365_Select_6_i3_2_lut_4_lut_LC_18_15_5  (
            .in0(N__51443),
            .in1(N__50658),
            .in2(N__47359),
            .in3(N__50961),
            .lcout(\c0.n3_adj_4467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1574_LC_18_15_6 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1574_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1574_LC_18_15_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i11_4_lut_adj_1574_LC_18_15_6  (
            .in0(N__47355),
            .in1(N__45225),
            .in2(N__47401),
            .in3(N__45534),
            .lcout(\c0.n28_adj_4381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i17_LC_18_15_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i17_LC_18_15_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i17_LC_18_15_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i17_LC_18_15_7  (
            .in0(N__60755),
            .in1(N__69213),
            .in2(N__44448),
            .in3(N__69558),
            .lcout(\c0.data_in_frame_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66703),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i204_LC_18_16_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i204_LC_18_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i204_LC_18_16_0 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i204_LC_18_16_0  (
            .in0(N__64698),
            .in1(N__53626),
            .in2(N__69866),
            .in3(N__67611),
            .lcout(\c0.data_in_frame_25_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66717),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i50_LC_18_16_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i50_LC_18_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i50_LC_18_16_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i50_LC_18_16_1  (
            .in0(N__63781),
            .in1(N__49703),
            .in2(_gnd_net_),
            .in3(N__44415),
            .lcout(data_in_frame_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66717),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i177_LC_18_16_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i177_LC_18_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i177_LC_18_16_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i177_LC_18_16_2  (
            .in0(N__69486),
            .in1(N__62815),
            .in2(_gnd_net_),
            .in3(N__59169),
            .lcout(data_in_frame_22_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66717),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i36_LC_18_16_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i36_LC_18_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i36_LC_18_16_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i36_LC_18_16_3  (
            .in0(N__64818),
            .in1(N__60714),
            .in2(N__49642),
            .in3(N__64531),
            .lcout(\c0.data_in_frame_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66717),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_1176_LC_18_16_4 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_1176_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_1176_LC_18_16_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.rx.i1_2_lut_adj_1176_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(N__59883),
            .in2(_gnd_net_),
            .in3(N__57105),
            .lcout(n4),
            .ltout(n4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i2_LC_18_16_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i2_LC_18_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i2_LC_18_16_5 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.rx.r_Rx_Byte_i2_LC_18_16_5  (
            .in0(N__59694),
            .in1(N__68289),
            .in2(N__44545),
            .in3(N__59944),
            .lcout(rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66717),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i39_LC_18_16_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i39_LC_18_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i39_LC_18_16_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i39_LC_18_16_6  (
            .in0(N__60713),
            .in1(N__65697),
            .in2(N__64556),
            .in3(N__44534),
            .lcout(\c0.data_in_frame_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66717),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i3_LC_18_16_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i3_LC_18_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i3_LC_18_16_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i3_LC_18_16_7  (
            .in0(N__44518),
            .in1(N__64699),
            .in2(N__59710),
            .in3(N__56221),
            .lcout(rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66717),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_16_i3_2_lut_4_lut_LC_18_17_1 .C_ON=1'b0;
    defparam \c0.select_365_Select_16_i3_2_lut_4_lut_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_16_i3_2_lut_4_lut_LC_18_17_1 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_16_i3_2_lut_4_lut_LC_18_17_1  (
            .in0(N__51448),
            .in1(N__50954),
            .in2(N__49897),
            .in3(N__50651),
            .lcout(\c0.n3_adj_4450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1466_LC_18_17_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1466_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1466_LC_18_17_2 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_adj_1466_LC_18_17_2  (
            .in0(N__46049),
            .in1(N__45064),
            .in2(N__47321),
            .in3(N__44723),
            .lcout(\c0.n21758 ),
            .ltout(\c0.n21758_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i162_LC_18_17_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i162_LC_18_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i162_LC_18_17_3 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i162_LC_18_17_3  (
            .in0(N__63814),
            .in1(N__64527),
            .in2(N__44509),
            .in3(N__53241),
            .lcout(\c0.data_in_frame_20_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66731),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1457_LC_18_17_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1457_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1457_LC_18_17_4 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_adj_1457_LC_18_17_4  (
            .in0(N__46050),
            .in1(N__45065),
            .in2(N__47322),
            .in3(N__44724),
            .lcout(\c0.n21749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1240_LC_18_17_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1240_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1240_LC_18_17_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1240_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(N__55432),
            .in2(_gnd_net_),
            .in3(N__61430),
            .lcout(\c0.n22308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i212_LC_18_17_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i212_LC_18_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i212_LC_18_17_7 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i212_LC_18_17_7  (
            .in0(N__64700),
            .in1(N__57987),
            .in2(N__69253),
            .in3(N__67678),
            .lcout(\c0.data_in_frame_26_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66731),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i234_LC_18_18_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i234_LC_18_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i234_LC_18_18_0 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i234_LC_18_18_0  (
            .in0(N__67609),
            .in1(N__44880),
            .in2(N__62190),
            .in3(N__63825),
            .lcout(\c0.data_in_frame_29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66745),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1571_LC_18_18_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1571_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1571_LC_18_18_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_1571_LC_18_18_1  (
            .in0(N__45327),
            .in1(N__45174),
            .in2(N__45385),
            .in3(N__45435),
            .lcout(\c0.n17_adj_4378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i141_LC_18_18_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i141_LC_18_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i141_LC_18_18_3 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i141_LC_18_18_3  (
            .in0(N__63145),
            .in1(N__67912),
            .in2(N__69881),
            .in3(N__55375),
            .lcout(\c0.data_in_frame_17_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66745),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i0_LC_18_18_4 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i0_LC_18_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i0_LC_18_18_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i0_LC_18_18_4  (
            .in0(N__44591),
            .in1(N__44710),
            .in2(_gnd_net_),
            .in3(N__44660),
            .lcout(control_mode_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66745),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_97_i9_2_lut_3_lut_LC_18_18_5 .C_ON=1'b0;
    defparam \c0.equal_97_i9_2_lut_3_lut_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.equal_97_i9_2_lut_3_lut_LC_18_18_5 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \c0.equal_97_i9_2_lut_3_lut_LC_18_18_5  (
            .in0(N__56467),
            .in1(_gnd_net_),
            .in2(N__56744),
            .in3(N__56600),
            .lcout(\c0.n9_adj_4278 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i137_LC_18_18_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i137_LC_18_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i137_LC_18_18_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i137_LC_18_18_7  (
            .in0(N__69860),
            .in1(N__67911),
            .in2(N__55627),
            .in3(N__69491),
            .lcout(\c0.data_in_frame_17_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66745),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1376_LC_18_19_0 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1376_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1376_LC_18_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_1376_LC_18_19_0  (
            .in0(N__56057),
            .in1(N__56279),
            .in2(N__44560),
            .in3(N__53743),
            .lcout(\c0.n23523 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1362_LC_18_19_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1362_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1362_LC_18_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1362_LC_18_19_1  (
            .in0(N__58609),
            .in1(N__65326),
            .in2(N__44803),
            .in3(N__64990),
            .lcout(),
            .ltout(\c0.n10_adj_4286_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1374_LC_18_19_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1374_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1374_LC_18_19_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i5_3_lut_adj_1374_LC_18_19_2  (
            .in0(N__54016),
            .in1(_gnd_net_),
            .in2(N__44806),
            .in3(N__59983),
            .lcout(\c0.n23389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i190_LC_18_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i190_LC_18_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i190_LC_18_19_3 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \c0.data_in_frame_0__i190_LC_18_19_3  (
            .in0(N__68632),
            .in1(N__67206),
            .in2(N__68044),
            .in3(N__49919),
            .lcout(\c0.data_in_frame_23_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66759),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i227_LC_18_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i227_LC_18_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i227_LC_18_19_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i227_LC_18_19_4  (
            .in0(N__67731),
            .in1(N__44802),
            .in2(N__64567),
            .in3(N__68394),
            .lcout(\c0.data_in_frame_28_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66759),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i230_LC_18_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i230_LC_18_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i230_LC_18_19_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i230_LC_18_19_5  (
            .in0(N__64566),
            .in1(N__67207),
            .in2(N__58377),
            .in3(N__67733),
            .lcout(\c0.data_in_frame_28_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66759),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i203_LC_18_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i203_LC_18_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i203_LC_18_19_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i203_LC_18_19_7  (
            .in0(N__68393),
            .in1(N__69865),
            .in2(N__53694),
            .in3(N__67732),
            .lcout(\c0.data_in_frame_25_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66759),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1375_LC_18_20_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1375_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1375_LC_18_20_0 .LUT_INIT=16'b1101111011101101;
    LogicCell40 \c0.i1_4_lut_adj_1375_LC_18_20_0  (
            .in0(N__44790),
            .in1(N__44773),
            .in2(N__53533),
            .in3(N__58866),
            .lcout(),
            .ltout(\c0.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1378_LC_18_20_1 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1378_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1378_LC_18_20_1 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i14_4_lut_adj_1378_LC_18_20_1  (
            .in0(N__59461),
            .in1(N__56233),
            .in2(N__44755),
            .in3(N__44752),
            .lcout(),
            .ltout(\c0.n32_adj_4295_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1386_LC_18_20_2 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1386_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1386_LC_18_20_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i16_4_lut_adj_1386_LC_18_20_2  (
            .in0(N__58357),
            .in1(N__54070),
            .in2(N__44746),
            .in3(N__44743),
            .lcout(\c0.n34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1367_LC_18_20_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1367_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1367_LC_18_20_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_1367_LC_18_20_3  (
            .in0(N__58867),
            .in1(N__55798),
            .in2(N__44898),
            .in3(N__50205),
            .lcout(),
            .ltout(\c0.n23388_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1385_LC_18_20_4 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1385_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1385_LC_18_20_4 .LUT_INIT=16'b1111111111110110;
    LogicCell40 \c0.i12_4_lut_adj_1385_LC_18_20_4  (
            .in0(N__53532),
            .in1(N__44881),
            .in2(N__44866),
            .in3(N__64972),
            .lcout(\c0.n30_adj_4299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1577_LC_18_21_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1577_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1577_LC_18_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i10_4_lut_adj_1577_LC_18_21_0  (
            .in0(N__49822),
            .in1(N__45838),
            .in2(N__45802),
            .in3(N__45715),
            .lcout(\c0.n27_adj_4383 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_adj_1568_LC_18_21_2 .C_ON=1'b0;
    defparam \c0.i5_2_lut_adj_1568_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_adj_1568_LC_18_21_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i5_2_lut_adj_1568_LC_18_21_2  (
            .in0(N__45877),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45279),
            .lcout(),
            .ltout(\c0.n15_adj_4376_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1572_LC_18_21_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1572_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1572_LC_18_21_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_4_lut_adj_1572_LC_18_21_3  (
            .in0(N__50157),
            .in1(N__49873),
            .in2(N__44857),
            .in3(N__44854),
            .lcout(),
            .ltout(\c0.n18_adj_4379_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1573_LC_18_21_4 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1573_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1573_LC_18_21_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i13_4_lut_adj_1573_LC_18_21_4  (
            .in0(N__45630),
            .in1(N__45498),
            .in2(N__44845),
            .in3(N__45579),
            .lcout(),
            .ltout(\c0.n30_adj_4380_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1579_LC_18_21_5 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1579_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1579_LC_18_21_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i16_4_lut_adj_1579_LC_18_21_5  (
            .in0(N__44842),
            .in1(N__44965),
            .in2(N__44836),
            .in3(N__44833),
            .lcout(\c0.n13000 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_adj_1731_LC_18_22_0 .C_ON=1'b0;
    defparam \c0.i20_4_lut_adj_1731_LC_18_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_adj_1731_LC_18_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_4_lut_adj_1731_LC_18_22_0  (
            .in0(N__66136),
            .in1(N__59117),
            .in2(N__56149),
            .in3(N__53560),
            .lcout(\c0.n49_adj_4488 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_22_i3_2_lut_4_lut_LC_18_22_1 .C_ON=1'b0;
    defparam \c0.select_365_Select_22_i3_2_lut_4_lut_LC_18_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_22_i3_2_lut_4_lut_LC_18_22_1 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \c0.select_365_Select_22_i3_2_lut_4_lut_LC_18_22_1  (
            .in0(N__50646),
            .in1(N__51412),
            .in2(N__51070),
            .in3(N__45675),
            .lcout(\c0.n3_adj_4438 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_21_i3_2_lut_4_lut_LC_18_22_2 .C_ON=1'b0;
    defparam \c0.select_365_Select_21_i3_2_lut_4_lut_LC_18_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_21_i3_2_lut_4_lut_LC_18_22_2 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_21_i3_2_lut_4_lut_LC_18_22_2  (
            .in0(N__51413),
            .in1(N__50987),
            .in2(N__45640),
            .in3(N__50647),
            .lcout(\c0.n3_adj_4440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i220_LC_18_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i220_LC_18_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i220_LC_18_22_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i220_LC_18_22_3  (
            .in0(N__67403),
            .in1(N__64823),
            .in2(N__56284),
            .in3(N__67762),
            .lcout(\c0.data_in_frame_27_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66796),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i211_LC_18_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i211_LC_18_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i211_LC_18_22_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i211_LC_18_22_4  (
            .in0(N__67760),
            .in1(N__59118),
            .in2(N__69234),
            .in3(N__68359),
            .lcout(\c0.data_in_frame_26_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66796),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i219_LC_18_22_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i219_LC_18_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i219_LC_18_22_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i219_LC_18_22_5  (
            .in0(N__68358),
            .in1(N__67452),
            .in2(N__56058),
            .in3(N__67761),
            .lcout(\c0.data_in_frame_27_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66796),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1213_LC_18_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1213_LC_18_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1213_LC_18_23_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1213_LC_18_23_5  (
            .in0(_gnd_net_),
            .in1(N__59306),
            .in2(_gnd_net_),
            .in3(N__44921),
            .lcout(\c0.n22191 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_23_i3_2_lut_4_lut_LC_18_24_1 .C_ON=1'b0;
    defparam \c0.select_365_Select_23_i3_2_lut_4_lut_LC_18_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_23_i3_2_lut_4_lut_LC_18_24_1 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_23_i3_2_lut_4_lut_LC_18_24_1  (
            .in0(N__51450),
            .in1(N__51068),
            .in2(N__45714),
            .in3(N__50649),
            .lcout(\c0.n3_adj_4436 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i18920_2_lut_3_lut_LC_18_24_3 .C_ON=1'b0;
    defparam \c0.rx.i18920_2_lut_3_lut_LC_18_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i18920_2_lut_3_lut_LC_18_24_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.rx.i18920_2_lut_3_lut_LC_18_24_3  (
            .in0(N__56826),
            .in1(N__59655),
            .in2(_gnd_net_),
            .in3(N__56187),
            .lcout(),
            .ltout(\c0.rx.n22611_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_adj_1172_LC_18_24_4 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_1172_LC_18_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_1172_LC_18_24_4 .LUT_INIT=16'b0000000010001011;
    LogicCell40 \c0.rx.i1_4_lut_adj_1172_LC_18_24_4  (
            .in0(N__57061),
            .in1(N__56927),
            .in2(N__44905),
            .in3(N__57007),
            .lcout(\c0.rx.n17411 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3_3_lut_4_lut_LC_18_24_5 .C_ON=1'b0;
    defparam \c0.rx.i3_3_lut_4_lut_LC_18_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3_3_lut_4_lut_LC_18_24_5 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.rx.i3_3_lut_4_lut_LC_18_24_5  (
            .in0(N__56827),
            .in1(N__59653),
            .in2(N__56938),
            .in3(N__56188),
            .lcout(),
            .ltout(\c0.rx.n8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i18819_4_lut_LC_18_24_6 .C_ON=1'b0;
    defparam \c0.rx.i18819_4_lut_LC_18_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i18819_4_lut_LC_18_24_6 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \c0.rx.i18819_4_lut_LC_18_24_6  (
            .in0(N__59654),
            .in1(N__57008),
            .in2(N__44902),
            .in3(N__56828),
            .lcout(\c0.rx.n14391 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_24_i3_2_lut_4_lut_LC_18_24_7 .C_ON=1'b0;
    defparam \c0.select_365_Select_24_i3_2_lut_4_lut_LC_18_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_24_i3_2_lut_4_lut_LC_18_24_7 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_24_i3_2_lut_4_lut_LC_18_24_7  (
            .in0(N__51449),
            .in1(N__51067),
            .in2(N__45760),
            .in3(N__50648),
            .lcout(\c0.n3_adj_4435 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_30_i3_2_lut_4_lut_LC_18_25_2 .C_ON=1'b0;
    defparam \c0.select_365_Select_30_i3_2_lut_4_lut_LC_18_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_30_i3_2_lut_4_lut_LC_18_25_2 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \c0.select_365_Select_30_i3_2_lut_4_lut_LC_18_25_2  (
            .in0(N__51403),
            .in1(N__50969),
            .in2(N__50679),
            .in3(N__45943),
            .lcout(\c0.n3_adj_4426 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1576_LC_18_25_4 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1576_LC_18_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1576_LC_18_25_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i12_4_lut_adj_1576_LC_18_25_4  (
            .in0(N__45676),
            .in1(N__45903),
            .in2(N__45759),
            .in3(N__45942),
            .lcout(\c0.n29_adj_4382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_31_i3_2_lut_4_lut_LC_18_25_7 .C_ON=1'b0;
    defparam \c0.select_365_Select_31_i3_2_lut_4_lut_LC_18_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_31_i3_2_lut_4_lut_LC_18_25_7 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \c0.select_365_Select_31_i3_2_lut_4_lut_LC_18_25_7  (
            .in0(N__50667),
            .in1(N__46147),
            .in2(N__51065),
            .in3(N__51402),
            .lcout(\c0.n3_adj_4421 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_18_26_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_18_26_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_18_26_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_18_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_25_i3_2_lut_4_lut_LC_18_26_6 .C_ON=1'b0;
    defparam \c0.select_365_Select_25_i3_2_lut_4_lut_LC_18_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_25_i3_2_lut_4_lut_LC_18_26_6 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_25_i3_2_lut_4_lut_LC_18_26_6  (
            .in0(N__51410),
            .in1(N__50973),
            .in2(N__45798),
            .in3(N__50669),
            .lcout(\c0.n3_adj_4434 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_29_i3_2_lut_4_lut_LC_18_26_7 .C_ON=1'b0;
    defparam \c0.select_365_Select_29_i3_2_lut_4_lut_LC_18_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_29_i3_2_lut_4_lut_LC_18_26_7 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \c0.select_365_Select_29_i3_2_lut_4_lut_LC_18_26_7  (
            .in0(N__50668),
            .in1(N__51409),
            .in2(N__51066),
            .in3(N__45904),
            .lcout(\c0.n3_adj_4428 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_26_i3_2_lut_4_lut_LC_18_27_5 .C_ON=1'b0;
    defparam \c0.select_365_Select_26_i3_2_lut_4_lut_LC_18_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_26_i3_2_lut_4_lut_LC_18_27_5 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \c0.select_365_Select_26_i3_2_lut_4_lut_LC_18_27_5  (
            .in0(N__50980),
            .in1(N__51411),
            .in2(N__45837),
            .in3(N__50674),
            .lcout(\c0.n3_adj_4433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_27_i3_2_lut_4_lut_LC_18_28_0 .C_ON=1'b0;
    defparam \c0.select_365_Select_27_i3_2_lut_4_lut_LC_18_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_27_i3_2_lut_4_lut_LC_18_28_0 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_27_i3_2_lut_4_lut_LC_18_28_0  (
            .in0(N__51475),
            .in1(N__50974),
            .in2(N__45876),
            .in3(N__50673),
            .lcout(\c0.n3_adj_4432 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i0_LC_19_1_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i0_LC_19_1_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i0_LC_19_1_0 .LUT_INIT=16'b1001011000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i0_LC_19_1_0  (
            .in0(_gnd_net_),
            .in1(N__56630),
            .in2(N__44953),
            .in3(N__51173),
            .lcout(\c0.FRAME_MATCHER_i_0 ),
            .ltout(),
            .carryin(bfn_19_1_0_),
            .carryout(\c0.n19442 ),
            .clk(N__66630),
            .ce(),
            .sr(N__44980));
    defparam \c0.add_49_2_THRU_CRY_0_LC_19_1_1 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_0_LC_19_1_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_0_LC_19_1_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_0_LC_19_1_1  (
            .in0(_gnd_net_),
            .in1(N__47190),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19442 ),
            .carryout(\c0.n19442_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_1_LC_19_1_2 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_1_LC_19_1_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_1_LC_19_1_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_1_LC_19_1_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47215),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19442_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19442_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_2_LC_19_1_3 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_2_LC_19_1_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_2_LC_19_1_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_2_LC_19_1_3  (
            .in0(_gnd_net_),
            .in1(N__47194),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19442_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19442_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_3_LC_19_1_4 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_3_LC_19_1_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_3_LC_19_1_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_3_LC_19_1_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47216),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19442_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19442_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_4_LC_19_1_5 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_4_LC_19_1_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_4_LC_19_1_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_4_LC_19_1_5  (
            .in0(_gnd_net_),
            .in1(N__47198),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19442_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19442_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_5_LC_19_1_6 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_5_LC_19_1_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_5_LC_19_1_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_5_LC_19_1_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47217),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19442_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19442_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_6_LC_19_1_7 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_6_LC_19_1_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_6_LC_19_1_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_6_LC_19_1_7  (
            .in0(_gnd_net_),
            .in1(N__47202),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19442_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19442_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i1_LC_19_2_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i1_LC_19_2_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i1_LC_19_2_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i1_LC_19_2_0  (
            .in0(N__51100),
            .in1(N__56495),
            .in2(_gnd_net_),
            .in3(N__44968),
            .lcout(\c0.FRAME_MATCHER_i_1 ),
            .ltout(),
            .carryin(bfn_19_2_0_),
            .carryout(\c0.n19443 ),
            .clk(N__66631),
            .ce(),
            .sr(N__46060));
    defparam \c0.add_49_3_THRU_CRY_0_LC_19_2_1 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_0_LC_19_2_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_0_LC_19_2_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_0_LC_19_2_1  (
            .in0(_gnd_net_),
            .in1(N__47177),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19443 ),
            .carryout(\c0.n19443_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_1_LC_19_2_2 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_1_LC_19_2_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_1_LC_19_2_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_1_LC_19_2_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47212),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19443_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19443_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_2_LC_19_2_3 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_2_LC_19_2_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_2_LC_19_2_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_2_LC_19_2_3  (
            .in0(_gnd_net_),
            .in1(N__47181),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19443_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19443_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_3_LC_19_2_4 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_3_LC_19_2_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_3_LC_19_2_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_3_LC_19_2_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47213),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19443_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19443_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_4_LC_19_2_5 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_4_LC_19_2_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_4_LC_19_2_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_4_LC_19_2_5  (
            .in0(_gnd_net_),
            .in1(N__47185),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19443_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19443_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_5_LC_19_2_6 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_5_LC_19_2_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_5_LC_19_2_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_5_LC_19_2_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47214),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19443_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19443_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_6_LC_19_2_7 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_6_LC_19_2_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_6_LC_19_2_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_6_LC_19_2_7  (
            .in0(_gnd_net_),
            .in1(N__47189),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19443_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19443_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i2_LC_19_3_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i2_LC_19_3_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i2_LC_19_3_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i2_LC_19_3_0  (
            .in0(N__51191),
            .in1(N__56353),
            .in2(_gnd_net_),
            .in3(N__44983),
            .lcout(\c0.FRAME_MATCHER_i_2 ),
            .ltout(),
            .carryin(bfn_19_3_0_),
            .carryout(\c0.n19444 ),
            .clk(N__66632),
            .ce(),
            .sr(N__47413));
    defparam \c0.add_49_4_THRU_CRY_0_LC_19_3_1 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_0_LC_19_3_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_0_LC_19_3_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_0_LC_19_3_1  (
            .in0(_gnd_net_),
            .in1(N__47164),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19444 ),
            .carryout(\c0.n19444_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_1_LC_19_3_2 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_1_LC_19_3_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_1_LC_19_3_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_1_LC_19_3_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47209),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19444_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19444_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_2_LC_19_3_3 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_2_LC_19_3_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_2_LC_19_3_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_2_LC_19_3_3  (
            .in0(_gnd_net_),
            .in1(N__47168),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19444_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19444_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_3_LC_19_3_4 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_3_LC_19_3_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_3_LC_19_3_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_3_LC_19_3_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47210),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19444_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19444_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_4_LC_19_3_5 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_4_LC_19_3_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_4_LC_19_3_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_4_LC_19_3_5  (
            .in0(_gnd_net_),
            .in1(N__47172),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19444_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19444_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_5_LC_19_3_6 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_5_LC_19_3_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_5_LC_19_3_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_5_LC_19_3_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47211),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19444_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19444_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_6_LC_19_3_7 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_6_LC_19_3_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_6_LC_19_3_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_6_LC_19_3_7  (
            .in0(_gnd_net_),
            .in1(N__47176),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19444_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19444_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i3_LC_19_4_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i3_LC_19_4_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i3_LC_19_4_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i3_LC_19_4_0  (
            .in0(N__51160),
            .in1(N__45999),
            .in2(_gnd_net_),
            .in3(N__44986),
            .lcout(\c0.FRAME_MATCHER_i_3 ),
            .ltout(),
            .carryin(bfn_19_4_0_),
            .carryout(\c0.n19445 ),
            .clk(N__66633),
            .ce(),
            .sr(N__45964));
    defparam \c0.add_49_5_THRU_CRY_0_LC_19_4_1 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_0_LC_19_4_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_0_LC_19_4_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_0_LC_19_4_1  (
            .in0(_gnd_net_),
            .in1(N__47151),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19445 ),
            .carryout(\c0.n19445_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_1_LC_19_4_2 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_1_LC_19_4_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_1_LC_19_4_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_1_LC_19_4_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47206),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19445_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19445_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_2_LC_19_4_3 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_2_LC_19_4_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_2_LC_19_4_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_2_LC_19_4_3  (
            .in0(_gnd_net_),
            .in1(N__47155),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19445_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19445_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_3_LC_19_4_4 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_3_LC_19_4_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_3_LC_19_4_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_3_LC_19_4_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47207),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19445_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19445_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_4_LC_19_4_5 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_4_LC_19_4_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_4_LC_19_4_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_4_LC_19_4_5  (
            .in0(_gnd_net_),
            .in1(N__47159),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19445_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19445_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_5_LC_19_4_6 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_5_LC_19_4_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_5_LC_19_4_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_5_LC_19_4_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47208),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19445_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19445_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_6_LC_19_4_7 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_6_LC_19_4_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_6_LC_19_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_6_LC_19_4_7  (
            .in0(_gnd_net_),
            .in1(N__47163),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19445_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19445_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i4_LC_19_5_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i4_LC_19_5_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i4_LC_19_5_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i4_LC_19_5_0  (
            .in0(N__51175),
            .in1(N__45018),
            .in2(_gnd_net_),
            .in3(N__45007),
            .lcout(\c0.FRAME_MATCHER_i_4 ),
            .ltout(),
            .carryin(bfn_19_5_0_),
            .carryout(\c0.n19446 ),
            .clk(N__66635),
            .ce(),
            .sr(N__45004));
    defparam \c0.add_49_6_THRU_CRY_0_LC_19_5_1 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_0_LC_19_5_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_0_LC_19_5_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_0_LC_19_5_1  (
            .in0(_gnd_net_),
            .in1(N__47063),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19446 ),
            .carryout(\c0.n19446_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_1_LC_19_5_2 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_1_LC_19_5_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_1_LC_19_5_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_1_LC_19_5_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47148),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19446_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19446_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_2_LC_19_5_3 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_2_LC_19_5_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_2_LC_19_5_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_2_LC_19_5_3  (
            .in0(_gnd_net_),
            .in1(N__47067),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19446_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19446_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_3_LC_19_5_4 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_3_LC_19_5_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_3_LC_19_5_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_3_LC_19_5_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47149),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19446_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19446_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_4_LC_19_5_5 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_4_LC_19_5_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_4_LC_19_5_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_4_LC_19_5_5  (
            .in0(_gnd_net_),
            .in1(N__47071),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19446_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19446_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_5_LC_19_5_6 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_5_LC_19_5_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_5_LC_19_5_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_5_LC_19_5_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47150),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19446_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19446_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_6_LC_19_5_7 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_6_LC_19_5_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_6_LC_19_5_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_6_LC_19_5_7  (
            .in0(_gnd_net_),
            .in1(N__47075),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19446_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19446_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i5_LC_19_6_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i5_LC_19_6_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i5_LC_19_6_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i5_LC_19_6_0  (
            .in0(N__51174),
            .in1(N__47380),
            .in2(_gnd_net_),
            .in3(N__45100),
            .lcout(\c0.FRAME_MATCHER_i_5 ),
            .ltout(),
            .carryin(bfn_19_6_0_),
            .carryout(\c0.n19447 ),
            .clk(N__66637),
            .ce(),
            .sr(N__45097));
    defparam \c0.add_49_7_THRU_CRY_0_LC_19_6_1 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_0_LC_19_6_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_0_LC_19_6_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_0_LC_19_6_1  (
            .in0(_gnd_net_),
            .in1(N__47050),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19447 ),
            .carryout(\c0.n19447_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_1_LC_19_6_2 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_1_LC_19_6_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_1_LC_19_6_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_1_LC_19_6_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47145),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19447_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19447_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_2_LC_19_6_3 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_2_LC_19_6_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_2_LC_19_6_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_2_LC_19_6_3  (
            .in0(_gnd_net_),
            .in1(N__47054),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19447_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19447_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_3_LC_19_6_4 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_3_LC_19_6_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_3_LC_19_6_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_3_LC_19_6_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47146),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19447_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19447_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_4_LC_19_6_5 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_4_LC_19_6_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_4_LC_19_6_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_4_LC_19_6_5  (
            .in0(_gnd_net_),
            .in1(N__47058),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19447_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19447_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_5_LC_19_6_6 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_5_LC_19_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_5_LC_19_6_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_5_LC_19_6_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47147),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19447_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19447_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_6_LC_19_6_7 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_6_LC_19_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_6_LC_19_6_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_6_LC_19_6_7  (
            .in0(_gnd_net_),
            .in1(N__47062),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19447_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19447_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i6_LC_19_7_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i6_LC_19_7_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i6_LC_19_7_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i6_LC_19_7_0  (
            .in0(N__51172),
            .in1(N__47348),
            .in2(_gnd_net_),
            .in3(N__45118),
            .lcout(\c0.FRAME_MATCHER_i_6 ),
            .ltout(),
            .carryin(bfn_19_7_0_),
            .carryout(\c0.n19448 ),
            .clk(N__66642),
            .ce(),
            .sr(N__45115));
    defparam \c0.add_49_8_THRU_CRY_0_LC_19_7_1 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_0_LC_19_7_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_0_LC_19_7_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_0_LC_19_7_1  (
            .in0(_gnd_net_),
            .in1(N__47037),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19448 ),
            .carryout(\c0.n19448_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_1_LC_19_7_2 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_1_LC_19_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_1_LC_19_7_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_1_LC_19_7_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47142),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19448_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19448_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_2_LC_19_7_3 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_2_LC_19_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_2_LC_19_7_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_2_LC_19_7_3  (
            .in0(_gnd_net_),
            .in1(N__47041),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19448_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19448_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_3_LC_19_7_4 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_3_LC_19_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_3_LC_19_7_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_3_LC_19_7_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47143),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19448_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19448_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_4_LC_19_7_5 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_4_LC_19_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_4_LC_19_7_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_4_LC_19_7_5  (
            .in0(_gnd_net_),
            .in1(N__47045),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19448_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19448_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_5_LC_19_7_6 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_5_LC_19_7_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_5_LC_19_7_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_5_LC_19_7_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47144),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19448_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19448_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_6_LC_19_7_7 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_6_LC_19_7_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_6_LC_19_7_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_6_LC_19_7_7  (
            .in0(_gnd_net_),
            .in1(N__47049),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19448_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19448_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i7_LC_19_8_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i7_LC_19_8_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i7_LC_19_8_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i7_LC_19_8_0  (
            .in0(N__51064),
            .in1(N__45155),
            .in2(_gnd_net_),
            .in3(N__45139),
            .lcout(\c0.FRAME_MATCHER_i_7 ),
            .ltout(),
            .carryin(bfn_19_8_0_),
            .carryout(\c0.n19449 ),
            .clk(N__66649),
            .ce(),
            .sr(N__45136));
    defparam \c0.add_49_9_THRU_CRY_0_LC_19_8_1 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_0_LC_19_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_0_LC_19_8_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_0_LC_19_8_1  (
            .in0(_gnd_net_),
            .in1(N__47024),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19449 ),
            .carryout(\c0.n19449_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_1_LC_19_8_2 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_1_LC_19_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_1_LC_19_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_1_LC_19_8_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47139),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19449_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19449_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_2_LC_19_8_3 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_2_LC_19_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_2_LC_19_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_2_LC_19_8_3  (
            .in0(_gnd_net_),
            .in1(N__47028),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19449_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19449_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_3_LC_19_8_4 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_3_LC_19_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_3_LC_19_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_3_LC_19_8_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47140),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19449_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19449_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_4_LC_19_8_5 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_4_LC_19_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_4_LC_19_8_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_4_LC_19_8_5  (
            .in0(_gnd_net_),
            .in1(N__47032),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19449_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19449_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_5_LC_19_8_6 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_5_LC_19_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_5_LC_19_8_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_5_LC_19_8_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47141),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19449_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19449_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_6_LC_19_8_7 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_6_LC_19_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_6_LC_19_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_6_LC_19_8_7  (
            .in0(_gnd_net_),
            .in1(N__47036),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19449_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19449_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i8_LC_19_9_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i8_LC_19_9_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i8_LC_19_9_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i8_LC_19_9_0  (
            .in0(N__51193),
            .in1(N__45215),
            .in2(_gnd_net_),
            .in3(N__45196),
            .lcout(\c0.FRAME_MATCHER_i_8 ),
            .ltout(),
            .carryin(bfn_19_9_0_),
            .carryout(\c0.n19450 ),
            .clk(N__66656),
            .ce(),
            .sr(N__45193));
    defparam \c0.add_49_10_THRU_CRY_0_LC_19_9_1 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_0_LC_19_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_0_LC_19_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_0_LC_19_9_1  (
            .in0(_gnd_net_),
            .in1(N__46927),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19450 ),
            .carryout(\c0.n19450_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_1_LC_19_9_2 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_1_LC_19_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_1_LC_19_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_1_LC_19_9_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47021),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19450_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19450_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_2_LC_19_9_3 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_2_LC_19_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_2_LC_19_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_2_LC_19_9_3  (
            .in0(_gnd_net_),
            .in1(N__46931),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19450_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19450_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_3_LC_19_9_4 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_3_LC_19_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_3_LC_19_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_3_LC_19_9_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47022),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19450_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19450_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_4_LC_19_9_5 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_4_LC_19_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_4_LC_19_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_4_LC_19_9_5  (
            .in0(_gnd_net_),
            .in1(N__46935),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19450_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19450_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_5_LC_19_9_6 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_5_LC_19_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_5_LC_19_9_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_5_LC_19_9_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47023),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19450_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19450_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_6_LC_19_9_7 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_6_LC_19_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_6_LC_19_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_6_LC_19_9_7  (
            .in0(_gnd_net_),
            .in1(N__46939),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19450_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19450_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i9_LC_19_10_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i9_LC_19_10_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i9_LC_19_10_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i9_LC_19_10_0  (
            .in0(N__51192),
            .in1(N__45266),
            .in2(_gnd_net_),
            .in3(N__45250),
            .lcout(\c0.FRAME_MATCHER_i_9 ),
            .ltout(),
            .carryin(bfn_19_10_0_),
            .carryout(\c0.n19451 ),
            .clk(N__66661),
            .ce(),
            .sr(N__45247));
    defparam \c0.add_49_11_THRU_CRY_0_LC_19_10_1 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_0_LC_19_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_0_LC_19_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_0_LC_19_10_1  (
            .in0(_gnd_net_),
            .in1(N__46914),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19451 ),
            .carryout(\c0.n19451_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_1_LC_19_10_2 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_1_LC_19_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_1_LC_19_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_1_LC_19_10_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47018),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19451_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19451_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_2_LC_19_10_3 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_2_LC_19_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_2_LC_19_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_2_LC_19_10_3  (
            .in0(_gnd_net_),
            .in1(N__46918),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19451_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19451_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_3_LC_19_10_4 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_3_LC_19_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_3_LC_19_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_3_LC_19_10_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47019),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19451_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19451_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_4_LC_19_10_5 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_4_LC_19_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_4_LC_19_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_4_LC_19_10_5  (
            .in0(_gnd_net_),
            .in1(N__46922),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19451_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19451_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_5_LC_19_10_6 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_5_LC_19_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_5_LC_19_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_5_LC_19_10_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47020),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19451_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19451_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_6_LC_19_10_7 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_6_LC_19_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_6_LC_19_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_6_LC_19_10_7  (
            .in0(_gnd_net_),
            .in1(N__46926),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19451_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19451_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i10_LC_19_11_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i10_LC_19_11_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i10_LC_19_11_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i10_LC_19_11_0  (
            .in0(N__51204),
            .in1(N__50138),
            .in2(_gnd_net_),
            .in3(N__45232),
            .lcout(\c0.FRAME_MATCHER_i_10 ),
            .ltout(),
            .carryin(bfn_19_11_0_),
            .carryout(\c0.n19452 ),
            .clk(N__66667),
            .ce(),
            .sr(N__50122));
    defparam \c0.add_49_12_THRU_CRY_0_LC_19_11_1 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_0_LC_19_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_0_LC_19_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_0_LC_19_11_1  (
            .in0(_gnd_net_),
            .in1(N__46901),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19452 ),
            .carryout(\c0.n19452_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_1_LC_19_11_2 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_1_LC_19_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_1_LC_19_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_1_LC_19_11_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47015),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19452_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19452_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_2_LC_19_11_3 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_2_LC_19_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_2_LC_19_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_2_LC_19_11_3  (
            .in0(_gnd_net_),
            .in1(N__46905),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19452_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19452_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_3_LC_19_11_4 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_3_LC_19_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_3_LC_19_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_3_LC_19_11_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47016),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19452_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19452_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_4_LC_19_11_5 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_4_LC_19_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_4_LC_19_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_4_LC_19_11_5  (
            .in0(_gnd_net_),
            .in1(N__46909),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19452_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19452_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_5_LC_19_11_6 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_5_LC_19_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_5_LC_19_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_5_LC_19_11_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47017),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19452_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19452_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_6_LC_19_11_7 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_6_LC_19_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_6_LC_19_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_6_LC_19_11_7  (
            .in0(_gnd_net_),
            .in1(N__46913),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19452_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19452_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i11_LC_19_12_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i11_LC_19_12_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i11_LC_19_12_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i11_LC_19_12_0  (
            .in0(N__51203),
            .in1(N__45314),
            .in2(_gnd_net_),
            .in3(N__45301),
            .lcout(\c0.FRAME_MATCHER_i_11 ),
            .ltout(),
            .carryin(bfn_19_12_0_),
            .carryout(\c0.n19453 ),
            .clk(N__66678),
            .ce(),
            .sr(N__45298));
    defparam \c0.add_49_13_THRU_CRY_0_LC_19_12_1 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_0_LC_19_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_0_LC_19_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_0_LC_19_12_1  (
            .in0(_gnd_net_),
            .in1(N__46888),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19453 ),
            .carryout(\c0.n19453_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_1_LC_19_12_2 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_1_LC_19_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_1_LC_19_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_1_LC_19_12_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47012),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19453_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19453_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_2_LC_19_12_3 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_2_LC_19_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_2_LC_19_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_2_LC_19_12_3  (
            .in0(_gnd_net_),
            .in1(N__46892),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19453_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19453_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_3_LC_19_12_4 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_3_LC_19_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_3_LC_19_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_3_LC_19_12_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47013),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19453_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19453_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_4_LC_19_12_5 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_4_LC_19_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_4_LC_19_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_4_LC_19_12_5  (
            .in0(_gnd_net_),
            .in1(N__46896),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19453_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19453_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_5_LC_19_12_6 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_5_LC_19_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_5_LC_19_12_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_5_LC_19_12_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__47014),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19453_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19453_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_6_LC_19_12_7 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_6_LC_19_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_6_LC_19_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_6_LC_19_12_7  (
            .in0(_gnd_net_),
            .in1(N__46900),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19453_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19453_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i12_LC_19_13_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i12_LC_19_13_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i12_LC_19_13_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i12_LC_19_13_0  (
            .in0(N__51205),
            .in1(N__45362),
            .in2(_gnd_net_),
            .in3(N__45346),
            .lcout(\c0.FRAME_MATCHER_i_12 ),
            .ltout(),
            .carryin(bfn_19_13_0_),
            .carryout(\c0.n19454 ),
            .clk(N__66690),
            .ce(),
            .sr(N__45343));
    defparam \c0.add_49_14_THRU_CRY_0_LC_19_13_1 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_0_LC_19_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_0_LC_19_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_0_LC_19_13_1  (
            .in0(_gnd_net_),
            .in1(N__46789),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19454 ),
            .carryout(\c0.n19454_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_1_LC_19_13_2 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_1_LC_19_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_1_LC_19_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_1_LC_19_13_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46885),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19454_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19454_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_2_LC_19_13_3 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_2_LC_19_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_2_LC_19_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_2_LC_19_13_3  (
            .in0(_gnd_net_),
            .in1(N__46793),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19454_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19454_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_3_LC_19_13_4 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_3_LC_19_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_3_LC_19_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_3_LC_19_13_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46886),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19454_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19454_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_4_LC_19_13_5 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_4_LC_19_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_4_LC_19_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_4_LC_19_13_5  (
            .in0(_gnd_net_),
            .in1(N__46797),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19454_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19454_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_5_LC_19_13_6 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_5_LC_19_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_5_LC_19_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_5_LC_19_13_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46887),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19454_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19454_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_6_LC_19_13_7 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_6_LC_19_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_6_LC_19_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_6_LC_19_13_7  (
            .in0(_gnd_net_),
            .in1(N__46801),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19454_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19454_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i13_LC_19_14_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i13_LC_19_14_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i13_LC_19_14_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i13_LC_19_14_0  (
            .in0(N__51113),
            .in1(N__49851),
            .in2(_gnd_net_),
            .in3(N__45388),
            .lcout(\c0.FRAME_MATCHER_i_13 ),
            .ltout(),
            .carryin(bfn_19_14_0_),
            .carryout(\c0.n19455 ),
            .clk(N__66704),
            .ce(),
            .sr(N__49837));
    defparam \c0.add_49_15_THRU_CRY_0_LC_19_14_1 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_0_LC_19_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_0_LC_19_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_0_LC_19_14_1  (
            .in0(_gnd_net_),
            .in1(N__46776),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19455 ),
            .carryout(\c0.n19455_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_1_LC_19_14_2 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_1_LC_19_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_1_LC_19_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_1_LC_19_14_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46882),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19455_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19455_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_2_LC_19_14_3 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_2_LC_19_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_2_LC_19_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_2_LC_19_14_3  (
            .in0(_gnd_net_),
            .in1(N__46780),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19455_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19455_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_3_LC_19_14_4 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_3_LC_19_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_3_LC_19_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_3_LC_19_14_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46883),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19455_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19455_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_4_LC_19_14_5 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_4_LC_19_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_4_LC_19_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_4_LC_19_14_5  (
            .in0(_gnd_net_),
            .in1(N__46784),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19455_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19455_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_5_LC_19_14_6 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_5_LC_19_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_5_LC_19_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_5_LC_19_14_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46884),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19455_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19455_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_6_LC_19_14_7 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_6_LC_19_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_6_LC_19_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_6_LC_19_14_7  (
            .in0(_gnd_net_),
            .in1(N__46788),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19455_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19455_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i14_LC_19_15_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i14_LC_19_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i14_LC_19_15_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i14_LC_19_15_0  (
            .in0(N__51097),
            .in1(N__45425),
            .in2(_gnd_net_),
            .in3(N__45406),
            .lcout(\c0.FRAME_MATCHER_i_14 ),
            .ltout(),
            .carryin(bfn_19_15_0_),
            .carryout(\c0.n19456 ),
            .clk(N__66718),
            .ce(),
            .sr(N__45403));
    defparam \c0.add_49_16_THRU_CRY_0_LC_19_15_1 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_0_LC_19_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_0_LC_19_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_0_LC_19_15_1  (
            .in0(_gnd_net_),
            .in1(N__46763),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19456 ),
            .carryout(\c0.n19456_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_1_LC_19_15_2 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_1_LC_19_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_1_LC_19_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_1_LC_19_15_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46879),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19456_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19456_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_2_LC_19_15_3 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_2_LC_19_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_2_LC_19_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_2_LC_19_15_3  (
            .in0(_gnd_net_),
            .in1(N__46767),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19456_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19456_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_3_LC_19_15_4 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_3_LC_19_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_3_LC_19_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_3_LC_19_15_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46880),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19456_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19456_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_4_LC_19_15_5 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_4_LC_19_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_4_LC_19_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_4_LC_19_15_5  (
            .in0(_gnd_net_),
            .in1(N__46771),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19456_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19456_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_5_LC_19_15_6 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_5_LC_19_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_5_LC_19_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_5_LC_19_15_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46881),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19456_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19456_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_6_LC_19_15_7 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_6_LC_19_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_6_LC_19_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_6_LC_19_15_7  (
            .in0(_gnd_net_),
            .in1(N__46775),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19456_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19456_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i15_LC_19_16_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i15_LC_19_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i15_LC_19_16_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i15_LC_19_16_0  (
            .in0(N__51112),
            .in1(N__49814),
            .in2(_gnd_net_),
            .in3(N__45442),
            .lcout(\c0.FRAME_MATCHER_i_15 ),
            .ltout(),
            .carryin(bfn_19_16_0_),
            .carryout(\c0.n19457 ),
            .clk(N__66732),
            .ce(),
            .sr(N__49795));
    defparam \c0.add_49_17_THRU_CRY_0_LC_19_16_1 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_0_LC_19_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_0_LC_19_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_0_LC_19_16_1  (
            .in0(_gnd_net_),
            .in1(N__46750),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19457 ),
            .carryout(\c0.n19457_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_1_LC_19_16_2 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_1_LC_19_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_1_LC_19_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_1_LC_19_16_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46876),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19457_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19457_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_2_LC_19_16_3 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_2_LC_19_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_2_LC_19_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_2_LC_19_16_3  (
            .in0(_gnd_net_),
            .in1(N__46754),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19457_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19457_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_3_LC_19_16_4 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_3_LC_19_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_3_LC_19_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_3_LC_19_16_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46877),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19457_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19457_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_4_LC_19_16_5 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_4_LC_19_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_4_LC_19_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_4_LC_19_16_5  (
            .in0(_gnd_net_),
            .in1(N__46758),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19457_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19457_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_5_LC_19_16_6 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_5_LC_19_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_5_LC_19_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_5_LC_19_16_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46878),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19457_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19457_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_6_LC_19_16_7 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_6_LC_19_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_6_LC_19_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_6_LC_19_16_7  (
            .in0(_gnd_net_),
            .in1(N__46762),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19457_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19457_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i16_LC_19_17_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i16_LC_19_17_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i16_LC_19_17_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i16_LC_19_17_0  (
            .in0(N__50955),
            .in1(N__49889),
            .in2(_gnd_net_),
            .in3(N__45454),
            .lcout(\c0.FRAME_MATCHER_i_16 ),
            .ltout(),
            .carryin(bfn_19_17_0_),
            .carryout(\c0.n19458 ),
            .clk(N__66746),
            .ce(),
            .sr(N__45451));
    defparam \c0.add_49_18_THRU_CRY_0_LC_19_17_1 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_0_LC_19_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_0_LC_19_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_0_LC_19_17_1  (
            .in0(_gnd_net_),
            .in1(N__46654),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19458 ),
            .carryout(\c0.n19458_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_1_LC_19_17_2 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_1_LC_19_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_1_LC_19_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_1_LC_19_17_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46747),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19458_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19458_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_2_LC_19_17_3 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_2_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_2_LC_19_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_2_LC_19_17_3  (
            .in0(_gnd_net_),
            .in1(N__46658),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19458_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19458_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_3_LC_19_17_4 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_3_LC_19_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_3_LC_19_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_3_LC_19_17_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46748),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19458_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19458_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_4_LC_19_17_5 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_4_LC_19_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_4_LC_19_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_4_LC_19_17_5  (
            .in0(_gnd_net_),
            .in1(N__46662),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19458_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19458_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_5_LC_19_17_6 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_5_LC_19_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_5_LC_19_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_5_LC_19_17_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46749),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19458_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19458_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_6_LC_19_17_7 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_6_LC_19_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_6_LC_19_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_6_LC_19_17_7  (
            .in0(_gnd_net_),
            .in1(N__46666),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19458_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19458_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i17_LC_19_18_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i17_LC_19_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i17_LC_19_18_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i17_LC_19_18_0  (
            .in0(N__51054),
            .in1(N__45491),
            .in2(_gnd_net_),
            .in3(N__45472),
            .lcout(\c0.FRAME_MATCHER_i_17 ),
            .ltout(),
            .carryin(bfn_19_18_0_),
            .carryout(\c0.n19459 ),
            .clk(N__66760),
            .ce(),
            .sr(N__45469));
    defparam \c0.add_49_19_THRU_CRY_0_LC_19_18_1 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_0_LC_19_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_0_LC_19_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_0_LC_19_18_1  (
            .in0(_gnd_net_),
            .in1(N__46641),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19459 ),
            .carryout(\c0.n19459_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_1_LC_19_18_2 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_1_LC_19_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_1_LC_19_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_1_LC_19_18_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46744),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19459_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19459_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_2_LC_19_18_3 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_2_LC_19_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_2_LC_19_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_2_LC_19_18_3  (
            .in0(_gnd_net_),
            .in1(N__46645),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19459_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19459_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_3_LC_19_18_4 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_3_LC_19_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_3_LC_19_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_3_LC_19_18_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46745),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19459_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19459_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_4_LC_19_18_5 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_4_LC_19_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_4_LC_19_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_4_LC_19_18_5  (
            .in0(_gnd_net_),
            .in1(N__46649),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19459_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19459_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_5_LC_19_18_6 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_5_LC_19_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_5_LC_19_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_5_LC_19_18_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46746),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19459_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19459_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_6_LC_19_18_7 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_6_LC_19_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_6_LC_19_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_6_LC_19_18_7  (
            .in0(_gnd_net_),
            .in1(N__46653),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19459_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19459_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i18_LC_19_19_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i18_LC_19_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i18_LC_19_19_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i18_LC_19_19_0  (
            .in0(N__51053),
            .in1(N__45569),
            .in2(_gnd_net_),
            .in3(N__45550),
            .lcout(\c0.FRAME_MATCHER_i_18 ),
            .ltout(),
            .carryin(bfn_19_19_0_),
            .carryout(\c0.n19460 ),
            .clk(N__66772),
            .ce(),
            .sr(N__45547));
    defparam \c0.add_49_20_THRU_CRY_0_LC_19_19_1 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_0_LC_19_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_0_LC_19_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_0_LC_19_19_1  (
            .in0(_gnd_net_),
            .in1(N__46628),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19460 ),
            .carryout(\c0.n19460_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_1_LC_19_19_2 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_1_LC_19_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_1_LC_19_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_1_LC_19_19_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46741),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19460_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19460_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_2_LC_19_19_3 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_2_LC_19_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_2_LC_19_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_2_LC_19_19_3  (
            .in0(_gnd_net_),
            .in1(N__46632),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19460_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19460_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_3_LC_19_19_4 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_3_LC_19_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_3_LC_19_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_3_LC_19_19_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46742),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19460_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19460_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_4_LC_19_19_5 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_4_LC_19_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_4_LC_19_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_4_LC_19_19_5  (
            .in0(_gnd_net_),
            .in1(N__46636),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19460_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19460_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_5_LC_19_19_6 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_5_LC_19_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_5_LC_19_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_5_LC_19_19_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46743),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19460_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19460_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_6_LC_19_19_7 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_6_LC_19_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_6_LC_19_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_6_LC_19_19_7  (
            .in0(_gnd_net_),
            .in1(N__46640),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19460_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19460_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i19_LC_19_20_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i19_LC_19_20_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i19_LC_19_20_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i19_LC_19_20_0  (
            .in0(N__51052),
            .in1(N__45524),
            .in2(_gnd_net_),
            .in3(N__45505),
            .lcout(\c0.FRAME_MATCHER_i_19 ),
            .ltout(),
            .carryin(bfn_19_20_0_),
            .carryout(\c0.n19461 ),
            .clk(N__66786),
            .ce(),
            .sr(N__45601));
    defparam \c0.add_49_21_THRU_CRY_0_LC_19_20_1 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_0_LC_19_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_0_LC_19_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_0_LC_19_20_1  (
            .in0(_gnd_net_),
            .in1(N__46495),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19461 ),
            .carryout(\c0.n19461_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_1_LC_19_20_2 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_1_LC_19_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_1_LC_19_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_1_LC_19_20_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46619),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19461_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19461_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_2_LC_19_20_3 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_2_LC_19_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_2_LC_19_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_2_LC_19_20_3  (
            .in0(_gnd_net_),
            .in1(N__46499),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19461_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19461_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_3_LC_19_20_4 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_3_LC_19_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_3_LC_19_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_3_LC_19_20_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46620),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19461_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19461_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_4_LC_19_20_5 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_4_LC_19_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_4_LC_19_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_4_LC_19_20_5  (
            .in0(_gnd_net_),
            .in1(N__46503),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19461_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19461_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_5_LC_19_20_6 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_5_LC_19_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_5_LC_19_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_5_LC_19_20_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46621),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19461_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19461_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_6_LC_19_20_7 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_6_LC_19_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_6_LC_19_20_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_6_LC_19_20_7  (
            .in0(_gnd_net_),
            .in1(N__46507),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19461_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19461_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i20_LC_19_21_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i20_LC_19_21_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i20_LC_19_21_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i20_LC_19_21_0  (
            .in0(N__51055),
            .in1(N__49992),
            .in2(_gnd_net_),
            .in3(N__45586),
            .lcout(\c0.FRAME_MATCHER_i_20 ),
            .ltout(),
            .carryin(bfn_19_21_0_),
            .carryout(\c0.n19462 ),
            .clk(N__66797),
            .ce(),
            .sr(N__49981));
    defparam \c0.add_49_22_THRU_CRY_0_LC_19_21_1 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_0_LC_19_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_0_LC_19_21_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_0_LC_19_21_1  (
            .in0(_gnd_net_),
            .in1(N__46545),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19462 ),
            .carryout(\c0.n19462_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_1_LC_19_21_2 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_1_LC_19_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_1_LC_19_21_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_1_LC_19_21_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46625),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19462_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19462_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_2_LC_19_21_3 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_2_LC_19_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_2_LC_19_21_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_2_LC_19_21_3  (
            .in0(_gnd_net_),
            .in1(N__46549),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19462_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19462_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_3_LC_19_21_4 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_3_LC_19_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_3_LC_19_21_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_3_LC_19_21_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46626),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19462_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19462_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_4_LC_19_21_5 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_4_LC_19_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_4_LC_19_21_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_4_LC_19_21_5  (
            .in0(_gnd_net_),
            .in1(N__46553),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19462_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19462_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_5_LC_19_21_6 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_5_LC_19_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_5_LC_19_21_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_5_LC_19_21_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46627),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19462_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19462_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_6_LC_19_21_7 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_6_LC_19_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_6_LC_19_21_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_6_LC_19_21_7  (
            .in0(_gnd_net_),
            .in1(N__46557),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19462_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19462_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i21_LC_19_22_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i21_LC_19_22_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i21_LC_19_22_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i21_LC_19_22_0  (
            .in0(N__51010),
            .in1(N__45629),
            .in2(_gnd_net_),
            .in3(N__45613),
            .lcout(\c0.FRAME_MATCHER_i_21 ),
            .ltout(),
            .carryin(bfn_19_22_0_),
            .carryout(\c0.n19463 ),
            .clk(N__66806),
            .ce(),
            .sr(N__45610));
    defparam \c0.add_49_23_THRU_CRY_0_LC_19_22_1 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_0_LC_19_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_0_LC_19_22_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_0_LC_19_22_1  (
            .in0(_gnd_net_),
            .in1(N__46532),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19463 ),
            .carryout(\c0.n19463_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_1_LC_19_22_2 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_1_LC_19_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_1_LC_19_22_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_1_LC_19_22_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46622),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19463_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19463_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_2_LC_19_22_3 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_2_LC_19_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_2_LC_19_22_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_2_LC_19_22_3  (
            .in0(_gnd_net_),
            .in1(N__46536),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19463_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19463_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_3_LC_19_22_4 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_3_LC_19_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_3_LC_19_22_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_3_LC_19_22_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46623),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19463_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19463_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_4_LC_19_22_5 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_4_LC_19_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_4_LC_19_22_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_4_LC_19_22_5  (
            .in0(_gnd_net_),
            .in1(N__46540),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19463_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19463_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_5_LC_19_22_6 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_5_LC_19_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_5_LC_19_22_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_5_LC_19_22_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46624),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19463_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19463_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_6_LC_19_22_7 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_6_LC_19_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_6_LC_19_22_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_6_LC_19_22_7  (
            .in0(_gnd_net_),
            .in1(N__46544),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19463_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19463_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i22_LC_19_23_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i22_LC_19_23_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i22_LC_19_23_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i22_LC_19_23_0  (
            .in0(N__51088),
            .in1(N__45674),
            .in2(_gnd_net_),
            .in3(N__45655),
            .lcout(\c0.FRAME_MATCHER_i_22 ),
            .ltout(),
            .carryin(bfn_19_23_0_),
            .carryout(\c0.n19464 ),
            .clk(N__66818),
            .ce(),
            .sr(N__45652));
    defparam \c0.add_49_24_THRU_CRY_0_LC_19_23_1 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_0_LC_19_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_0_LC_19_23_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_0_LC_19_23_1  (
            .in0(_gnd_net_),
            .in1(N__46479),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19464 ),
            .carryout(\c0.n19464_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_1_LC_19_23_2 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_1_LC_19_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_1_LC_19_23_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_1_LC_19_23_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46616),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19464_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19464_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_2_LC_19_23_3 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_2_LC_19_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_2_LC_19_23_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_2_LC_19_23_3  (
            .in0(_gnd_net_),
            .in1(N__46483),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19464_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19464_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_3_LC_19_23_4 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_3_LC_19_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_3_LC_19_23_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_3_LC_19_23_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46617),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19464_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19464_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_4_LC_19_23_5 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_4_LC_19_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_4_LC_19_23_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_4_LC_19_23_5  (
            .in0(_gnd_net_),
            .in1(N__46487),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19464_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19464_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_5_LC_19_23_6 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_5_LC_19_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_5_LC_19_23_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_5_LC_19_23_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46618),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19464_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19464_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_6_LC_19_23_7 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_6_LC_19_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_6_LC_19_23_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_6_LC_19_23_7  (
            .in0(_gnd_net_),
            .in1(N__46491),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19464_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19464_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i23_LC_19_24_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i23_LC_19_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i23_LC_19_24_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i23_LC_19_24_0  (
            .in0(N__51087),
            .in1(N__45707),
            .in2(_gnd_net_),
            .in3(N__45688),
            .lcout(\c0.FRAME_MATCHER_i_23 ),
            .ltout(),
            .carryin(bfn_19_24_0_),
            .carryout(\c0.n19465 ),
            .clk(N__66830),
            .ce(),
            .sr(N__45685));
    defparam \c0.add_49_25_THRU_CRY_0_LC_19_24_1 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_0_LC_19_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_0_LC_19_24_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_0_LC_19_24_1  (
            .in0(_gnd_net_),
            .in1(N__46351),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19465 ),
            .carryout(\c0.n19465_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_1_LC_19_24_2 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_1_LC_19_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_1_LC_19_24_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_1_LC_19_24_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46492),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19465_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19465_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_2_LC_19_24_3 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_2_LC_19_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_2_LC_19_24_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_2_LC_19_24_3  (
            .in0(_gnd_net_),
            .in1(N__46355),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19465_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19465_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_3_LC_19_24_4 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_3_LC_19_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_3_LC_19_24_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_3_LC_19_24_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46493),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19465_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19465_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_4_LC_19_24_5 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_4_LC_19_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_4_LC_19_24_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_4_LC_19_24_5  (
            .in0(_gnd_net_),
            .in1(N__46359),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19465_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19465_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_5_LC_19_24_6 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_5_LC_19_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_5_LC_19_24_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_5_LC_19_24_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46494),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19465_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19465_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_6_LC_19_24_7 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_6_LC_19_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_6_LC_19_24_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_6_LC_19_24_7  (
            .in0(_gnd_net_),
            .in1(N__46363),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19465_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19465_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i24_LC_19_25_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i24_LC_19_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i24_LC_19_25_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i24_LC_19_25_0  (
            .in0(N__51085),
            .in1(N__45749),
            .in2(_gnd_net_),
            .in3(N__45730),
            .lcout(\c0.FRAME_MATCHER_i_24 ),
            .ltout(),
            .carryin(bfn_19_25_0_),
            .carryout(\c0.n19466 ),
            .clk(N__66842),
            .ce(),
            .sr(N__45727));
    defparam \c0.add_49_26_THRU_CRY_0_LC_19_25_1 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_0_LC_19_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_0_LC_19_25_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_0_LC_19_25_1  (
            .in0(_gnd_net_),
            .in1(N__46269),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19466 ),
            .carryout(\c0.n19466_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_1_LC_19_25_2 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_1_LC_19_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_1_LC_19_25_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_1_LC_19_25_2  (
            .in0(_gnd_net_),
            .in1(N__46273),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19466_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19466_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_2_LC_19_25_3 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_2_LC_19_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_2_LC_19_25_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_2_LC_19_25_3  (
            .in0(_gnd_net_),
            .in1(N__46270),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19466_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19466_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_3_LC_19_25_4 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_3_LC_19_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_3_LC_19_25_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_3_LC_19_25_4  (
            .in0(_gnd_net_),
            .in1(N__46274),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19466_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19466_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_4_LC_19_25_5 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_4_LC_19_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_4_LC_19_25_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_4_LC_19_25_5  (
            .in0(_gnd_net_),
            .in1(N__46271),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19466_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19466_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_5_LC_19_25_6 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_5_LC_19_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_5_LC_19_25_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_5_LC_19_25_6  (
            .in0(_gnd_net_),
            .in1(N__46275),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19466_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19466_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_6_LC_19_25_7 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_6_LC_19_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_6_LC_19_25_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_6_LC_19_25_7  (
            .in0(_gnd_net_),
            .in1(N__46272),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19466_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19466_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i25_LC_19_26_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i25_LC_19_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i25_LC_19_26_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i25_LC_19_26_0  (
            .in0(N__51086),
            .in1(N__45791),
            .in2(_gnd_net_),
            .in3(N__45772),
            .lcout(\c0.FRAME_MATCHER_i_25 ),
            .ltout(),
            .carryin(bfn_19_26_0_),
            .carryout(\c0.n19467 ),
            .clk(N__66851),
            .ce(),
            .sr(N__45769));
    defparam \c0.add_49_27_THRU_CRY_0_LC_19_26_1 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_0_LC_19_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_0_LC_19_26_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_0_LC_19_26_1  (
            .in0(_gnd_net_),
            .in1(N__46262),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19467 ),
            .carryout(\c0.n19467_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_1_LC_19_26_2 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_1_LC_19_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_1_LC_19_26_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_1_LC_19_26_2  (
            .in0(_gnd_net_),
            .in1(N__46266),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19467_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19467_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_2_LC_19_26_3 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_2_LC_19_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_2_LC_19_26_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_2_LC_19_26_3  (
            .in0(_gnd_net_),
            .in1(N__46263),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19467_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19467_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_3_LC_19_26_4 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_3_LC_19_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_3_LC_19_26_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_3_LC_19_26_4  (
            .in0(_gnd_net_),
            .in1(N__46267),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19467_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19467_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_4_LC_19_26_5 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_4_LC_19_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_4_LC_19_26_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_4_LC_19_26_5  (
            .in0(_gnd_net_),
            .in1(N__46264),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19467_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19467_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_5_LC_19_26_6 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_5_LC_19_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_5_LC_19_26_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_5_LC_19_26_6  (
            .in0(_gnd_net_),
            .in1(N__46268),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19467_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19467_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_6_LC_19_26_7 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_6_LC_19_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_6_LC_19_26_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_6_LC_19_26_7  (
            .in0(_gnd_net_),
            .in1(N__46265),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19467_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19467_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i26_LC_19_27_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i26_LC_19_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i26_LC_19_27_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i26_LC_19_27_0  (
            .in0(N__51099),
            .in1(N__45830),
            .in2(_gnd_net_),
            .in3(N__45811),
            .lcout(\c0.FRAME_MATCHER_i_26 ),
            .ltout(),
            .carryin(bfn_19_27_0_),
            .carryout(\c0.n19468 ),
            .clk(N__66860),
            .ce(),
            .sr(N__45808));
    defparam \c0.add_49_28_THRU_CRY_0_LC_19_27_1 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_0_LC_19_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_0_LC_19_27_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_0_LC_19_27_1  (
            .in0(_gnd_net_),
            .in1(N__46276),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19468 ),
            .carryout(\c0.n19468_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_1_LC_19_27_2 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_1_LC_19_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_1_LC_19_27_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_1_LC_19_27_2  (
            .in0(_gnd_net_),
            .in1(N__46280),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19468_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19468_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_2_LC_19_27_3 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_2_LC_19_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_2_LC_19_27_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_2_LC_19_27_3  (
            .in0(_gnd_net_),
            .in1(N__46277),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19468_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19468_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_3_LC_19_27_4 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_3_LC_19_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_3_LC_19_27_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_3_LC_19_27_4  (
            .in0(_gnd_net_),
            .in1(N__46281),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19468_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19468_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_4_LC_19_27_5 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_4_LC_19_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_4_LC_19_27_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_4_LC_19_27_5  (
            .in0(_gnd_net_),
            .in1(N__46278),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19468_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19468_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_5_LC_19_27_6 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_5_LC_19_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_5_LC_19_27_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_5_LC_19_27_6  (
            .in0(_gnd_net_),
            .in1(N__46282),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19468_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19468_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_6_LC_19_27_7 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_6_LC_19_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_6_LC_19_27_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_6_LC_19_27_7  (
            .in0(_gnd_net_),
            .in1(N__46279),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19468_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19468_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i27_LC_19_28_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i27_LC_19_28_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i27_LC_19_28_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i27_LC_19_28_0  (
            .in0(N__51130),
            .in1(N__45869),
            .in2(_gnd_net_),
            .in3(N__45850),
            .lcout(\c0.FRAME_MATCHER_i_27 ),
            .ltout(),
            .carryin(bfn_19_28_0_),
            .carryout(\c0.n19469 ),
            .clk(N__66866),
            .ce(),
            .sr(N__45847));
    defparam \c0.add_49_29_THRU_CRY_0_LC_19_28_1 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_0_LC_19_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_0_LC_19_28_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_0_LC_19_28_1  (
            .in0(_gnd_net_),
            .in1(N__46379),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19469 ),
            .carryout(\c0.n19469_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_1_LC_19_28_2 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_1_LC_19_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_1_LC_19_28_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_1_LC_19_28_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46508),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19469_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19469_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_2_LC_19_28_3 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_2_LC_19_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_2_LC_19_28_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_2_LC_19_28_3  (
            .in0(_gnd_net_),
            .in1(N__46383),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19469_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19469_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_3_LC_19_28_4 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_3_LC_19_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_3_LC_19_28_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_3_LC_19_28_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46509),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19469_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19469_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_4_LC_19_28_5 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_4_LC_19_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_4_LC_19_28_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_4_LC_19_28_5  (
            .in0(_gnd_net_),
            .in1(N__46387),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19469_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19469_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_5_LC_19_28_6 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_5_LC_19_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_5_LC_19_28_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_5_LC_19_28_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__46510),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19469_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19469_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_6_LC_19_28_7 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_6_LC_19_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_6_LC_19_28_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_6_LC_19_28_7  (
            .in0(_gnd_net_),
            .in1(N__46391),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19469_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19469_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i28_LC_19_29_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i28_LC_19_29_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i28_LC_19_29_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i28_LC_19_29_0  (
            .in0(N__51123),
            .in1(N__50699),
            .in2(_gnd_net_),
            .in3(N__45907),
            .lcout(\c0.FRAME_MATCHER_i_28 ),
            .ltout(),
            .carryin(bfn_19_29_0_),
            .carryout(\c0.n19470 ),
            .clk(N__66868),
            .ce(),
            .sr(N__50455));
    defparam \c0.add_49_30_THRU_CRY_0_LC_19_29_1 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_0_LC_19_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_0_LC_19_29_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_0_LC_19_29_1  (
            .in0(_gnd_net_),
            .in1(N__46511),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19470 ),
            .carryout(\c0.n19470_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_1_LC_19_29_2 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_1_LC_19_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_1_LC_19_29_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_1_LC_19_29_2  (
            .in0(_gnd_net_),
            .in1(N__46515),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19470_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19470_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_2_LC_19_29_3 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_2_LC_19_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_2_LC_19_29_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_2_LC_19_29_3  (
            .in0(_gnd_net_),
            .in1(N__46512),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19470_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19470_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_3_LC_19_29_4 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_3_LC_19_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_3_LC_19_29_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_3_LC_19_29_4  (
            .in0(_gnd_net_),
            .in1(N__46516),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19470_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19470_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_4_LC_19_29_5 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_4_LC_19_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_4_LC_19_29_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_4_LC_19_29_5  (
            .in0(_gnd_net_),
            .in1(N__46513),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19470_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19470_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_5_LC_19_29_6 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_5_LC_19_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_5_LC_19_29_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_5_LC_19_29_6  (
            .in0(_gnd_net_),
            .in1(N__46517),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19470_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19470_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_6_LC_19_29_7 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_6_LC_19_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_6_LC_19_29_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_6_LC_19_29_7  (
            .in0(_gnd_net_),
            .in1(N__46514),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19470_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19470_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i29_LC_19_30_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i29_LC_19_30_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i29_LC_19_30_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i29_LC_19_30_0  (
            .in0(N__51131),
            .in1(N__45896),
            .in2(_gnd_net_),
            .in3(N__45880),
            .lcout(\c0.FRAME_MATCHER_i_29 ),
            .ltout(),
            .carryin(bfn_19_30_0_),
            .carryout(\c0.n19471 ),
            .clk(N__66871),
            .ce(),
            .sr(N__45955));
    defparam \c0.add_49_31_THRU_CRY_0_LC_19_30_1 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_0_LC_19_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_0_LC_19_30_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_0_LC_19_30_1  (
            .in0(_gnd_net_),
            .in1(N__46518),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19471 ),
            .carryout(\c0.n19471_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_1_LC_19_30_2 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_1_LC_19_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_1_LC_19_30_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_1_LC_19_30_2  (
            .in0(_gnd_net_),
            .in1(N__46522),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19471_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19471_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_2_LC_19_30_3 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_2_LC_19_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_2_LC_19_30_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_2_LC_19_30_3  (
            .in0(_gnd_net_),
            .in1(N__46519),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19471_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19471_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_3_LC_19_30_4 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_3_LC_19_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_3_LC_19_30_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_3_LC_19_30_4  (
            .in0(_gnd_net_),
            .in1(N__46523),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19471_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19471_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_4_LC_19_30_5 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_4_LC_19_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_4_LC_19_30_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_4_LC_19_30_5  (
            .in0(_gnd_net_),
            .in1(N__46520),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19471_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19471_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_5_LC_19_30_6 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_5_LC_19_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_5_LC_19_30_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_5_LC_19_30_6  (
            .in0(_gnd_net_),
            .in1(N__46524),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19471_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19471_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_6_LC_19_30_7 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_6_LC_19_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_6_LC_19_30_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_6_LC_19_30_7  (
            .in0(_gnd_net_),
            .in1(N__46521),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19471_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19471_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i30_LC_19_31_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i30_LC_19_31_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i30_LC_19_31_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i30_LC_19_31_0  (
            .in0(N__51161),
            .in1(N__45936),
            .in2(_gnd_net_),
            .in3(N__45922),
            .lcout(\c0.FRAME_MATCHER_i_30 ),
            .ltout(),
            .carryin(bfn_19_31_0_),
            .carryout(\c0.n19472 ),
            .clk(N__66875),
            .ce(),
            .sr(N__45919));
    defparam \c0.add_49_32_THRU_CRY_0_LC_19_31_1 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_0_LC_19_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_0_LC_19_31_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_0_LC_19_31_1  (
            .in0(_gnd_net_),
            .in1(N__46525),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19472 ),
            .carryout(\c0.n19472_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_1_LC_19_31_2 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_1_LC_19_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_1_LC_19_31_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_1_LC_19_31_2  (
            .in0(_gnd_net_),
            .in1(N__46529),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19472_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19472_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_2_LC_19_31_3 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_2_LC_19_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_2_LC_19_31_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_2_LC_19_31_3  (
            .in0(_gnd_net_),
            .in1(N__46526),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19472_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19472_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_3_LC_19_31_4 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_3_LC_19_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_3_LC_19_31_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_3_LC_19_31_4  (
            .in0(_gnd_net_),
            .in1(N__46530),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19472_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19472_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_4_LC_19_31_5 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_4_LC_19_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_4_LC_19_31_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_4_LC_19_31_5  (
            .in0(_gnd_net_),
            .in1(N__46527),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19472_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19472_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_5_LC_19_31_6 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_5_LC_19_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_5_LC_19_31_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_5_LC_19_31_6  (
            .in0(_gnd_net_),
            .in1(N__46531),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19472_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19472_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_6_LC_19_31_7 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_6_LC_19_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_6_LC_19_31_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_6_LC_19_31_7  (
            .in0(_gnd_net_),
            .in1(N__46528),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19472_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19472_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i31_LC_19_32_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i31_LC_19_32_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i31_LC_19_32_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i31_LC_19_32_0  (
            .in0(N__51162),
            .in1(N__46109),
            .in2(_gnd_net_),
            .in3(N__46180),
            .lcout(\c0.FRAME_MATCHER_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66876),
            .ce(),
            .sr(N__46075));
    defparam \c0.select_365_Select_1_i3_2_lut_4_lut_LC_20_3_4 .C_ON=1'b0;
    defparam \c0.select_365_Select_1_i3_2_lut_4_lut_LC_20_3_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_1_i3_2_lut_4_lut_LC_20_3_4 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_1_i3_2_lut_4_lut_LC_20_3_4  (
            .in0(N__51472),
            .in1(N__51189),
            .in2(N__56544),
            .in3(N__50663),
            .lcout(\c0.n3_adj_4475 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_3_i3_2_lut_4_lut_LC_20_4_2 .C_ON=1'b0;
    defparam \c0.select_365_Select_3_i3_2_lut_4_lut_LC_20_4_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_3_i3_2_lut_4_lut_LC_20_4_2 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_3_i3_2_lut_4_lut_LC_20_4_2  (
            .in0(N__51474),
            .in1(N__51159),
            .in2(N__46014),
            .in3(N__50662),
            .lcout(\c0.n3_adj_4472 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_2_i3_2_lut_4_lut_LC_20_4_6 .C_ON=1'b0;
    defparam \c0.select_365_Select_2_i3_2_lut_4_lut_LC_20_4_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_2_i3_2_lut_4_lut_LC_20_4_6 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_2_i3_2_lut_4_lut_LC_20_4_6  (
            .in0(N__51473),
            .in1(N__51158),
            .in2(N__56403),
            .in3(N__50661),
            .lcout(\c0.n3_adj_4474 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_96_i9_2_lut_3_lut_LC_20_5_4 .C_ON=1'b0;
    defparam \c0.equal_96_i9_2_lut_3_lut_LC_20_5_4 .SEQ_MODE=4'b0000;
    defparam \c0.equal_96_i9_2_lut_3_lut_LC_20_5_4 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \c0.equal_96_i9_2_lut_3_lut_LC_20_5_4  (
            .in0(N__56568),
            .in1(N__56394),
            .in2(_gnd_net_),
            .in3(N__56708),
            .lcout(\c0.n9_adj_4302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_86_i9_2_lut_3_lut_LC_20_6_6 .C_ON=1'b0;
    defparam \c0.equal_86_i9_2_lut_3_lut_LC_20_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.equal_86_i9_2_lut_3_lut_LC_20_6_6 .LUT_INIT=16'b1111111101011111;
    LogicCell40 \c0.equal_86_i9_2_lut_3_lut_LC_20_6_6  (
            .in0(N__56569),
            .in1(_gnd_net_),
            .in2(N__56743),
            .in3(N__56419),
            .lcout(\c0.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_92_i11_2_lut_LC_20_7_6 .C_ON=1'b0;
    defparam \c0.equal_92_i11_2_lut_LC_20_7_6 .SEQ_MODE=4'b0000;
    defparam \c0.equal_92_i11_2_lut_LC_20_7_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.equal_92_i11_2_lut_LC_20_7_6  (
            .in0(_gnd_net_),
            .in1(N__47384),
            .in2(_gnd_net_),
            .in3(N__47347),
            .lcout(\c0.n11_adj_4326 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_LC_20_8_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_LC_20_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_LC_20_8_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_LC_20_8_0  (
            .in0(N__52105),
            .in1(N__52179),
            .in2(N__60154),
            .in3(N__52143),
            .lcout(\c0.n13697 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1622_LC_20_8_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1622_LC_20_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1622_LC_20_8_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i2_2_lut_adj_1622_LC_20_8_1  (
            .in0(N__52144),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48451),
            .lcout(\c0.n10_adj_4399 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1312_LC_20_8_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1312_LC_20_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1312_LC_20_8_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1312_LC_20_8_2  (
            .in0(_gnd_net_),
            .in1(N__48401),
            .in2(_gnd_net_),
            .in3(N__47253),
            .lcout(\c0.n6_adj_4258 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i60_LC_20_8_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i60_LC_20_8_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i60_LC_20_8_3 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i60_LC_20_8_3  (
            .in0(N__60889),
            .in1(N__68568),
            .in2(N__52275),
            .in3(N__64879),
            .lcout(\c0.data_in_frame_7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66657),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1258_LC_20_8_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1258_LC_20_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1258_LC_20_8_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1258_LC_20_8_4  (
            .in0(_gnd_net_),
            .in1(N__54193),
            .in2(_gnd_net_),
            .in3(N__60191),
            .lcout(\c0.n6_adj_4241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i71_LC_20_8_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i71_LC_20_8_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i71_LC_20_8_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i71_LC_20_8_6  (
            .in0(N__62509),
            .in1(N__52106),
            .in2(N__66028),
            .in3(N__65648),
            .lcout(\c0.data_in_frame_8_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66657),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i70_LC_20_8_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i70_LC_20_8_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i70_LC_20_8_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i70_LC_20_8_7  (
            .in0(N__67186),
            .in1(N__66008),
            .in2(N__48410),
            .in3(N__62510),
            .lcout(\c0.data_in_frame_8_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66657),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i88_LC_20_9_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i88_LC_20_9_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i88_LC_20_9_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i88_LC_20_9_0  (
            .in0(N__62374),
            .in1(N__69064),
            .in2(N__49753),
            .in3(N__68954),
            .lcout(\c0.data_in_frame_10_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66662),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i87_LC_20_9_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i87_LC_20_9_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i87_LC_20_9_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i87_LC_20_9_1  (
            .in0(N__69063),
            .in1(N__65576),
            .in2(N__60094),
            .in3(N__62376),
            .lcout(\c0.data_in_frame_10_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66662),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1316_LC_20_9_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1316_LC_20_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1316_LC_20_9_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1316_LC_20_9_2  (
            .in0(_gnd_net_),
            .in1(N__60081),
            .in2(_gnd_net_),
            .in3(N__49736),
            .lcout(\c0.n21925 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1666_LC_20_9_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1666_LC_20_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1666_LC_20_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1666_LC_20_9_3  (
            .in0(N__47548),
            .in1(N__51753),
            .in2(N__47524),
            .in3(N__51700),
            .lcout(\c0.n6_adj_4395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i22_LC_20_9_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i22_LC_20_9_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i22_LC_20_9_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i22_LC_20_9_4  (
            .in0(N__67219),
            .in1(N__60888),
            .in2(N__48204),
            .in3(N__69065),
            .lcout(\c0.data_in_frame_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66662),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i82_LC_20_9_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i82_LC_20_9_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i82_LC_20_9_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i82_LC_20_9_5  (
            .in0(N__69062),
            .in1(N__62375),
            .in2(N__51547),
            .in3(N__63862),
            .lcout(\c0.data_in_frame_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66662),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1311_LC_20_9_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1311_LC_20_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1311_LC_20_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1311_LC_20_9_6  (
            .in0(N__52098),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57712),
            .lcout(),
            .ltout(\c0.n21861_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1313_LC_20_9_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1313_LC_20_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1313_LC_20_9_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1313_LC_20_9_7  (
            .in0(N__47455),
            .in1(N__52206),
            .in2(N__47422),
            .in3(N__47419),
            .lcout(\c0.n21940 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_LC_20_10_0 .C_ON=1'b0;
    defparam \c0.i3_3_lut_LC_20_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_LC_20_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_3_lut_LC_20_10_0  (
            .in0(N__50439),
            .in1(N__51622),
            .in2(_gnd_net_),
            .in3(N__51567),
            .lcout(),
            .ltout(\c0.n8_adj_4254_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1290_LC_20_10_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1290_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1290_LC_20_10_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1290_LC_20_10_1  (
            .in0(N__52274),
            .in1(N__47827),
            .in2(N__47809),
            .in3(N__47806),
            .lcout(\c0.n13865 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i46_LC_20_10_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i46_LC_20_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i46_LC_20_10_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i46_LC_20_10_2  (
            .in0(N__60881),
            .in1(N__62148),
            .in2(N__47787),
            .in3(N__67217),
            .lcout(\c0.data_in_frame_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66668),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1614_LC_20_10_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1614_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1614_LC_20_10_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1614_LC_20_10_3  (
            .in0(N__47766),
            .in1(N__47737),
            .in2(N__47688),
            .in3(N__47707),
            .lcout(\c0.n12484 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i10_LC_20_10_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i10_LC_20_10_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i10_LC_20_10_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i10_LC_20_10_5  (
            .in0(N__69806),
            .in1(N__60882),
            .in2(N__47689),
            .in3(N__63849),
            .lcout(data_in_frame_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66668),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i72_LC_20_10_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i72_LC_20_10_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i72_LC_20_10_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i72_LC_20_10_6  (
            .in0(N__66020),
            .in1(N__62542),
            .in2(N__57731),
            .in3(N__68988),
            .lcout(\c0.data_in_frame_8_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66668),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i6_LC_20_10_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i6_LC_20_10_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i6_LC_20_10_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i6_LC_20_10_7  (
            .in0(N__67216),
            .in1(N__60883),
            .in2(N__51773),
            .in3(N__66021),
            .lcout(\c0.data_in_frame_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66668),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1662_LC_20_11_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1662_LC_20_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1662_LC_20_11_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1662_LC_20_11_0  (
            .in0(N__50341),
            .in1(N__48197),
            .in2(N__48170),
            .in3(N__47640),
            .lcout(),
            .ltout(\c0.n13848_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1630_LC_20_11_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1630_LC_20_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1630_LC_20_11_1 .LUT_INIT=16'b1111111110010110;
    LogicCell40 \c0.i3_4_lut_adj_1630_LC_20_11_1  (
            .in0(N__47968),
            .in1(N__47578),
            .in2(N__47566),
            .in3(N__51970),
            .lcout(\c0.n13_adj_4405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1310_LC_20_11_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1310_LC_20_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1310_LC_20_11_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1310_LC_20_11_2  (
            .in0(N__48233),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47949),
            .lcout(\c0.n13652 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1667_LC_20_11_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1667_LC_20_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1667_LC_20_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1667_LC_20_11_3  (
            .in0(N__48196),
            .in1(N__48158),
            .in2(_gnd_net_),
            .in3(N__50340),
            .lcout(\c0.n13398 ),
            .ltout(\c0.n13398_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1717_LC_20_11_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1717_LC_20_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1717_LC_20_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1717_LC_20_11_4  (
            .in0(N__48048),
            .in1(N__48001),
            .in2(N__47971),
            .in3(N__47967),
            .lcout(\c0.n21794 ),
            .ltout(\c0.n21794_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1824_LC_20_11_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1824_LC_20_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1824_LC_20_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1824_LC_20_11_5  (
            .in0(_gnd_net_),
            .in1(N__47938),
            .in2(N__47911),
            .in3(N__48232),
            .lcout(\c0.n22239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_LC_20_11_6 .C_ON=1'b0;
    defparam \c0.i21_4_lut_LC_20_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_LC_20_11_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i21_4_lut_LC_20_11_6  (
            .in0(N__51508),
            .in1(N__48364),
            .in2(N__52291),
            .in3(N__48340),
            .lcout(\c0.n44_adj_4262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i64_LC_20_11_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i64_LC_20_11_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i64_LC_20_11_7 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.data_in_frame_0__i64_LC_20_11_7  (
            .in0(N__68989),
            .in1(N__68569),
            .in2(N__51919),
            .in3(N__60897),
            .lcout(\c0.data_in_frame_7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66679),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1905_LC_20_12_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1905_LC_20_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1905_LC_20_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1905_LC_20_12_0  (
            .in0(N__47902),
            .in1(N__51974),
            .in2(_gnd_net_),
            .in3(N__48351),
            .lcout(),
            .ltout(\c0.n6_adj_4257_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1308_LC_20_12_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1308_LC_20_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1308_LC_20_12_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1308_LC_20_12_1  (
            .in0(N__51914),
            .in1(N__48279),
            .in2(N__47848),
            .in3(N__47845),
            .lcout(\c0.n13771 ),
            .ltout(\c0.n13771_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1314_LC_20_12_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1314_LC_20_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1314_LC_20_12_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1314_LC_20_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48355),
            .in3(N__54999),
            .lcout(\c0.n4 ),
            .ltout(\c0.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_LC_20_12_3 .C_ON=1'b0;
    defparam \c0.i14_4_lut_LC_20_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_LC_20_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_LC_20_12_3  (
            .in0(N__48352),
            .in1(N__48383),
            .in2(N__48343),
            .in3(N__60054),
            .lcout(\c0.n37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1220_LC_20_12_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1220_LC_20_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1220_LC_20_12_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i2_2_lut_adj_1220_LC_20_12_4  (
            .in0(N__52443),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60435),
            .lcout(\c0.n21967 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1300_LC_20_12_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1300_LC_20_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1300_LC_20_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1300_LC_20_12_5  (
            .in0(N__48334),
            .in1(N__48384),
            .in2(N__48322),
            .in3(N__48292),
            .lcout(\c0.n13425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1402_LC_20_12_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1402_LC_20_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1402_LC_20_12_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1402_LC_20_12_6  (
            .in0(N__61468),
            .in1(N__54175),
            .in2(N__54478),
            .in3(N__48286),
            .lcout(\c0.n21170 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i84_LC_20_12_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i84_LC_20_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i84_LC_20_12_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i84_LC_20_12_7  (
            .in0(N__64836),
            .in1(N__62543),
            .in2(N__69191),
            .in3(N__48280),
            .lcout(\c0.data_in_frame_10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66691),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1252_LC_20_13_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1252_LC_20_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1252_LC_20_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1252_LC_20_13_0  (
            .in0(N__48414),
            .in1(N__60367),
            .in2(N__48271),
            .in3(N__51856),
            .lcout(\c0.n21979 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1302_LC_20_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1302_LC_20_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1302_LC_20_13_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1302_LC_20_13_1  (
            .in0(_gnd_net_),
            .in1(N__48448),
            .in2(_gnd_net_),
            .in3(N__52171),
            .lcout(\c0.n21964 ),
            .ltout(\c0.n21964_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1320_LC_20_13_2 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1320_LC_20_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1320_LC_20_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_1320_LC_20_13_2  (
            .in0(N__60973),
            .in1(N__48262),
            .in2(N__48244),
            .in3(N__48240),
            .lcout(\c0.n40_adj_4261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1259_LC_20_13_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1259_LC_20_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1259_LC_20_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1259_LC_20_13_3  (
            .in0(N__49755),
            .in1(N__49779),
            .in2(N__48466),
            .in3(N__63969),
            .lcout(\c0.n21864 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1328_LC_20_13_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1328_LC_20_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1328_LC_20_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1328_LC_20_13_4  (
            .in0(N__48449),
            .in1(N__60520),
            .in2(N__48415),
            .in3(N__49754),
            .lcout(\c0.n22415 ),
            .ltout(\c0.n22415_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1833_LC_20_13_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1833_LC_20_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1833_LC_20_13_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1833_LC_20_13_5  (
            .in0(N__52107),
            .in1(_gnd_net_),
            .in2(N__48388),
            .in3(N__57730),
            .lcout(\c0.n6_adj_4256 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i73_LC_20_13_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i73_LC_20_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i73_LC_20_13_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i73_LC_20_13_6  (
            .in0(N__69750),
            .in1(N__62554),
            .in2(N__52207),
            .in3(N__69557),
            .lcout(\c0.data_in_frame_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66705),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1275_LC_20_14_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1275_LC_20_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1275_LC_20_14_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1275_LC_20_14_2  (
            .in0(_gnd_net_),
            .in1(N__61807),
            .in2(_gnd_net_),
            .in3(N__55326),
            .lcout(\c0.n13681 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i61_LC_20_14_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i61_LC_20_14_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i61_LC_20_14_3 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \c0.data_in_frame_0__i61_LC_20_14_3  (
            .in0(N__63205),
            .in1(N__50438),
            .in2(N__60887),
            .in3(N__68674),
            .lcout(\c0.data_in_frame_7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66719),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1841_LC_20_14_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1841_LC_20_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1841_LC_20_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1841_LC_20_14_4  (
            .in0(N__61813),
            .in1(N__55327),
            .in2(_gnd_net_),
            .in3(N__57490),
            .lcout(\c0.n22355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i135_LC_20_14_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i135_LC_20_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i135_LC_20_14_5 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0__i135_LC_20_14_5  (
            .in0(N__52375),
            .in1(N__68095),
            .in2(N__66019),
            .in3(N__65661),
            .lcout(\c0.data_in_frame_16_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66719),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i86_LC_20_14_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i86_LC_20_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i86_LC_20_14_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i86_LC_20_14_6  (
            .in0(N__69125),
            .in1(N__62396),
            .in2(N__48385),
            .in3(N__67163),
            .lcout(\c0.data_in_frame_10_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66719),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_3_lut_4_lut_LC_20_14_7 .C_ON=1'b0;
    defparam \c0.i12_3_lut_4_lut_LC_20_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i12_3_lut_4_lut_LC_20_14_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_3_lut_4_lut_LC_20_14_7  (
            .in0(N__52534),
            .in1(N__54709),
            .in2(N__54893),
            .in3(N__54561),
            .lcout(\c0.n35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i142_LC_20_15_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i142_LC_20_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i142_LC_20_15_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i142_LC_20_15_0  (
            .in0(N__69695),
            .in1(N__68092),
            .in2(N__55338),
            .in3(N__67162),
            .lcout(\c0.data_in_frame_17_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66733),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i77_LC_20_15_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i77_LC_20_15_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i77_LC_20_15_1 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i77_LC_20_15_1  (
            .in0(N__63143),
            .in1(N__69697),
            .in2(N__52480),
            .in3(N__62430),
            .lcout(\c0.data_in_frame_9_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66733),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1263_LC_20_15_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1263_LC_20_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1263_LC_20_15_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1263_LC_20_15_2  (
            .in0(_gnd_net_),
            .in1(N__52476),
            .in2(_gnd_net_),
            .in3(N__57643),
            .lcout(\c0.n6_adj_4243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i143_LC_20_15_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i143_LC_20_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i143_LC_20_15_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i143_LC_20_15_3  (
            .in0(N__68091),
            .in1(N__69696),
            .in2(N__61823),
            .in3(N__65563),
            .lcout(\c0.data_in_frame_17_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66733),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i53_LC_20_15_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i53_LC_20_15_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i53_LC_20_15_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i53_LC_20_15_4  (
            .in0(N__49708),
            .in1(N__63144),
            .in2(_gnd_net_),
            .in3(N__49608),
            .lcout(data_in_frame_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66733),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1584_LC_20_15_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1584_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1584_LC_20_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1584_LC_20_15_5  (
            .in0(N__49654),
            .in1(N__49641),
            .in2(N__49609),
            .in3(N__49589),
            .lcout(\c0.n13605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i35_LC_20_15_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i35_LC_20_15_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i35_LC_20_15_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i35_LC_20_15_6  (
            .in0(N__68373),
            .in1(N__64518),
            .in2(N__49596),
            .in3(N__60727),
            .lcout(\c0.data_in_frame_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66733),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__6__5471_LC_20_15_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__6__5471_LC_20_15_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__6__5471_LC_20_15_7 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_6__6__5471_LC_20_15_7  (
            .in0(N__49356),
            .in1(N__49012),
            .in2(N__48571),
            .in3(N__48480),
            .lcout(data_out_frame_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66733),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1329_LC_20_16_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1329_LC_20_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1329_LC_20_16_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1329_LC_20_16_0  (
            .in0(_gnd_net_),
            .in1(N__60399),
            .in2(_gnd_net_),
            .in3(N__60196),
            .lcout(),
            .ltout(\c0.n22440_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1235_LC_20_16_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1235_LC_20_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1235_LC_20_16_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1235_LC_20_16_1  (
            .in0(N__52629),
            .in1(N__49783),
            .in2(N__49762),
            .in3(N__52608),
            .lcout(),
            .ltout(\c0.n10_adj_4229_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1860_LC_20_16_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1860_LC_20_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1860_LC_20_16_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1860_LC_20_16_2  (
            .in0(N__60101),
            .in1(N__49759),
            .in2(N__49720),
            .in3(N__55015),
            .lcout(\c0.n5943 ),
            .ltout(\c0.n5943_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1754_LC_20_16_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1754_LC_20_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1754_LC_20_16_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1754_LC_20_16_3  (
            .in0(N__55328),
            .in1(N__55217),
            .in2(N__49717),
            .in3(N__55303),
            .lcout(\c0.n22081 ),
            .ltout(\c0.n22081_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1273_LC_20_16_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1273_LC_20_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1273_LC_20_16_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_3_lut_adj_1273_LC_20_16_4  (
            .in0(N__61615),
            .in1(_gnd_net_),
            .in2(N__49714),
            .in3(N__55395),
            .lcout(\c0.n13457 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1894_LC_20_16_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1894_LC_20_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1894_LC_20_16_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1894_LC_20_16_5  (
            .in0(N__55396),
            .in1(N__61616),
            .in2(N__61216),
            .in3(N__53218),
            .lcout(\c0.n13443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1221_LC_20_16_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1221_LC_20_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1221_LC_20_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1221_LC_20_16_6  (
            .in0(N__52378),
            .in1(N__55126),
            .in2(_gnd_net_),
            .in3(N__52348),
            .lcout(\c0.n21187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1580_LC_20_17_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1580_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1580_LC_20_17_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1580_LC_20_17_0  (
            .in0(N__55624),
            .in1(N__63356),
            .in2(N__64030),
            .in3(N__61603),
            .lcout(\c0.n22349 ),
            .ltout(\c0.n22349_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1616_LC_20_17_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1616_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1616_LC_20_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1616_LC_20_17_1  (
            .in0(N__57446),
            .in1(N__61420),
            .in2(N__49711),
            .in3(N__55431),
            .lcout(\c0.n6_adj_4224 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1857_LC_20_17_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1857_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1857_LC_20_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1857_LC_20_17_2  (
            .in0(N__55430),
            .in1(N__61415),
            .in2(_gnd_net_),
            .in3(N__57445),
            .lcout(),
            .ltout(\c0.n21858_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1247_LC_20_17_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1247_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1247_LC_20_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1247_LC_20_17_3  (
            .in0(N__55385),
            .in1(N__64017),
            .in2(N__49900),
            .in3(N__55623),
            .lcout(\c0.n21989 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i159_LC_20_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i159_LC_20_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i159_LC_20_17_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i159_LC_20_17_4  (
            .in0(N__68007),
            .in1(N__67339),
            .in2(N__61617),
            .in3(N__65568),
            .lcout(\c0.data_in_frame_19_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66761),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i215_LC_20_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i215_LC_20_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i215_LC_20_17_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i215_LC_20_17_5  (
            .in0(N__65567),
            .in1(N__69249),
            .in2(N__59439),
            .in3(N__67677),
            .lcout(\c0.data_in_frame_26_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66761),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i139_LC_20_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i139_LC_20_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i139_LC_20_17_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i139_LC_20_17_6  (
            .in0(N__68006),
            .in1(N__69802),
            .in2(N__68436),
            .in3(N__61416),
            .lcout(\c0.data_in_frame_17_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66761),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i138_LC_20_17_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i138_LC_20_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i138_LC_20_17_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i138_LC_20_17_7  (
            .in0(N__69801),
            .in1(N__68008),
            .in2(N__64035),
            .in3(N__63764),
            .lcout(\c0.data_in_frame_17_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66761),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1567_LC_20_18_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1567_LC_20_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1567_LC_20_18_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_1567_LC_20_18_0  (
            .in0(N__50710),
            .in1(N__49890),
            .in2(N__50010),
            .in3(N__49857),
            .lcout(\c0.n16_adj_4375 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_13_i3_2_lut_4_lut_LC_20_18_1 .C_ON=1'b0;
    defparam \c0.select_365_Select_13_i3_2_lut_4_lut_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_13_i3_2_lut_4_lut_LC_20_18_1 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_13_i3_2_lut_4_lut_LC_20_18_1  (
            .in0(N__51433),
            .in1(N__51041),
            .in2(N__49861),
            .in3(N__50609),
            .lcout(\c0.n3_adj_4454 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i172_LC_20_18_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i172_LC_20_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i172_LC_20_18_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i172_LC_20_18_2  (
            .in0(N__62184),
            .in1(N__68067),
            .in2(N__49939),
            .in3(N__64871),
            .lcout(\c0.data_in_frame_21_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66773),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1211_LC_20_18_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1211_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1211_LC_20_18_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1211_LC_20_18_3  (
            .in0(N__63486),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65248),
            .lcout(\c0.n22028 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_15_i3_2_lut_4_lut_LC_20_18_4 .C_ON=1'b0;
    defparam \c0.select_365_Select_15_i3_2_lut_4_lut_LC_20_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_15_i3_2_lut_4_lut_LC_20_18_4 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \c0.select_365_Select_15_i3_2_lut_4_lut_LC_20_18_4  (
            .in0(N__50610),
            .in1(N__49821),
            .in2(N__51111),
            .in3(N__51435),
            .lcout(\c0.n3_adj_4452 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i185_LC_20_18_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i185_LC_20_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i185_LC_20_18_5 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i185_LC_20_18_5  (
            .in0(N__68065),
            .in1(N__68670),
            .in2(N__63268),
            .in3(N__69503),
            .lcout(\c0.data_in_frame_23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66773),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i171_LC_20_18_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i171_LC_20_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i171_LC_20_18_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i171_LC_20_18_6  (
            .in0(N__62183),
            .in1(N__68066),
            .in2(N__53818),
            .in3(N__68369),
            .lcout(\c0.data_in_frame_21_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66773),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_20_i3_2_lut_4_lut_LC_20_18_7 .C_ON=1'b0;
    defparam \c0.select_365_Select_20_i3_2_lut_4_lut_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_20_i3_2_lut_4_lut_LC_20_18_7 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_20_i3_2_lut_4_lut_LC_20_18_7  (
            .in0(N__51434),
            .in1(N__51042),
            .in2(N__50011),
            .in3(N__50611),
            .lcout(\c0.n3_adj_4442 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1369_LC_20_19_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1369_LC_20_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1369_LC_20_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1369_LC_20_19_0  (
            .in0(N__53602),
            .in1(N__65322),
            .in2(N__49969),
            .in3(N__53788),
            .lcout(\c0.n12_adj_4290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1214_LC_20_19_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1214_LC_20_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1214_LC_20_19_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1214_LC_20_19_1  (
            .in0(_gnd_net_),
            .in1(N__53809),
            .in2(_gnd_net_),
            .in3(N__49934),
            .lcout(\c0.n21870 ),
            .ltout(\c0.n21870_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1192_LC_20_19_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1192_LC_20_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1192_LC_20_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1192_LC_20_19_2  (
            .in0(N__50073),
            .in1(N__55486),
            .in2(N__49942),
            .in3(N__55540),
            .lcout(\c0.n13761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1350_LC_20_19_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1350_LC_20_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1350_LC_20_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1350_LC_20_19_3  (
            .in0(N__55919),
            .in1(N__50072),
            .in2(_gnd_net_),
            .in3(N__49920),
            .lcout(\c0.n22396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_LC_20_19_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_LC_20_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_LC_20_19_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i2_2_lut_LC_20_19_4  (
            .in0(N__49935),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49921),
            .lcout(\c0.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i207_LC_20_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i207_LC_20_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i207_LC_20_19_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i207_LC_20_19_5  (
            .in0(N__69730),
            .in1(N__65573),
            .in2(N__58610),
            .in3(N__67707),
            .lcout(\c0.data_in_frame_25_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66787),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i191_LC_20_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i191_LC_20_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i191_LC_20_19_6 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \c0.data_in_frame_0__i191_LC_20_19_6  (
            .in0(N__65572),
            .in1(N__55920),
            .in2(N__68679),
            .in3(N__68069),
            .lcout(\c0.data_in_frame_23_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66787),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i189_LC_20_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i189_LC_20_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i189_LC_20_19_7 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_in_frame_0__i189_LC_20_19_7  (
            .in0(N__68068),
            .in1(N__68669),
            .in2(N__63172),
            .in3(N__50074),
            .lcout(\c0.data_in_frame_23_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66787),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1195_LC_20_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1195_LC_20_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1195_LC_20_20_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1195_LC_20_20_0  (
            .in0(N__53601),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53728),
            .lcout(\c0.n13266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1363_LC_20_20_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1363_LC_20_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1363_LC_20_20_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1363_LC_20_20_1  (
            .in0(N__56059),
            .in1(N__54135),
            .in2(N__53941),
            .in3(N__59023),
            .lcout(),
            .ltout(\c0.n10_adj_4287_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1384_LC_20_20_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1384_LC_20_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1384_LC_20_20_2 .LUT_INIT=16'b1101111011101101;
    LogicCell40 \c0.i4_4_lut_adj_1384_LC_20_20_2  (
            .in0(N__50204),
            .in1(N__50017),
            .in2(N__50062),
            .in3(N__56326),
            .lcout(\c0.n22_adj_4298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i157_LC_20_20_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i157_LC_20_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i157_LC_20_20_4 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i157_LC_20_20_4  (
            .in0(N__63058),
            .in1(N__68070),
            .in2(N__67402),
            .in3(N__55876),
            .lcout(\c0.data_in_frame_19_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66798),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1721_LC_20_20_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1721_LC_20_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1721_LC_20_20_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_1721_LC_20_20_5  (
            .in0(_gnd_net_),
            .in1(N__53600),
            .in2(_gnd_net_),
            .in3(N__54007),
            .lcout(\c0.n10_adj_4483 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1899_LC_20_21_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1899_LC_20_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1899_LC_20_21_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1899_LC_20_21_0  (
            .in0(N__53654),
            .in1(N__53979),
            .in2(N__66913),
            .in3(N__53767),
            .lcout(\c0.n21233 ),
            .ltout(\c0.n21233_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1364_LC_20_21_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1364_LC_20_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1364_LC_20_21_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_1364_LC_20_21_1  (
            .in0(N__50047),
            .in1(N__50038),
            .in2(N__50020),
            .in3(N__53986),
            .lcout(\c0.n23506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i239_LC_20_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i239_LC_20_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i239_LC_20_21_3 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i239_LC_20_21_3  (
            .in0(N__65562),
            .in1(N__54112),
            .in2(N__62202),
            .in3(N__67708),
            .lcout(\c0.data_in_frame_29_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66807),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1727_LC_20_21_7 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1727_LC_20_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1727_LC_20_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_1727_LC_20_21_7  (
            .in0(N__50206),
            .in1(N__58770),
            .in2(N__65103),
            .in3(N__59419),
            .lcout(\c0.n45_adj_4486 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i158_LC_20_22_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i158_LC_20_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i158_LC_20_22_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i158_LC_20_22_5  (
            .in0(N__68140),
            .in1(N__67392),
            .in2(N__58835),
            .in3(N__67218),
            .lcout(\c0.data_in_frame_19_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66819),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_365_Select_10_i3_2_lut_4_lut_LC_20_22_6 .C_ON=1'b0;
    defparam \c0.select_365_Select_10_i3_2_lut_4_lut_LC_20_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_10_i3_2_lut_4_lut_LC_20_22_6 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_10_i3_2_lut_4_lut_LC_20_22_6  (
            .in0(N__51436),
            .in1(N__51069),
            .in2(N__50167),
            .in3(N__50620),
            .lcout(\c0.n3_adj_4460 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i155_LC_20_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i155_LC_20_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i155_LC_20_22_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i155_LC_20_22_7  (
            .in0(N__68139),
            .in1(N__67391),
            .in2(N__56006),
            .in3(N__68412),
            .lcout(\c0.data_in_frame_19_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66819),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i1_LC_20_23_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i1_LC_20_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i1_LC_20_23_0 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.rx.r_Rx_Byte_i1_LC_20_23_0  (
            .in0(N__63643),
            .in1(N__50106),
            .in2(N__59716),
            .in3(N__56207),
            .lcout(rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66831),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i221_LC_20_23_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i221_LC_20_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i221_LC_20_23_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i221_LC_20_23_2  (
            .in0(N__67348),
            .in1(N__63092),
            .in2(N__55839),
            .in3(N__67752),
            .lcout(\c0.data_in_frame_27_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66831),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_LC_20_23_3 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_LC_20_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_LC_20_23_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.rx.i2_3_lut_LC_20_23_3  (
            .in0(N__50229),
            .in1(N__50259),
            .in2(_gnd_net_),
            .in3(N__50244),
            .lcout(\c0.rx.n18655 ),
            .ltout(\c0.rx.n18655_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3_4_lut_LC_20_23_4 .C_ON=1'b0;
    defparam \c0.rx.i3_4_lut_LC_20_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3_4_lut_LC_20_23_4 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \c0.rx.i3_4_lut_LC_20_23_4  (
            .in0(N__54261),
            .in1(N__54284),
            .in2(N__50080),
            .in3(N__54321),
            .lcout(\c0.rx.n21704 ),
            .ltout(\c0.rx.n21704_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i18882_2_lut_LC_20_23_5 .C_ON=1'b0;
    defparam \c0.rx.i18882_2_lut_LC_20_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i18882_2_lut_LC_20_23_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \c0.rx.i18882_2_lut_LC_20_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50077),
            .in3(N__59711),
            .lcout(),
            .ltout(\c0.rx.n22573_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i25_4_lut_LC_20_23_6 .C_ON=1'b0;
    defparam \c0.rx.i25_4_lut_LC_20_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i25_4_lut_LC_20_23_6 .LUT_INIT=16'b0100011111001100;
    LogicCell40 \c0.rx.i25_4_lut_LC_20_23_6  (
            .in0(N__57059),
            .in1(N__56898),
            .in2(N__50269),
            .in3(N__56835),
            .lcout(),
            .ltout(\c0.rx.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i1_LC_20_23_7 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i1_LC_20_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i1_LC_20_23_7 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \c0.rx.r_SM_Main_i1_LC_20_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50266),
            .in3(N__57003),
            .lcout(r_SM_Main_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66831),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i0_LC_20_24_0 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i0_LC_20_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i0_LC_20_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i0_LC_20_24_0  (
            .in0(_gnd_net_),
            .in1(N__54285),
            .in2(_gnd_net_),
            .in3(N__50263),
            .lcout(\c0.rx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(bfn_20_24_0_),
            .carryout(\c0.rx.n19533 ),
            .clk(N__66843),
            .ce(N__51499),
            .sr(N__51484));
    defparam \c0.rx.r_Clock_Count__i1_LC_20_24_1 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i1_LC_20_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i1_LC_20_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i1_LC_20_24_1  (
            .in0(_gnd_net_),
            .in1(N__50260),
            .in2(_gnd_net_),
            .in3(N__50248),
            .lcout(\c0.rx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\c0.rx.n19533 ),
            .carryout(\c0.rx.n19534 ),
            .clk(N__66843),
            .ce(N__51499),
            .sr(N__51484));
    defparam \c0.rx.r_Clock_Count__i2_LC_20_24_2 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i2_LC_20_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i2_LC_20_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i2_LC_20_24_2  (
            .in0(_gnd_net_),
            .in1(N__50245),
            .in2(_gnd_net_),
            .in3(N__50233),
            .lcout(\c0.rx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\c0.rx.n19534 ),
            .carryout(\c0.rx.n19535 ),
            .clk(N__66843),
            .ce(N__51499),
            .sr(N__51484));
    defparam \c0.rx.r_Clock_Count__i3_LC_20_24_3 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i3_LC_20_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i3_LC_20_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i3_LC_20_24_3  (
            .in0(_gnd_net_),
            .in1(N__50230),
            .in2(_gnd_net_),
            .in3(N__50218),
            .lcout(\c0.rx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\c0.rx.n19535 ),
            .carryout(\c0.rx.n19536 ),
            .clk(N__66843),
            .ce(N__51499),
            .sr(N__51484));
    defparam \c0.rx.r_Clock_Count__i4_LC_20_24_4 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i4_LC_20_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i4_LC_20_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i4_LC_20_24_4  (
            .in0(_gnd_net_),
            .in1(N__54322),
            .in2(_gnd_net_),
            .in3(N__50215),
            .lcout(\c0.rx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\c0.rx.n19536 ),
            .carryout(\c0.rx.n19537 ),
            .clk(N__66843),
            .ce(N__51499),
            .sr(N__51484));
    defparam \c0.rx.r_Clock_Count__i5_LC_20_24_5 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i5_LC_20_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i5_LC_20_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i5_LC_20_24_5  (
            .in0(_gnd_net_),
            .in1(N__54043),
            .in2(_gnd_net_),
            .in3(N__50212),
            .lcout(\c0.rx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\c0.rx.n19537 ),
            .carryout(\c0.rx.n19538 ),
            .clk(N__66843),
            .ce(N__51499),
            .sr(N__51484));
    defparam \c0.rx.r_Clock_Count__i6_LC_20_24_6 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i6_LC_20_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i6_LC_20_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i6_LC_20_24_6  (
            .in0(_gnd_net_),
            .in1(N__54031),
            .in2(_gnd_net_),
            .in3(N__50209),
            .lcout(\c0.rx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\c0.rx.n19538 ),
            .carryout(\c0.rx.n19539 ),
            .clk(N__66843),
            .ce(N__51499),
            .sr(N__51484));
    defparam \c0.rx.r_Clock_Count__i7_LC_20_24_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i7_LC_20_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i7_LC_20_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i7_LC_20_24_7  (
            .in0(_gnd_net_),
            .in1(N__54055),
            .in2(_gnd_net_),
            .in3(N__51502),
            .lcout(\c0.rx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66843),
            .ce(N__51499),
            .sr(N__51484));
    defparam \c0.select_365_Select_28_i3_2_lut_4_lut_LC_20_27_4 .C_ON=1'b0;
    defparam \c0.select_365_Select_28_i3_2_lut_4_lut_LC_20_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_365_Select_28_i3_2_lut_4_lut_LC_20_27_4 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.select_365_Select_28_i3_2_lut_4_lut_LC_20_27_4  (
            .in0(N__51466),
            .in1(N__51098),
            .in2(N__50709),
            .in3(N__50621),
            .lcout(\c0.n3_adj_4430 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1617_LC_21_8_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1617_LC_21_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1617_LC_21_8_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1617_LC_21_8_1  (
            .in0(N__51623),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51571),
            .lcout(\c0.n13555 ),
            .ltout(\c0.n13555_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1285_LC_21_8_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1285_LC_21_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1285_LC_21_8_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1285_LC_21_8_2  (
            .in0(N__52510),
            .in1(N__50443),
            .in2(N__50416),
            .in3(N__52229),
            .lcout(\c0.n22043 ),
            .ltout(\c0.n22043_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1837_LC_21_8_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1837_LC_21_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1837_LC_21_8_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1837_LC_21_8_3  (
            .in0(N__50403),
            .in1(N__51596),
            .in2(N__50392),
            .in3(N__54683),
            .lcout(\c0.n21097 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_87_i9_2_lut_3_lut_LC_21_8_5 .C_ON=1'b0;
    defparam \c0.equal_87_i9_2_lut_3_lut_LC_21_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.equal_87_i9_2_lut_3_lut_LC_21_8_5 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.equal_87_i9_2_lut_3_lut_LC_21_8_5  (
            .in0(N__56729),
            .in1(N__56582),
            .in2(_gnd_net_),
            .in3(N__56455),
            .lcout(\c0.n9_adj_4341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i33_LC_21_9_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i33_LC_21_9_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i33_LC_21_9_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i33_LC_21_9_0  (
            .in0(N__64549),
            .in1(N__60892),
            .in2(N__54436),
            .in3(N__69568),
            .lcout(\c0.data_in_frame_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66669),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i62_LC_21_9_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i62_LC_21_9_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i62_LC_21_9_1 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \c0.data_in_frame_0__i62_LC_21_9_1  (
            .in0(N__60891),
            .in1(N__67142),
            .in2(N__51598),
            .in3(N__68600),
            .lcout(\c0.data_in_frame_7_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66669),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_LC_21_9_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_LC_21_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_LC_21_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_LC_21_9_3  (
            .in0(N__50389),
            .in1(N__50349),
            .in2(N__50281),
            .in3(N__51754),
            .lcout(\c0.n13488 ),
            .ltout(\c0.n13488_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1321_LC_21_9_4 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1321_LC_21_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1321_LC_21_9_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_1321_LC_21_9_4  (
            .in0(N__51820),
            .in1(N__51592),
            .in2(N__51805),
            .in3(N__51802),
            .lcout(\c0.n39_adj_4263 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i44_LC_21_9_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i44_LC_21_9_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i44_LC_21_9_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i44_LC_21_9_5  (
            .in0(N__60890),
            .in1(N__62088),
            .in2(N__51630),
            .in3(N__64888),
            .lcout(\c0.data_in_frame_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66669),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20132_2_lut_LC_21_9_7 .C_ON=1'b0;
    defparam \c0.i20132_2_lut_LC_21_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i20132_2_lut_LC_21_9_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i20132_2_lut_LC_21_9_7  (
            .in0(_gnd_net_),
            .in1(N__51755),
            .in2(_gnd_net_),
            .in3(N__51710),
            .lcout(\c0.n23827 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1821_LC_21_10_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1821_LC_21_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1821_LC_21_10_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1821_LC_21_10_0  (
            .in0(N__51631),
            .in1(N__54682),
            .in2(N__51597),
            .in3(N__51566),
            .lcout(),
            .ltout(\c0.n20368_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1745_LC_21_10_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1745_LC_21_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1745_LC_21_10_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1745_LC_21_10_1  (
            .in0(N__51997),
            .in1(N__52006),
            .in2(N__51550),
            .in3(N__51837),
            .lcout(\c0.n22133 ),
            .ltout(\c0.n22133_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1315_LC_21_10_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1315_LC_21_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1315_LC_21_10_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1315_LC_21_10_2  (
            .in0(N__57369),
            .in1(N__51543),
            .in2(N__51526),
            .in3(N__51892),
            .lcout(\c0.n20927 ),
            .ltout(\c0.n20927_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1319_LC_21_10_3 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1319_LC_21_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1319_LC_21_10_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1319_LC_21_10_3  (
            .in0(N__51523),
            .in1(N__52330),
            .in2(N__51517),
            .in3(N__51514),
            .lcout(\c0.n36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1317_LC_21_10_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1317_LC_21_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1317_LC_21_10_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_1317_LC_21_10_4  (
            .in0(N__54777),
            .in1(_gnd_net_),
            .in2(N__51918),
            .in3(_gnd_net_),
            .lcout(\c0.n22379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1555_LC_21_10_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1555_LC_21_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1555_LC_21_10_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1555_LC_21_10_5  (
            .in0(_gnd_net_),
            .in1(N__52050),
            .in2(_gnd_net_),
            .in3(N__54399),
            .lcout(\c0.n22334 ),
            .ltout(\c0.n22334_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_1408_i15_2_lut_3_lut_LC_21_10_6 .C_ON=1'b0;
    defparam \c0.equal_1408_i15_2_lut_3_lut_LC_21_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.equal_1408_i15_2_lut_3_lut_LC_21_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.equal_1408_i15_2_lut_3_lut_LC_21_10_6  (
            .in0(_gnd_net_),
            .in1(N__51836),
            .in2(N__52000),
            .in3(N__51996),
            .lcout(\c0.n15_adj_4404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1809_LC_21_10_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1809_LC_21_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1809_LC_21_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1809_LC_21_10_7  (
            .in0(N__51943),
            .in1(N__51910),
            .in2(_gnd_net_),
            .in3(N__54776),
            .lcout(\c0.n6_adj_4259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1296_LC_21_11_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1296_LC_21_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1296_LC_21_11_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1296_LC_21_11_0  (
            .in0(N__51855),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54214),
            .lcout(\c0.n22270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1318_LC_21_11_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1318_LC_21_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1318_LC_21_11_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1318_LC_21_11_1  (
            .in0(_gnd_net_),
            .in1(N__59244),
            .in2(_gnd_net_),
            .in3(N__57889),
            .lcout(\c0.n22060 ),
            .ltout(\c0.n22060_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1323_LC_21_11_2 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1323_LC_21_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1323_LC_21_11_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_4_lut_adj_1323_LC_21_11_2  (
            .in0(N__51886),
            .in1(N__51877),
            .in2(N__51868),
            .in3(N__51865),
            .lcout(),
            .ltout(\c0.n11_adj_4266_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1324_LC_21_11_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1324_LC_21_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1324_LC_21_11_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1324_LC_21_11_3  (
            .in0(N__54588),
            .in1(N__57655),
            .in2(N__51859),
            .in3(N__51854),
            .lcout(),
            .ltout(\c0.n22842_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1326_LC_21_11_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1326_LC_21_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1326_LC_21_11_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_1326_LC_21_11_4  (
            .in0(N__60363),
            .in1(N__52309),
            .in2(N__51841),
            .in3(N__52596),
            .lcout(\c0.n15_adj_4269 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i47_LC_21_11_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i47_LC_21_11_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i47_LC_21_11_5 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i47_LC_21_11_5  (
            .in0(N__65689),
            .in1(N__51838),
            .in2(N__62177),
            .in3(N__60807),
            .lcout(\c0.data_in_frame_5_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66692),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1298_LC_21_11_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1298_LC_21_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1298_LC_21_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1298_LC_21_11_6  (
            .in0(_gnd_net_),
            .in1(N__59579),
            .in2(_gnd_net_),
            .in3(N__57581),
            .lcout(\c0.n22245 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_LC_21_12_0 .C_ON=1'b0;
    defparam \c0.i15_4_lut_LC_21_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_LC_21_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_LC_21_12_0  (
            .in0(N__52461),
            .in1(N__52132),
            .in2(N__52303),
            .in3(N__52505),
            .lcout(\c0.n38_adj_4260 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1294_LC_21_12_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1294_LC_21_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1294_LC_21_12_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1294_LC_21_12_1  (
            .in0(N__61062),
            .in1(N__52282),
            .in2(N__57619),
            .in3(N__54601),
            .lcout(\c0.n5810 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1332_LC_21_12_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1332_LC_21_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1332_LC_21_12_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1332_LC_21_12_2  (
            .in0(_gnd_net_),
            .in1(N__52276),
            .in2(_gnd_net_),
            .in3(N__52233),
            .lcout(\c0.n22139 ),
            .ltout(\c0.n22139_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1336_LC_21_12_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1336_LC_21_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1336_LC_21_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1336_LC_21_12_3  (
            .in0(N__54859),
            .in1(N__52462),
            .in2(N__52210),
            .in3(N__61024),
            .lcout(\c0.n20135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1339_LC_21_12_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1339_LC_21_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1339_LC_21_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1339_LC_21_12_5  (
            .in0(N__52133),
            .in1(N__54894),
            .in2(N__52329),
            .in3(N__57732),
            .lcout(\c0.n10_adj_4274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1230_LC_21_12_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1230_LC_21_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1230_LC_21_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1230_LC_21_12_6  (
            .in0(N__52202),
            .in1(N__52178),
            .in2(_gnd_net_),
            .in3(N__52134),
            .lcout(\c0.n21822 ),
            .ltout(\c0.n21822_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1292_LC_21_12_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1292_LC_21_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1292_LC_21_12_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1292_LC_21_12_7  (
            .in0(N__57615),
            .in1(N__52111),
            .in2(N__52072),
            .in3(N__54600),
            .lcout(\c0.n22221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1239_LC_21_13_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1239_LC_21_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1239_LC_21_13_0 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i1_2_lut_adj_1239_LC_21_13_0  (
            .in0(N__52377),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52344),
            .lcout(\c0.n22242 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1397_LC_21_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1397_LC_21_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1397_LC_21_13_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1397_LC_21_13_1  (
            .in0(N__54174),
            .in1(_gnd_net_),
            .in2(N__61501),
            .in3(N__54477),
            .lcout(\c0.n22296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1261_LC_21_13_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1261_LC_21_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1261_LC_21_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1261_LC_21_13_2  (
            .in0(N__52426),
            .in1(N__57346),
            .in2(N__57244),
            .in3(N__61496),
            .lcout(),
            .ltout(\c0.n10_adj_4242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1907_LC_21_13_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1907_LC_21_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1907_LC_21_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1907_LC_21_13_3  (
            .in0(N__52535),
            .in1(N__54710),
            .in2(N__52411),
            .in3(N__52408),
            .lcout(\c0.n13786 ),
            .ltout(\c0.n13786_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_LC_21_13_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_LC_21_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_LC_21_13_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_2_lut_4_lut_LC_21_13_4  (
            .in0(N__52376),
            .in1(N__57285),
            .in2(N__52351),
            .in3(N__52343),
            .lcout(\c0.n7_adj_4235 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i184_LC_21_13_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i184_LC_21_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i184_LC_21_13_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i184_LC_21_13_5  (
            .in0(N__60310),
            .in1(N__68987),
            .in2(_gnd_net_),
            .in3(N__59199),
            .lcout(data_in_frame_22_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66720),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i74_LC_21_13_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i74_LC_21_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i74_LC_21_13_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i74_LC_21_13_6  (
            .in0(N__69839),
            .in1(N__63779),
            .in2(N__54633),
            .in3(N__62501),
            .lcout(\c0.data_in_frame_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66720),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1337_LC_21_13_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1337_LC_21_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1337_LC_21_13_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1337_LC_21_13_7  (
            .in0(_gnd_net_),
            .in1(N__60007),
            .in2(_gnd_net_),
            .in3(N__54626),
            .lcout(\c0.n13974 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i58_LC_21_14_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i58_LC_21_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i58_LC_21_14_0 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i58_LC_21_14_0  (
            .in0(N__68672),
            .in1(N__60806),
            .in2(N__54895),
            .in3(N__63800),
            .lcout(\c0.data_in_frame_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66734),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1873_LC_21_14_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1873_LC_21_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1873_LC_21_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1873_LC_21_14_1  (
            .in0(N__55102),
            .in1(N__55064),
            .in2(_gnd_net_),
            .in3(N__54500),
            .lcout(\c0.n6_adj_4221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i81_LC_21_14_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i81_LC_21_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i81_LC_21_14_2 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i81_LC_21_14_2  (
            .in0(N__69480),
            .in1(N__62498),
            .in2(N__69192),
            .in3(N__54714),
            .lcout(\c0.data_in_frame_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66734),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i121_LC_21_14_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i121_LC_21_14_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i121_LC_21_14_3 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i121_LC_21_14_3  (
            .in0(N__62496),
            .in1(N__68673),
            .in2(N__54507),
            .in3(N__69481),
            .lcout(\c0.data_in_frame_15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66734),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i83_LC_21_14_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i83_LC_21_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i83_LC_21_14_4 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i83_LC_21_14_4  (
            .in0(N__68356),
            .in1(N__62499),
            .in2(N__69193),
            .in3(N__52539),
            .lcout(\c0.data_in_frame_10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66734),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1854_LC_21_14_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1854_LC_21_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1854_LC_21_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1854_LC_21_14_5  (
            .in0(N__58162),
            .in1(N__55118),
            .in2(_gnd_net_),
            .in3(N__57291),
            .lcout(\c0.n20402 ),
            .ltout(\c0.n20402_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1898_LC_21_14_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1898_LC_21_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1898_LC_21_14_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1898_LC_21_14_6  (
            .in0(N__57292),
            .in1(N__57325),
            .in2(N__52513),
            .in3(N__58216),
            .lcout(\c0.n21834 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i79_LC_21_14_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i79_LC_21_14_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i79_LC_21_14_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i79_LC_21_14_7  (
            .in0(N__62497),
            .in1(N__69883),
            .in2(N__52509),
            .in3(N__65670),
            .lcout(\c0.data_in_frame_9_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66734),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1333_LC_21_15_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1333_LC_21_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1333_LC_21_15_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1333_LC_21_15_0  (
            .in0(_gnd_net_),
            .in1(N__52475),
            .in2(_gnd_net_),
            .in3(N__57395),
            .lcout(\c0.n21873 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1720_LC_21_15_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1720_LC_21_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1720_LC_21_15_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1720_LC_21_15_1  (
            .in0(N__53656),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53695),
            .lcout(\c0.n22119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_LC_21_15_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_LC_21_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_LC_21_15_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_LC_21_15_3  (
            .in0(N__65761),
            .in1(N__52450),
            .in2(N__55027),
            .in3(N__60400),
            .lcout(),
            .ltout(\c0.n18_adj_4222_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_LC_21_15_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_LC_21_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_LC_21_15_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_LC_21_15_4  (
            .in0(N__52633),
            .in1(N__55668),
            .in2(N__52612),
            .in3(N__60103),
            .lcout(\c0.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i102_LC_21_15_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i102_LC_21_15_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i102_LC_21_15_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i102_LC_21_15_5  (
            .in0(N__64451),
            .in1(N__62428),
            .in2(N__60948),
            .in3(N__67171),
            .lcout(\c0.data_in_frame_12_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i76_LC_21_15_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i76_LC_21_15_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i76_LC_21_15_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i76_LC_21_15_6  (
            .in0(N__62427),
            .in1(N__57396),
            .in2(N__69877),
            .in3(N__64825),
            .lcout(\c0.data_in_frame_9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i122_LC_21_15_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i122_LC_21_15_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i122_LC_21_15_7 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \c0.data_in_frame_0__i122_LC_21_15_7  (
            .in0(N__63780),
            .in1(N__62429),
            .in2(N__68658),
            .in3(N__61382),
            .lcout(\c0.data_in_frame_15_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1217_LC_21_16_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1217_LC_21_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1217_LC_21_16_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1217_LC_21_16_0  (
            .in0(N__54796),
            .in1(N__52609),
            .in2(N__61360),
            .in3(N__52585),
            .lcout(\c0.n22003 ),
            .ltout(\c0.n22003_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1215_LC_21_16_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1215_LC_21_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1215_LC_21_16_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1215_LC_21_16_1  (
            .in0(N__52576),
            .in1(N__55210),
            .in2(N__52564),
            .in3(N__52561),
            .lcout(\c0.n6221 ),
            .ltout(\c0.n6221_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1216_LC_21_16_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1216_LC_21_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1216_LC_21_16_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1216_LC_21_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52555),
            .in3(N__55895),
            .lcout(\c0.n22084 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i150_LC_21_16_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i150_LC_21_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i150_LC_21_16_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i150_LC_21_16_4  (
            .in0(N__68093),
            .in1(N__69124),
            .in2(N__61579),
            .in3(N__67122),
            .lcout(\c0.data_in_frame_18_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66762),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i169_LC_21_16_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i169_LC_21_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i169_LC_21_16_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i169_LC_21_16_5  (
            .in0(N__62150),
            .in1(N__68094),
            .in2(N__55728),
            .in3(N__69537),
            .lcout(\c0.data_in_frame_21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66762),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1892_LC_21_16_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1892_LC_21_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1892_LC_21_16_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1892_LC_21_16_6  (
            .in0(N__55626),
            .in1(N__55557),
            .in2(N__64034),
            .in3(N__52552),
            .lcout(\c0.n22311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1866_LC_21_17_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1866_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1866_LC_21_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1866_LC_21_17_0  (
            .in0(N__58838),
            .in1(N__58691),
            .in2(_gnd_net_),
            .in3(N__59278),
            .lcout(\c0.n22099 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i205_LC_21_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i205_LC_21_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i205_LC_21_17_1 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i205_LC_21_17_1  (
            .in0(N__63107),
            .in1(N__53719),
            .in2(N__69882),
            .in3(N__67675),
            .lcout(\c0.data_in_frame_25_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66774),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1861_LC_21_17_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1861_LC_21_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1861_LC_21_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1861_LC_21_17_3  (
            .in0(N__54951),
            .in1(N__61747),
            .in2(_gnd_net_),
            .in3(N__58543),
            .lcout(),
            .ltout(\c0.n6_adj_4226_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1231_LC_21_17_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1231_LC_21_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1231_LC_21_17_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1231_LC_21_17_4  (
            .in0(N__53242),
            .in1(N__55156),
            .in2(N__53227),
            .in3(N__63357),
            .lcout(\c0.n23615 ),
            .ltout(\c0.n23615_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1232_LC_21_17_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1232_LC_21_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1232_LC_21_17_5 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \c0.i1_2_lut_adj_1232_LC_21_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53224),
            .in3(N__65073),
            .lcout(\c0.n22100 ),
            .ltout(\c0.n22100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1278_LC_21_17_6 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1278_LC_21_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1278_LC_21_17_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_1278_LC_21_17_6  (
            .in0(N__58278),
            .in1(N__53286),
            .in2(N__53221),
            .in3(N__53901),
            .lcout(\c0.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1226_LC_21_17_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1226_LC_21_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1226_LC_21_17_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1226_LC_21_17_7  (
            .in0(N__53217),
            .in1(N__55155),
            .in2(N__53206),
            .in3(N__58542),
            .lcout(\c0.n12594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1767_LC_21_18_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1767_LC_21_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1767_LC_21_18_0 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1767_LC_21_18_0  (
            .in0(N__52649),
            .in1(N__53196),
            .in2(_gnd_net_),
            .in3(N__53029),
            .lcout(\c0.n21366 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i20_LC_21_18_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i20_LC_21_18_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i20_LC_21_18_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i20_LC_21_18_1  (
            .in0(_gnd_net_),
            .in1(N__52650),
            .in2(_gnd_net_),
            .in3(N__52867),
            .lcout(\c0.FRAME_MATCHER_state_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66788),
            .ce(),
            .sr(N__53518));
    defparam \c0.i2_3_lut_LC_21_18_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_LC_21_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_LC_21_18_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_3_lut_LC_21_18_5  (
            .in0(N__53810),
            .in1(N__53786),
            .in2(_gnd_net_),
            .in3(N__55535),
            .lcout(\c0.n21043 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1455_LC_21_18_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1455_LC_21_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1455_LC_21_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1455_LC_21_18_7  (
            .in0(N__53503),
            .in1(N__53475),
            .in2(_gnd_net_),
            .in3(N__53416),
            .lcout(\c0.n13379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_LC_21_19_0 .C_ON=1'b0;
    defparam \c0.i11_4_lut_LC_21_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_LC_21_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_LC_21_19_0  (
            .in0(N__55228),
            .in1(N__53862),
            .in2(N__53335),
            .in3(N__55753),
            .lcout(),
            .ltout(\c0.n28_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_LC_21_19_1 .C_ON=1'b0;
    defparam \c0.i16_4_lut_LC_21_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_LC_21_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_LC_21_19_1  (
            .in0(N__62839),
            .in1(N__55261),
            .in2(N__53302),
            .in3(N__55678),
            .lcout(\c0.n23640 ),
            .ltout(\c0.n23640_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1903_LC_21_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1903_LC_21_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1903_LC_21_19_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1903_LC_21_19_2  (
            .in0(N__60489),
            .in1(_gnd_net_),
            .in2(N__53299),
            .in3(N__53292),
            .lcout(\c0.n22197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_LC_21_19_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_LC_21_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_LC_21_19_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_4_lut_LC_21_19_3  (
            .in0(N__55485),
            .in1(N__53256),
            .in2(N__57972),
            .in3(N__55684),
            .lcout(\c0.n22305 ),
            .ltout(\c0.n22305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1901_LC_21_19_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1901_LC_21_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1901_LC_21_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1901_LC_21_19_4  (
            .in0(_gnd_net_),
            .in1(N__60340),
            .in2(N__53296),
            .in3(N__60312),
            .lcout(\c0.n20137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_LC_21_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_LC_21_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_LC_21_19_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i1_2_lut_LC_21_19_5  (
            .in0(N__53293),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53257),
            .lcout(\c0.n21208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1200_LC_21_19_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1200_LC_21_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1200_LC_21_19_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1200_LC_21_19_6  (
            .in0(_gnd_net_),
            .in1(N__53848),
            .in2(_gnd_net_),
            .in3(N__53248),
            .lcout(),
            .ltout(\c0.n6_adj_4219_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1201_LC_21_19_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1201_LC_21_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1201_LC_21_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1201_LC_21_19_7  (
            .in0(N__60313),
            .in1(N__63257),
            .in2(N__53821),
            .in3(N__64257),
            .lcout(\c0.n21160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1902_LC_21_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1902_LC_21_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1902_LC_21_20_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1902_LC_21_20_0  (
            .in0(N__53817),
            .in1(N__53787),
            .in2(N__53727),
            .in3(N__55539),
            .lcout(\c0.n21949 ),
            .ltout(\c0.n21949_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1191_LC_21_20_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1191_LC_21_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1191_LC_21_20_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_3_lut_adj_1191_LC_21_20_1  (
            .in0(N__53650),
            .in1(_gnd_net_),
            .in2(N__53770),
            .in3(N__53762),
            .lcout(\c0.n23009 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1736_LC_21_20_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1736_LC_21_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1736_LC_21_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1736_LC_21_20_2  (
            .in0(N__53690),
            .in1(N__59541),
            .in2(N__53766),
            .in3(N__64189),
            .lcout(\c0.n22157 ),
            .ltout(\c0.n22157_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1733_LC_21_20_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1733_LC_21_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1733_LC_21_20_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_1733_LC_21_20_3  (
            .in0(N__58899),
            .in1(N__55807),
            .in2(N__53746),
            .in3(N__54130),
            .lcout(\c0.n20846 ),
            .ltout(\c0.n20846_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1734_LC_21_20_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1734_LC_21_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1734_LC_21_20_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i5_4_lut_adj_1734_LC_21_20_4  (
            .in0(N__54131),
            .in1(N__54008),
            .in2(N__53731),
            .in3(N__55794),
            .lcout(\c0.n12_adj_4491 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1655_LC_21_20_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1655_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1655_LC_21_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1655_LC_21_20_5  (
            .in0(N__53720),
            .in1(N__53689),
            .in2(N__53655),
            .in3(N__53599),
            .lcout(\c0.n22370 ),
            .ltout(\c0.n22370_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1735_LC_21_20_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1735_LC_21_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1735_LC_21_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1735_LC_21_20_6  (
            .in0(N__53548),
            .in1(N__53542),
            .in2(N__53536),
            .in3(N__56080),
            .lcout(\c0.n23356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1194_LC_21_21_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1194_LC_21_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1194_LC_21_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1194_LC_21_21_2  (
            .in0(N__53827),
            .in1(N__66097),
            .in2(_gnd_net_),
            .in3(N__54015),
            .lcout(\c0.n22145 ),
            .ltout(\c0.n22145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1381_LC_21_21_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1381_LC_21_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1381_LC_21_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1381_LC_21_21_3  (
            .in0(N__58614),
            .in1(N__53980),
            .in2(N__53968),
            .in3(N__66135),
            .lcout(\c0.n10_adj_4297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i238_LC_21_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i238_LC_21_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i238_LC_21_21_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i238_LC_21_21_4  (
            .in0(N__67705),
            .in1(N__62167),
            .in2(N__56308),
            .in3(N__67079),
            .lcout(\c0.data_in_frame_29_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66820),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1383_LC_21_21_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1383_LC_21_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1383_LC_21_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1383_LC_21_21_5  (
            .in0(N__59542),
            .in1(N__64588),
            .in2(N__59365),
            .in3(N__56065),
            .lcout(),
            .ltout(\c0.n23335_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1387_LC_21_21_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1387_LC_21_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1387_LC_21_21_6 .LUT_INIT=16'b0110111110011111;
    LogicCell40 \c0.i3_4_lut_adj_1387_LC_21_21_6  (
            .in0(N__53916),
            .in1(N__53965),
            .in2(N__53959),
            .in3(N__58717),
            .lcout(\c0.n21_adj_4300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i236_LC_21_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i236_LC_21_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i236_LC_21_21_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i236_LC_21_21_7  (
            .in0(N__62166),
            .in1(N__64887),
            .in2(N__53940),
            .in3(N__67706),
            .lcout(\c0.data_in_frame_29_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66820),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i225_LC_21_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i225_LC_21_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i225_LC_21_22_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i225_LC_21_22_1  (
            .in0(N__67751),
            .in1(N__64565),
            .in2(N__53920),
            .in3(N__69538),
            .lcout(\c0.data_in_frame_28_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66832),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1196_LC_21_22_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1196_LC_21_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1196_LC_21_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1196_LC_21_22_2  (
            .in0(N__53905),
            .in1(N__65428),
            .in2(N__55729),
            .in3(N__53866),
            .lcout(\c0.n22040 ),
            .ltout(\c0.n22040_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1193_LC_21_22_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1193_LC_21_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1193_LC_21_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1193_LC_21_22_3  (
            .in0(N__67818),
            .in1(N__64228),
            .in2(N__53839),
            .in3(N__53836),
            .lcout(\c0.n21099 ),
            .ltout(\c0.n21099_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1718_LC_21_22_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1718_LC_21_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1718_LC_21_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1718_LC_21_22_4  (
            .in0(N__54148),
            .in1(N__55829),
            .in2(N__54139),
            .in3(N__54136),
            .lcout(\c0.n22148 ),
            .ltout(\c0.n22148_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1377_LC_21_22_5 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1377_LC_21_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1377_LC_21_22_5 .LUT_INIT=16'b1110110111011110;
    LogicCell40 \c0.i8_4_lut_adj_1377_LC_21_22_5  (
            .in0(N__54111),
            .in1(N__54097),
            .in2(N__54079),
            .in3(N__54076),
            .lcout(\c0.n26_adj_4294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i173_LC_21_23_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i173_LC_21_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i173_LC_21_23_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i173_LC_21_23_0  (
            .in0(N__62160),
            .in1(N__68141),
            .in2(N__58337),
            .in3(N__63000),
            .lcout(\c0.data_in_frame_21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66844),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_1178_LC_21_23_1 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_1178_LC_21_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_1178_LC_21_23_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.rx.i1_2_lut_adj_1178_LC_21_23_1  (
            .in0(_gnd_net_),
            .in1(N__59749),
            .in2(_gnd_net_),
            .in3(N__56160),
            .lcout(n12977),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_LC_21_23_5 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_LC_21_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_LC_21_23_5 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_4_lut_LC_21_23_5  (
            .in0(N__56991),
            .in1(N__56808),
            .in2(N__56910),
            .in3(N__57054),
            .lcout(\c0.rx.n12862 ),
            .ltout(\c0.rx.n12862_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_1175_LC_21_23_6 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_1175_LC_21_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_1175_LC_21_23_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \c0.rx.i1_2_lut_adj_1175_LC_21_23_6  (
            .in0(N__59748),
            .in1(_gnd_net_),
            .in2(N__54058),
            .in3(_gnd_net_),
            .lcout(n12973),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_adj_1171_LC_21_24_1 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_adj_1171_LC_21_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_adj_1171_LC_21_24_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.rx.i2_3_lut_adj_1171_LC_21_24_1  (
            .in0(N__54054),
            .in1(N__54042),
            .in2(_gnd_net_),
            .in3(N__54030),
            .lcout(\c0.rx.n80 ),
            .ltout(\c0.rx.n80_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_LC_21_24_2 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_LC_21_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_LC_21_24_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \c0.rx.i1_4_lut_LC_21_24_2  (
            .in0(N__54283),
            .in1(N__54319),
            .in2(N__54019),
            .in3(N__54300),
            .lcout(r_SM_Main_2_N_3681_2),
            .ltout(r_SM_Main_2_N_3681_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_4_lut_LC_21_24_3.C_ON=1'b0;
    defparam i13_4_lut_4_lut_LC_21_24_3.SEQ_MODE=4'b0000;
    defparam i13_4_lut_4_lut_LC_21_24_3.LUT_INIT=16'b0010000001010101;
    LogicCell40 i13_4_lut_4_lut_LC_21_24_3 (
            .in0(N__56889),
            .in1(N__56993),
            .in2(N__54346),
            .in3(N__56818),
            .lcout(n14283),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i2_LC_21_24_5 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i2_LC_21_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i2_LC_21_24_5 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \c0.rx.r_SM_Main_i2_LC_21_24_5  (
            .in0(N__54320),
            .in1(N__54301),
            .in2(N__54289),
            .in3(N__54262),
            .lcout(r_SM_Main_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66852),
            .ce(),
            .sr(N__54250));
    defparam \c0.rx.r_Rx_Data_50_LC_22_7_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_50_LC_22_7_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_50_LC_22_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.rx.r_Rx_Data_50_LC_22_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54232),
            .lcout(r_Rx_Data),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66663),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i103_LC_22_8_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i103_LC_22_8_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i103_LC_22_8_1 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i103_LC_22_8_1  (
            .in0(N__65623),
            .in1(N__62432),
            .in2(N__54213),
            .in3(N__64346),
            .lcout(\c0.data_in_frame_12_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66670),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i124_LC_22_8_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i124_LC_22_8_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i124_LC_22_8_2 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_in_frame_0__i124_LC_22_8_2  (
            .in0(N__62431),
            .in1(N__68516),
            .in2(N__64892),
            .in3(N__54189),
            .lcout(\c0.data_in_frame_15_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66670),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1286_LC_22_8_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1286_LC_22_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1286_LC_22_8_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1286_LC_22_8_3  (
            .in0(N__54528),
            .in1(N__59245),
            .in2(N__56767),
            .in3(N__57909),
            .lcout(\c0.n22424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1242_LC_22_8_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1242_LC_22_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1242_LC_22_8_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1242_LC_22_8_4  (
            .in0(_gnd_net_),
            .in1(N__61389),
            .in2(_gnd_net_),
            .in3(N__54188),
            .lcout(\c0.n22430 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i133_LC_22_8_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i133_LC_22_8_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i133_LC_22_8_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i133_LC_22_8_5  (
            .in0(N__66007),
            .in1(N__68166),
            .in2(N__57324),
            .in3(N__63177),
            .lcout(\c0.data_in_frame_16_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66670),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1267_LC_22_9_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1267_LC_22_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1267_LC_22_9_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1267_LC_22_9_0  (
            .in0(_gnd_net_),
            .in1(N__54447),
            .in2(_gnd_net_),
            .in3(N__54164),
            .lcout(),
            .ltout(\c0.n6_adj_4244_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1268_LC_22_9_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1268_LC_22_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1268_LC_22_9_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1268_LC_22_9_1  (
            .in0(N__54541),
            .in1(N__57175),
            .in2(N__54532),
            .in3(N__54529),
            .lcout(\c0.n20240 ),
            .ltout(\c0.n20240_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1309_LC_22_9_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1309_LC_22_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1309_LC_22_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1309_LC_22_9_2  (
            .in0(_gnd_net_),
            .in1(N__58137),
            .in2(N__54514),
            .in3(N__57313),
            .lcout(\c0.n22385 ),
            .ltout(\c0.n22385_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1246_LC_22_9_3 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1246_LC_22_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1246_LC_22_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_1246_LC_22_9_3  (
            .in0(N__55219),
            .in1(N__54511),
            .in2(N__54481),
            .in3(N__61467),
            .lcout(\c0.n29_adj_4234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i118_LC_22_9_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i118_LC_22_9_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i118_LC_22_9_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i118_LC_22_9_4  (
            .in0(N__67123),
            .in1(N__57157),
            .in2(_gnd_net_),
            .in3(N__54467),
            .lcout(data_in_frame_14_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66680),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i80_LC_22_9_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i80_LC_22_9_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i80_LC_22_9_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i80_LC_22_9_5  (
            .in0(N__62377),
            .in1(N__69716),
            .in2(N__57370),
            .in3(N__68867),
            .lcout(\c0.data_in_frame_9_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66680),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i116_LC_22_10_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i116_LC_22_10_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i116_LC_22_10_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i116_LC_22_10_1  (
            .in0(N__64863),
            .in1(N__57158),
            .in2(_gnd_net_),
            .in3(N__54448),
            .lcout(data_in_frame_14_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66693),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i13_LC_22_10_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i13_LC_22_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i13_LC_22_10_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i13_LC_22_10_2  (
            .in0(N__63175),
            .in1(N__69871),
            .in2(N__54407),
            .in3(N__60898),
            .lcout(data_in_frame_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66693),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1548_LC_22_10_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1548_LC_22_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1548_LC_22_10_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1548_LC_22_10_3  (
            .in0(_gnd_net_),
            .in1(N__54432),
            .in2(_gnd_net_),
            .in3(N__54395),
            .lcout(\c0.n21797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i181_LC_22_10_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i181_LC_22_10_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i181_LC_22_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i181_LC_22_10_4  (
            .in0(N__63174),
            .in1(N__59811),
            .in2(_gnd_net_),
            .in3(N__59198),
            .lcout(data_in_frame_22_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66693),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1269_LC_22_10_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1269_LC_22_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1269_LC_22_10_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1269_LC_22_10_5  (
            .in0(N__57345),
            .in1(N__59581),
            .in2(N__57253),
            .in3(N__54778),
            .lcout(),
            .ltout(\c0.n10_adj_4245_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1853_LC_22_10_6 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1853_LC_22_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1853_LC_22_10_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1853_LC_22_10_6  (
            .in0(N__54751),
            .in1(N__54718),
            .in2(N__54688),
            .in3(N__54684),
            .lcout(\c0.n13598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i119_LC_22_10_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i119_LC_22_10_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i119_LC_22_10_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i119_LC_22_10_7  (
            .in0(N__65624),
            .in1(N__57159),
            .in2(_gnd_net_),
            .in3(N__55095),
            .lcout(data_in_frame_14_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66693),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1291_LC_22_11_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1291_LC_22_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1291_LC_22_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1291_LC_22_11_1  (
            .in0(N__60574),
            .in1(N__54634),
            .in2(_gnd_net_),
            .in3(N__54613),
            .lcout(\c0.n22233 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i127_LC_22_11_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i127_LC_22_11_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i127_LC_22_11_2 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_in_frame_0__i127_LC_22_11_2  (
            .in0(N__62538),
            .in1(N__68601),
            .in2(N__65696),
            .in3(N__57870),
            .lcout(\c0.data_in_frame_15_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66706),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i92_LC_22_11_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i92_LC_22_11_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i92_LC_22_11_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i92_LC_22_11_3  (
            .in0(N__67477),
            .in1(N__62540),
            .in2(N__54592),
            .in3(N__64862),
            .lcout(\c0.data_in_frame_11_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66706),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1340_LC_22_11_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1340_LC_22_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1340_LC_22_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1340_LC_22_11_4  (
            .in0(N__54587),
            .in1(N__54571),
            .in2(_gnd_net_),
            .in3(N__54565),
            .lcout(\c0.n4_adj_4240 ),
            .ltout(\c0.n4_adj_4240_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_4_lut_LC_22_11_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_4_lut_LC_22_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_4_lut_LC_22_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_4_lut_4_lut_LC_22_11_5  (
            .in0(_gnd_net_),
            .in1(N__57817),
            .in2(N__54544),
            .in3(N__57584),
            .lcout(\c0.n22781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1784_LC_22_11_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1784_LC_22_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1784_LC_22_11_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1784_LC_22_11_6  (
            .in0(N__57585),
            .in1(N__57217),
            .in2(N__61894),
            .in3(N__59580),
            .lcout(\c0.n21126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i110_LC_22_11_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i110_LC_22_11_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i110_LC_22_11_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i110_LC_22_11_7  (
            .in0(N__67124),
            .in1(N__62539),
            .in2(N__62149),
            .in3(N__61289),
            .lcout(\c0.data_in_frame_13_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66706),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i94_LC_22_12_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i94_LC_22_12_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i94_LC_22_12_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i94_LC_22_12_0  (
            .in0(N__67445),
            .in1(N__62500),
            .in2(N__57679),
            .in3(N__67157),
            .lcout(\c0.data_in_frame_11_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66721),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i120_LC_22_12_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i120_LC_22_12_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i120_LC_22_12_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i120_LC_22_12_1  (
            .in0(N__68865),
            .in1(N__57166),
            .in2(_gnd_net_),
            .in3(N__55057),
            .lcout(data_in_frame_14_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66721),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i202_LC_22_12_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i202_LC_22_12_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i202_LC_22_12_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i202_LC_22_12_2  (
            .in0(N__63826),
            .in1(N__69872),
            .in2(N__56138),
            .in3(N__67776),
            .lcout(\c0.data_in_frame_25_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66721),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1289_LC_22_12_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1289_LC_22_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1289_LC_22_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1289_LC_22_12_3  (
            .in0(N__57843),
            .in1(N__60937),
            .in2(_gnd_net_),
            .in3(N__57582),
            .lcout(\c0.n22236 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1335_LC_22_12_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1335_LC_22_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1335_LC_22_12_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1335_LC_22_12_4  (
            .in0(_gnd_net_),
            .in1(N__57674),
            .in2(_gnd_net_),
            .in3(N__54889),
            .lcout(\c0.n6_adj_4273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1264_LC_22_12_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1264_LC_22_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1264_LC_22_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1264_LC_22_12_5  (
            .in0(N__54853),
            .in1(N__60996),
            .in2(N__54847),
            .in3(N__54828),
            .lcout(\c0.n21982 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1293_LC_22_12_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1293_LC_22_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1293_LC_22_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1293_LC_22_12_6  (
            .in0(_gnd_net_),
            .in1(N__57842),
            .in2(_gnd_net_),
            .in3(N__55137),
            .lcout(\c0.n5813 ),
            .ltout(\c0.n5813_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1295_LC_22_12_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1295_LC_22_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1295_LC_22_12_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1295_LC_22_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__54799),
            .in3(N__54906),
            .lcout(\c0.n13728 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1223_LC_22_13_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1223_LC_22_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1223_LC_22_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1223_LC_22_13_0  (
            .in0(N__55097),
            .in1(N__54795),
            .in2(N__65404),
            .in3(N__54937),
            .lcout(\c0.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1338_LC_22_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1338_LC_22_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1338_LC_22_13_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1338_LC_22_13_1  (
            .in0(_gnd_net_),
            .in1(N__57583),
            .in2(_gnd_net_),
            .in3(N__57540),
            .lcout(),
            .ltout(\c0.n20222_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1243_LC_22_13_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1243_LC_22_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1243_LC_22_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1243_LC_22_13_2  (
            .in0(N__54927),
            .in1(N__60450),
            .in2(N__55018),
            .in3(N__55011),
            .lcout(),
            .ltout(\c0.n28_adj_4232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_3_lut_4_lut_adj_1858_LC_22_13_3 .C_ON=1'b0;
    defparam \c0.i14_3_lut_4_lut_adj_1858_LC_22_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_3_lut_4_lut_adj_1858_LC_22_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_3_lut_4_lut_adj_1858_LC_22_13_3  (
            .in0(N__58029),
            .in1(N__55096),
            .in2(N__54985),
            .in3(N__55047),
            .lcout(),
            .ltout(\c0.n32_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_LC_22_13_4 .C_ON=1'b0;
    defparam \c0.i17_4_lut_LC_22_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_LC_22_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_LC_22_13_4  (
            .in0(N__57199),
            .in1(N__57823),
            .in2(N__54982),
            .in3(N__54979),
            .lcout(\c0.n21238 ),
            .ltout(\c0.n21238_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_LC_22_13_5 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_LC_22_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_LC_22_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_3_lut_4_lut_LC_22_13_5  (
            .in0(N__65759),
            .in1(N__54970),
            .in2(N__54958),
            .in3(N__54955),
            .lcout(\c0.n8_adj_4236 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1392_LC_22_13_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1392_LC_22_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1392_LC_22_13_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1392_LC_22_13_6  (
            .in0(N__58172),
            .in1(N__65760),
            .in2(_gnd_net_),
            .in3(N__54936),
            .lcout(\c0.n21831 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i147_LC_22_14_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i147_LC_22_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i147_LC_22_14_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i147_LC_22_14_0  (
            .in0(N__69205),
            .in1(N__68111),
            .in2(N__57796),
            .in3(N__68357),
            .lcout(\c0.data_in_frame_18_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66748),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1228_LC_22_14_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1228_LC_22_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1228_LC_22_14_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1228_LC_22_14_2  (
            .in0(N__54928),
            .in1(N__57529),
            .in2(N__55065),
            .in3(N__61156),
            .lcout(\c0.n22480 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1238_LC_22_14_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1238_LC_22_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1238_LC_22_14_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1238_LC_22_14_3  (
            .in0(N__60030),
            .in1(N__61322),
            .in2(N__58498),
            .in3(N__54910),
            .lcout(\c0.n13719 ),
            .ltout(\c0.n13719_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1249_LC_22_14_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1249_LC_22_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1249_LC_22_14_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1249_LC_22_14_4  (
            .in0(N__61177),
            .in1(N__61824),
            .in2(N__55144),
            .in3(N__55141),
            .lcout(\c0.n14_adj_4238 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i149_LC_22_14_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i149_LC_22_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i149_LC_22_14_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i149_LC_22_14_5  (
            .in0(N__68109),
            .in1(N__69206),
            .in2(N__58236),
            .in3(N__63146),
            .lcout(\c0.data_in_frame_18_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66748),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i145_LC_22_14_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i145_LC_22_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i145_LC_22_14_6 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i145_LC_22_14_6  (
            .in0(N__69482),
            .in1(N__68110),
            .in2(N__69233),
            .in3(N__57756),
            .lcout(\c0.data_in_frame_18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66748),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1262_LC_22_14_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1262_LC_22_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1262_LC_22_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1262_LC_22_14_7  (
            .in0(_gnd_net_),
            .in1(N__55119),
            .in2(_gnd_net_),
            .in3(N__57284),
            .lcout(\c0.n20374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_1676_LC_22_15_0 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_1676_LC_22_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_1676_LC_22_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_1676_LC_22_15_0  (
            .in0(N__63918),
            .in1(N__63956),
            .in2(N__56014),
            .in3(N__55509),
            .lcout(\c0.n21067 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1233_LC_22_15_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1233_LC_22_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1233_LC_22_15_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1233_LC_22_15_1  (
            .in0(_gnd_net_),
            .in1(N__61763),
            .in2(_gnd_net_),
            .in3(N__61737),
            .lcout(\c0.n22113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3317_2_lut_LC_22_15_2 .C_ON=1'b0;
    defparam \c0.i3317_2_lut_LC_22_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3317_2_lut_LC_22_15_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3317_2_lut_LC_22_15_2  (
            .in0(_gnd_net_),
            .in1(N__55101),
            .in2(_gnd_net_),
            .in3(N__55066),
            .lcout(\c0.n5996 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i134_LC_22_15_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i134_LC_22_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i134_LC_22_15_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i134_LC_22_15_3  (
            .in0(N__65937),
            .in1(N__68162),
            .in2(N__58174),
            .in3(N__67170),
            .lcout(\c0.data_in_frame_16_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66763),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i195_LC_22_15_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i195_LC_22_15_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i195_LC_22_15_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i195_LC_22_15_4  (
            .in0(N__68417),
            .in1(N__65938),
            .in2(N__65192),
            .in3(N__67756),
            .lcout(\c0.data_in_frame_24_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66763),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i131_LC_22_15_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i131_LC_22_15_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i131_LC_22_15_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i131_LC_22_15_5  (
            .in0(N__65936),
            .in1(N__68161),
            .in2(N__58099),
            .in3(N__68418),
            .lcout(\c0.data_in_frame_16_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66763),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i163_LC_22_15_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i163_LC_22_15_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i163_LC_22_15_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i163_LC_22_15_7  (
            .in0(N__64517),
            .in1(N__68163),
            .in2(N__61773),
            .in3(N__68419),
            .lcout(\c0.data_in_frame_20_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66763),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i140_LC_22_16_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i140_LC_22_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i140_LC_22_16_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i140_LC_22_16_0  (
            .in0(N__69867),
            .in1(N__68043),
            .in2(N__55429),
            .in3(N__64748),
            .lcout(\c0.data_in_frame_17_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_LC_22_16_1 .C_ON=1'b0;
    defparam \c0.i2_4_lut_LC_22_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_LC_22_16_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_LC_22_16_1  (
            .in0(N__64152),
            .in1(N__55249),
            .in2(N__60037),
            .in3(N__55240),
            .lcout(\c0.n20203 ),
            .ltout(\c0.n20203_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1255_LC_22_16_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1255_LC_22_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1255_LC_22_16_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1255_LC_22_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__55231),
            .in3(N__61745),
            .lcout(\c0.n21120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i148_LC_22_16_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i148_LC_22_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i148_LC_22_16_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i148_LC_22_16_3  (
            .in0(N__68042),
            .in1(N__69210),
            .in2(N__64819),
            .in3(N__62900),
            .lcout(\c0.data_in_frame_18_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i125_LC_22_16_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i125_LC_22_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i125_LC_22_16_4 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \c0.data_in_frame_0__i125_LC_22_16_4  (
            .in0(N__63218),
            .in1(N__62505),
            .in2(N__68659),
            .in3(N__58483),
            .lcout(\c0.data_in_frame_15_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i123_LC_22_16_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i123_LC_22_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i123_LC_22_16_6 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i123_LC_22_16_6  (
            .in0(N__68628),
            .in1(N__62504),
            .in2(N__55218),
            .in3(N__68288),
            .lcout(\c0.data_in_frame_15_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1227_LC_22_16_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1227_LC_22_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1227_LC_22_16_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1227_LC_22_16_7  (
            .in0(N__57489),
            .in1(N__55183),
            .in2(N__55171),
            .in3(N__55641),
            .lcout(\c0.n20196 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1719_LC_22_17_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1719_LC_22_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1719_LC_22_17_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_1719_LC_22_17_0  (
            .in0(N__65153),
            .in1(N__55447),
            .in2(N__59797),
            .in3(N__59279),
            .lcout(\c0.n21054 ),
            .ltout(\c0.n21054_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1722_LC_22_17_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1722_LC_22_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1722_LC_22_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1722_LC_22_17_1  (
            .in0(N__62631),
            .in1(N__58972),
            .in2(N__55441),
            .in3(N__55438),
            .lcout(\c0.n14_adj_4484 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4028_2_lut_LC_22_17_2 .C_ON=1'b0;
    defparam \c0.i4028_2_lut_LC_22_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4028_2_lut_LC_22_17_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i4028_2_lut_LC_22_17_2  (
            .in0(N__59534),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59401),
            .lcout(\c0.n6707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1884_LC_22_17_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1884_LC_22_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1884_LC_22_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1884_LC_22_17_3  (
            .in0(N__59400),
            .in1(N__59533),
            .in2(N__63475),
            .in3(N__65230),
            .lcout(\c0.n22323 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1229_LC_22_17_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1229_LC_22_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1229_LC_22_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1229_LC_22_17_4  (
            .in0(N__55417),
            .in1(N__55394),
            .in2(_gnd_net_),
            .in3(N__55350),
            .lcout(\c0.n12596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1750_LC_22_17_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1750_LC_22_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1750_LC_22_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1750_LC_22_17_5  (
            .in0(N__55351),
            .in1(N__55339),
            .in2(_gnd_net_),
            .in3(N__55302),
            .lcout(\c0.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_LC_22_18_0 .C_ON=1'b0;
    defparam \c0.i13_4_lut_LC_22_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_LC_22_18_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_LC_22_18_0  (
            .in0(N__61848),
            .in1(N__55282),
            .in2(N__55276),
            .in3(N__55497),
            .lcout(\c0.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1661_LC_22_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1661_LC_22_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1661_LC_22_18_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1661_LC_22_18_2  (
            .in0(N__55964),
            .in1(N__55896),
            .in2(N__58846),
            .in3(N__58692),
            .lcout(\c0.n20266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1280_LC_22_18_3 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1280_LC_22_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1280_LC_22_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1280_LC_22_18_3  (
            .in0(N__55534),
            .in1(N__55255),
            .in2(N__62598),
            .in3(N__58504),
            .lcout(\c0.n23062 ),
            .ltout(\c0.n23062_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1282_LC_22_18_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1282_LC_22_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1282_LC_22_18_4 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.i5_3_lut_adj_1282_LC_22_18_4  (
            .in0(N__55749),
            .in1(_gnd_net_),
            .in2(N__55732),
            .in3(N__55724),
            .lcout(\c0.n14_adj_4251 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_1399_LC_22_18_6 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_1399_LC_22_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_1399_LC_22_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_1399_LC_22_18_6  (
            .in0(N__58429),
            .in1(N__55690),
            .in2(N__55945),
            .in3(N__58741),
            .lcout(\c0.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_LC_22_19_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_LC_22_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_LC_22_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_LC_22_19_0  (
            .in0(N__55564),
            .in1(N__61435),
            .in2(N__63957),
            .in3(N__58459),
            .lcout(\c0.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1222_LC_22_19_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1222_LC_22_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1222_LC_22_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1222_LC_22_19_1  (
            .in0(N__55672),
            .in1(N__60947),
            .in2(N__63421),
            .in3(N__55645),
            .lcout(),
            .ltout(\c0.n16_adj_4223_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1224_LC_22_19_2 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1224_LC_22_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1224_LC_22_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1224_LC_22_19_2  (
            .in0(N__55625),
            .in1(N__58189),
            .in2(N__55576),
            .in3(N__55573),
            .lcout(\c0.n22211 ),
            .ltout(\c0.n22211_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1225_LC_22_19_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1225_LC_22_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1225_LC_22_19_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i2_3_lut_adj_1225_LC_22_19_3  (
            .in0(_gnd_net_),
            .in1(N__55563),
            .in2(N__55543),
            .in3(N__64069),
            .lcout(\c0.n21140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1207_LC_22_19_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1207_LC_22_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1207_LC_22_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1207_LC_22_19_5  (
            .in0(N__56010),
            .in1(N__55513),
            .in2(_gnd_net_),
            .in3(N__55498),
            .lcout(\c0.n23298 ),
            .ltout(\c0.n23298_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1208_LC_22_19_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1208_LC_22_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1208_LC_22_19_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1208_LC_22_19_6  (
            .in0(N__55471),
            .in1(N__58341),
            .in2(N__55462),
            .in3(N__58426),
            .lcout(\c0.n21200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_4_lut_adj_1729_LC_22_20_0 .C_ON=1'b0;
    defparam \c0.i23_4_lut_adj_1729_LC_22_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i23_4_lut_adj_1729_LC_22_20_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i23_4_lut_adj_1729_LC_22_20_0  (
            .in0(N__55459),
            .in1(N__57952),
            .in2(N__55840),
            .in3(N__59067),
            .lcout(),
            .ltout(\c0.n52_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i26_4_lut_adj_1732_LC_22_20_1 .C_ON=1'b0;
    defparam \c0.i26_4_lut_adj_1732_LC_22_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i26_4_lut_adj_1732_LC_22_20_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i26_4_lut_adj_1732_LC_22_20_1  (
            .in0(N__63547),
            .in1(N__58898),
            .in2(N__55810),
            .in3(N__55774),
            .lcout(\c0.n55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1738_LC_22_20_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1738_LC_22_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1738_LC_22_20_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1738_LC_22_20_2  (
            .in0(_gnd_net_),
            .in1(N__58644),
            .in2(_gnd_net_),
            .in3(N__59393),
            .lcout(\c0.n13872 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1653_LC_22_20_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1653_LC_22_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1653_LC_22_20_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1653_LC_22_20_4  (
            .in0(N__58897),
            .in1(N__58645),
            .in2(N__59408),
            .in3(N__59019),
            .lcout(\c0.n12420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i199_LC_22_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i199_LC_22_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i199_LC_22_20_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i199_LC_22_20_5  (
            .in0(N__67758),
            .in1(N__65575),
            .in2(N__59407),
            .in3(N__65939),
            .lcout(\c0.data_in_frame_24_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66821),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1199_LC_22_20_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1199_LC_22_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1199_LC_22_20_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_1199_LC_22_20_6  (
            .in0(_gnd_net_),
            .in1(N__61642),
            .in2(_gnd_net_),
            .in3(N__55783),
            .lcout(\c0.n22468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_3_lut_4_lut_LC_22_20_7 .C_ON=1'b0;
    defparam \c0.i15_3_lut_4_lut_LC_22_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15_3_lut_4_lut_LC_22_20_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_3_lut_4_lut_LC_22_20_7  (
            .in0(N__62791),
            .in1(N__58713),
            .in2(N__58845),
            .in3(N__59289),
            .lcout(\c0.n44_adj_4490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_1725_LC_22_21_0 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_1725_LC_22_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_1725_LC_22_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_adj_1725_LC_22_21_0  (
            .in0(N__69280),
            .in1(N__58896),
            .in2(N__66096),
            .in3(N__59079),
            .lcout(),
            .ltout(\c0.n48_adj_4485_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_LC_22_21_1 .C_ON=1'b0;
    defparam \c0.i24_4_lut_LC_22_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_LC_22_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i24_4_lut_LC_22_21_1  (
            .in0(N__58561),
            .in1(N__56020),
            .in2(N__55768),
            .in3(N__66908),
            .lcout(\c0.n53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1371_LC_22_21_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1371_LC_22_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1371_LC_22_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1371_LC_22_21_2  (
            .in0(N__55938),
            .in1(N__66128),
            .in2(N__65275),
            .in3(N__55765),
            .lcout(\c0.n22719 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1654_LC_22_21_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1654_LC_22_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1654_LC_22_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1654_LC_22_21_3  (
            .in0(N__56142),
            .in1(N__63490),
            .in2(_gnd_net_),
            .in3(N__65247),
            .lcout(\c0.n20370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i28_4_lut_LC_22_21_4 .C_ON=1'b0;
    defparam \c0.i28_4_lut_LC_22_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i28_4_lut_LC_22_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i28_4_lut_LC_22_21_4  (
            .in0(N__56107),
            .in1(N__56092),
            .in2(N__58570),
            .in3(N__56086),
            .lcout(\c0.n23416 ),
            .ltout(\c0.n23416_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1380_LC_22_21_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1380_LC_22_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1380_LC_22_21_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i5_4_lut_adj_1380_LC_22_21_5  (
            .in0(N__59080),
            .in1(N__63439),
            .in2(N__56068),
            .in3(N__59071),
            .lcout(\c0.n12_adj_4296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_4_lut_adj_1829_LC_22_22_0 .C_ON=1'b0;
    defparam \c0.i7_3_lut_4_lut_adj_1829_LC_22_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_4_lut_adj_1829_LC_22_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_3_lut_4_lut_adj_1829_LC_22_22_0  (
            .in0(N__55966),
            .in1(N__56053),
            .in2(N__56283),
            .in3(N__55846),
            .lcout(\c0.n36_adj_4489 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1659_LC_22_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1659_LC_22_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1659_LC_22_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1659_LC_22_22_2  (
            .in0(N__55999),
            .in1(N__55890),
            .in2(N__58836),
            .in3(N__63900),
            .lcout(\c0.n22388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1782_LC_22_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1782_LC_22_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1782_LC_22_22_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1782_LC_22_22_3  (
            .in0(N__63901),
            .in1(N__55965),
            .in2(N__55897),
            .in3(N__63958),
            .lcout(\c0.n21037 ),
            .ltout(\c0.n21037_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1391_LC_22_22_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1391_LC_22_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1391_LC_22_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1391_LC_22_22_4  (
            .in0(N__58327),
            .in1(N__55924),
            .in2(N__55900),
            .in3(N__58427),
            .lcout(\c0.n13993 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1236_LC_22_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1236_LC_22_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1236_LC_22_22_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1236_LC_22_22_5  (
            .in0(N__55894),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58822),
            .lcout(\c0.n13282 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_adj_1370_LC_22_22_6 .C_ON=1'b0;
    defparam \c0.i3_3_lut_adj_1370_LC_22_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_adj_1370_LC_22_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_3_lut_adj_1370_LC_22_22_6  (
            .in0(N__56322),
            .in1(N__56304),
            .in2(_gnd_net_),
            .in3(N__56293),
            .lcout(),
            .ltout(\c0.n8_adj_4291_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20116_4_lut_LC_22_22_7 .C_ON=1'b0;
    defparam \c0.i20116_4_lut_LC_22_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i20116_4_lut_LC_22_22_7 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \c0.i20116_4_lut_LC_22_22_7  (
            .in0(N__56278),
            .in1(N__56248),
            .in2(N__56242),
            .in3(N__56239),
            .lcout(\c0.n23811 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i7_LC_22_23_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i7_LC_22_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i7_LC_22_23_1 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \c0.rx.r_Rx_Byte_i7_LC_22_23_1  (
            .in0(N__68784),
            .in1(N__59958),
            .in2(N__56220),
            .in3(N__59699),
            .lcout(rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66853),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i12_3_lut_LC_22_23_3 .C_ON=1'b0;
    defparam \c0.rx.i12_3_lut_LC_22_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i12_3_lut_LC_22_23_3 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \c0.rx.i12_3_lut_LC_22_23_3  (
            .in0(N__56810),
            .in1(N__59698),
            .in2(_gnd_net_),
            .in3(N__56186),
            .lcout(\c0.rx.n36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_4_lut_4_lut_LC_22_23_4 .C_ON=1'b0;
    defparam \c0.rx.i2_4_lut_4_lut_LC_22_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_4_lut_4_lut_LC_22_23_4 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \c0.rx.i2_4_lut_4_lut_LC_22_23_4  (
            .in0(N__56992),
            .in1(N__56809),
            .in2(N__56928),
            .in3(N__57058),
            .lcout(n14436),
            .ltout(n14436_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i11380_3_lut_4_lut_LC_22_23_5 .C_ON=1'b0;
    defparam \c0.rx.i11380_3_lut_4_lut_LC_22_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i11380_3_lut_4_lut_LC_22_23_5 .LUT_INIT=16'b1011000000110000;
    LogicCell40 \c0.rx.i11380_3_lut_4_lut_LC_22_23_5  (
            .in0(N__59747),
            .in1(N__56914),
            .in2(N__56164),
            .in3(N__59957),
            .lcout(n14917),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_adj_1174_LC_22_23_7 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_adj_1174_LC_22_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_adj_1174_LC_22_23_7 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \c0.rx.i2_3_lut_adj_1174_LC_22_23_7  (
            .in0(N__57091),
            .in1(N__59863),
            .in2(_gnd_net_),
            .in3(N__56161),
            .lcout(n12970),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i2_LC_22_24_0 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i2_LC_22_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i2_LC_22_24_0 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \c0.rx.r_Bit_Index_i2_LC_22_24_0  (
            .in0(N__59898),
            .in1(N__57115),
            .in2(N__57101),
            .in3(N__59911),
            .lcout(r_Bit_Index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66861),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i0_LC_22_24_1 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i0_LC_22_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i0_LC_22_24_1 .LUT_INIT=16'b0101000010101010;
    LogicCell40 \c0.rx.r_Bit_Index_i0_LC_22_24_1  (
            .in0(N__59752),
            .in1(_gnd_net_),
            .in2(N__56946),
            .in3(N__59897),
            .lcout(r_Bit_Index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66861),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15930_2_lut_LC_22_24_3 .C_ON=1'b0;
    defparam \c0.rx.i15930_2_lut_LC_22_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15930_2_lut_LC_22_24_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \c0.rx.i15930_2_lut_LC_22_24_3  (
            .in0(N__59751),
            .in1(_gnd_net_),
            .in2(N__59868),
            .in3(_gnd_net_),
            .lcout(n19619),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_LC_22_24_4 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_LC_22_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_LC_22_24_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i1_2_lut_LC_22_24_4  (
            .in0(_gnd_net_),
            .in1(N__59859),
            .in2(_gnd_net_),
            .in3(N__57090),
            .lcout(n91),
            .ltout(n91_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i28_3_lut_4_lut_LC_22_24_5 .C_ON=1'b0;
    defparam \c0.rx.i28_3_lut_4_lut_LC_22_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i28_3_lut_4_lut_LC_22_24_5 .LUT_INIT=16'b0010000011001100;
    LogicCell40 \c0.rx.i28_3_lut_4_lut_LC_22_24_5  (
            .in0(N__59750),
            .in1(N__56822),
            .in2(N__57064),
            .in3(N__57060),
            .lcout(),
            .ltout(\c0.rx.n14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i0_LC_22_24_6 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i0_LC_22_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i0_LC_22_24_6 .LUT_INIT=16'b0100000001010001;
    LogicCell40 \c0.rx.r_SM_Main_i0_LC_22_24_6  (
            .in0(N__57002),
            .in1(N__56939),
            .in2(N__56845),
            .in3(N__56842),
            .lcout(r_SM_Main_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66861),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_69_i9_2_lut_3_lut_LC_23_8_6 .C_ON=1'b0;
    defparam \c0.equal_69_i9_2_lut_3_lut_LC_23_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.equal_69_i9_2_lut_3_lut_LC_23_8_6 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \c0.equal_69_i9_2_lut_3_lut_LC_23_8_6  (
            .in0(N__56718),
            .in1(N__56598),
            .in2(_gnd_net_),
            .in3(N__56457),
            .lcout(\c0.n9_adj_4217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1260_LC_23_9_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1260_LC_23_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1260_LC_23_9_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1260_LC_23_9_0  (
            .in0(N__57126),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60234),
            .lcout(\c0.n22328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1664_LC_23_9_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1664_LC_23_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1664_LC_23_9_1 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1664_LC_23_9_1  (
            .in0(N__56692),
            .in1(N__56597),
            .in2(N__56458),
            .in3(N__62351),
            .lcout(n21755),
            .ltout(n21755_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i114_LC_23_9_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i114_LC_23_9_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i114_LC_23_9_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \c0.data_in_frame_0__i114_LC_23_9_2  (
            .in0(_gnd_net_),
            .in1(N__63831),
            .in2(N__56770),
            .in3(N__56763),
            .lcout(data_in_frame_14_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66694),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_68_i9_2_lut_3_lut_LC_23_9_3 .C_ON=1'b0;
    defparam \c0.equal_68_i9_2_lut_3_lut_LC_23_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.equal_68_i9_2_lut_3_lut_LC_23_9_3 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \c0.equal_68_i9_2_lut_3_lut_LC_23_9_3  (
            .in0(N__56691),
            .in1(N__56596),
            .in2(_gnd_net_),
            .in3(N__56439),
            .lcout(\c0.n9_adj_4237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1265_LC_23_9_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1265_LC_23_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1265_LC_23_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1265_LC_23_9_4  (
            .in0(_gnd_net_),
            .in1(N__57382),
            .in2(_gnd_net_),
            .in3(N__57365),
            .lcout(\c0.n22471 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1382_LC_23_9_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1382_LC_23_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1382_LC_23_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1382_LC_23_9_6  (
            .in0(N__57314),
            .in1(N__58205),
            .in2(_gnd_net_),
            .in3(N__57283),
            .lcout(\c0.n21069 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1266_LC_23_10_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1266_LC_23_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1266_LC_23_10_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1266_LC_23_10_0  (
            .in0(N__60255),
            .in1(N__57940),
            .in2(N__57187),
            .in3(N__57910),
            .lcout(\c0.n22446 ),
            .ltout(\c0.n22446_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1244_LC_23_10_1 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1244_LC_23_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1244_LC_23_10_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1244_LC_23_10_1  (
            .in0(N__58497),
            .in1(N__57234),
            .in2(N__57220),
            .in3(N__57216),
            .lcout(\c0.n30_adj_4233 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i115_LC_23_10_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i115_LC_23_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i115_LC_23_10_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i115_LC_23_10_2  (
            .in0(N__57186),
            .in1(N__57155),
            .in2(_gnd_net_),
            .in3(N__68443),
            .lcout(data_in_frame_14_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66707),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1304_LC_23_10_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1304_LC_23_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1304_LC_23_10_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1304_LC_23_10_3  (
            .in0(_gnd_net_),
            .in1(N__60233),
            .in2(_gnd_net_),
            .in3(N__60254),
            .lcout(\c0.n22340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i113_LC_23_10_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i113_LC_23_10_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i113_LC_23_10_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i113_LC_23_10_4  (
            .in0(N__57924),
            .in1(N__57154),
            .in2(_gnd_net_),
            .in3(N__69493),
            .lcout(data_in_frame_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66707),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i117_LC_23_10_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i117_LC_23_10_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i117_LC_23_10_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i117_LC_23_10_5  (
            .in0(N__57156),
            .in1(N__63176),
            .in2(_gnd_net_),
            .in3(N__57127),
            .lcout(data_in_frame_14_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66707),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i192_LC_23_10_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i192_LC_23_10_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i192_LC_23_10_6 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i192_LC_23_10_6  (
            .in0(N__68155),
            .in1(N__68591),
            .in2(N__65297),
            .in3(N__68979),
            .lcout(\c0.data_in_frame_23_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66707),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i146_LC_23_10_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i146_LC_23_10_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i146_LC_23_10_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i146_LC_23_10_7  (
            .in0(N__69203),
            .in1(N__68156),
            .in2(N__57469),
            .in3(N__63859),
            .lcout(\c0.data_in_frame_18_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66707),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_LC_23_11_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_LC_23_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_LC_23_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_LC_23_11_1  (
            .in0(N__57447),
            .in1(N__57869),
            .in2(_gnd_net_),
            .in3(N__61284),
            .lcout(\c0.n10_adj_4239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1327_LC_23_11_2 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1327_LC_23_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1327_LC_23_11_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_1327_LC_23_11_2  (
            .in0(N__60907),
            .in1(N__57498),
            .in2(N__61290),
            .in3(N__57523),
            .lcout(\c0.n22464 ),
            .ltout(\c0.n22464_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_1785_LC_23_11_3 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_1785_LC_23_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_1785_LC_23_11_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_1785_LC_23_11_3  (
            .in0(N__60383),
            .in1(N__60172),
            .in2(N__57514),
            .in3(N__57511),
            .lcout(\c0.n8_adj_4275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1788_LC_23_11_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1788_LC_23_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1788_LC_23_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1788_LC_23_11_4  (
            .in0(N__58067),
            .in1(N__60232),
            .in2(_gnd_net_),
            .in3(N__60253),
            .lcout(\c0.n10_adj_4267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1250_LC_23_11_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1250_LC_23_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1250_LC_23_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1250_LC_23_11_5  (
            .in0(N__57499),
            .in1(N__61329),
            .in2(N__58036),
            .in3(N__58068),
            .lcout(\c0.n14053 ),
            .ltout(\c0.n14053_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1347_LC_23_11_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1347_LC_23_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1347_LC_23_11_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_1347_LC_23_11_6  (
            .in0(N__57468),
            .in1(N__61242),
            .in2(N__57451),
            .in3(N__60531),
            .lcout(),
            .ltout(\c0.n23586_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1297_LC_23_11_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1297_LC_23_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1297_LC_23_11_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1297_LC_23_11_7  (
            .in0(N__62677),
            .in1(N__57448),
            .in2(N__57406),
            .in3(N__61285),
            .lcout(\c0.n23426 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1288_LC_23_12_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1288_LC_23_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1288_LC_23_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1288_LC_23_12_0  (
            .in0(N__61003),
            .in1(N__60002),
            .in2(_gnd_net_),
            .in3(N__57403),
            .lcout(\c0.n13210 ),
            .ltout(\c0.n13210_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1342_LC_23_12_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1342_LC_23_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1342_LC_23_12_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1342_LC_23_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__57736),
            .in3(N__57733),
            .lcout(),
            .ltout(\c0.n7_adj_4277_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1343_LC_23_12_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1343_LC_23_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1343_LC_23_12_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1343_LC_23_12_2  (
            .in0(N__60121),
            .in1(N__57691),
            .in2(N__57682),
            .in3(N__60406),
            .lcout(\c0.n21867 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i93_LC_23_12_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i93_LC_23_12_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i93_LC_23_12_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i93_LC_23_12_3  (
            .in0(N__67476),
            .in1(N__63124),
            .in2(N__61045),
            .in3(N__62531),
            .lcout(\c0.data_in_frame_11_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66735),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1789_LC_23_12_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1789_LC_23_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1789_LC_23_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1789_LC_23_12_4  (
            .in0(N__60139),
            .in1(N__57605),
            .in2(_gnd_net_),
            .in3(N__60511),
            .lcout(),
            .ltout(\c0.n10_adj_4264_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1322_LC_23_12_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1322_LC_23_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1322_LC_23_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1322_LC_23_12_5  (
            .in0(N__61040),
            .in1(N__57675),
            .in2(N__57658),
            .in3(N__57632),
            .lcout(\c0.n16_adj_4265 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i95_LC_23_12_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i95_LC_23_12_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i95_LC_23_12_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i95_LC_23_12_6  (
            .in0(N__62529),
            .in1(N__65569),
            .in2(N__57639),
            .in3(N__67451),
            .lcout(\c0.data_in_frame_11_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66735),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i91_LC_23_12_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i91_LC_23_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i91_LC_23_12_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i91_LC_23_12_7  (
            .in0(N__67475),
            .in1(N__68437),
            .in2(N__57614),
            .in3(N__62530),
            .lcout(\c0.data_in_frame_11_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66735),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1344_LC_23_13_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1344_LC_23_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1344_LC_23_13_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1344_LC_23_13_0  (
            .in0(_gnd_net_),
            .in1(N__61517),
            .in2(_gnd_net_),
            .in3(N__58098),
            .lcout(\c0.n21845 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1565_LC_23_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1565_LC_23_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1565_LC_23_13_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1565_LC_23_13_1  (
            .in0(N__57850),
            .in1(N__57592),
            .in2(N__57553),
            .in3(N__57541),
            .lcout(\c0.n6_adj_4225 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_LC_23_13_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_LC_23_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_LC_23_13_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_3_lut_LC_23_13_3  (
            .in0(N__57936),
            .in1(N__57925),
            .in2(_gnd_net_),
            .in3(N__57908),
            .lcout(\c0.n22352 ),
            .ltout(\c0.n22352_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1253_LC_23_13_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1253_LC_23_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1253_LC_23_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1253_LC_23_13_4  (
            .in0(N__57874),
            .in1(N__57849),
            .in2(N__57829),
            .in3(N__61235),
            .lcout(\c0.n22000 ),
            .ltout(\c0.n22000_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1245_LC_23_13_5 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1245_LC_23_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1245_LC_23_13_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1245_LC_23_13_5  (
            .in0(N__57809),
            .in1(N__61172),
            .in2(N__57826),
            .in3(N__60546),
            .lcout(\c0.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i128_LC_23_13_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i128_LC_23_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i128_LC_23_13_6 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \c0.data_in_frame_0__i128_LC_23_13_6  (
            .in0(N__62541),
            .in1(N__57810),
            .in2(N__68680),
            .in3(N__68908),
            .lcout(\c0.data_in_frame_15_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66749),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i100_LC_23_14_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i100_LC_23_14_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i100_LC_23_14_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i100_LC_23_14_1  (
            .in0(N__62557),
            .in1(N__64481),
            .in2(N__61500),
            .in3(N__64874),
            .lcout(\c0.data_in_frame_12_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66764),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_LC_23_14_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_LC_23_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_LC_23_14_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_LC_23_14_3  (
            .in0(N__61254),
            .in1(N__61518),
            .in2(N__57795),
            .in3(N__61884),
            .lcout(),
            .ltout(\c0.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1254_LC_23_14_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1254_LC_23_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1254_LC_23_14_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1254_LC_23_14_4  (
            .in0(N__64173),
            .in1(N__57778),
            .in2(N__57769),
            .in3(N__58062),
            .lcout(\c0.n20246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1251_LC_23_14_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1251_LC_23_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1251_LC_23_14_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1251_LC_23_14_5  (
            .in0(N__58061),
            .in1(N__57766),
            .in2(N__57757),
            .in3(N__57742),
            .lcout(\c0.n13544 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1237_LC_23_14_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1237_LC_23_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1237_LC_23_14_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1237_LC_23_14_6  (
            .in0(N__58243),
            .in1(N__61149),
            .in2(N__58237),
            .in3(N__58212),
            .lcout(\c0.n10_adj_4230 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_3_lut_4_lut_LC_23_15_1 .C_ON=1'b0;
    defparam \c0.i5_2_lut_3_lut_4_lut_LC_23_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_3_lut_4_lut_LC_23_15_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_2_lut_3_lut_4_lut_LC_23_15_1  (
            .in0(N__58018),
            .in1(N__58185),
            .in2(N__58173),
            .in3(N__58063),
            .lcout(\c0.n18_adj_4246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_LC_23_15_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_LC_23_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_LC_23_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_LC_23_15_2  (
            .in0(N__58141),
            .in1(N__58094),
            .in2(_gnd_net_),
            .in3(N__58075),
            .lcout(\c0.n22849 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i201_LC_23_15_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i201_LC_23_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i201_LC_23_15_3 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i201_LC_23_15_3  (
            .in0(N__69565),
            .in1(N__58637),
            .in2(N__69878),
            .in3(N__67757),
            .lcout(\c0.data_in_frame_25_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66776),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i109_LC_23_15_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i109_LC_23_15_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i109_LC_23_15_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i109_LC_23_15_4  (
            .in0(N__63139),
            .in1(N__62058),
            .in2(N__58069),
            .in3(N__62507),
            .lcout(\c0.data_in_frame_13_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66776),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i126_LC_23_15_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i126_LC_23_15_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i126_LC_23_15_6 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i126_LC_23_15_6  (
            .in0(N__68678),
            .in1(N__62506),
            .in2(N__58028),
            .in3(N__67070),
            .lcout(\c0.data_in_frame_15_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66776),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1190_LC_23_16_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1190_LC_23_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1190_LC_23_16_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1190_LC_23_16_1  (
            .in0(N__62787),
            .in1(N__65146),
            .in2(N__57997),
            .in3(N__57973),
            .lcout(\c0.n22402 ),
            .ltout(\c0.n22402_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_4_lut_LC_23_16_2 .C_ON=1'b0;
    defparam \c0.i4_3_lut_4_lut_LC_23_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_4_lut_LC_23_16_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_3_lut_4_lut_LC_23_16_2  (
            .in0(N__59488),
            .in1(N__65061),
            .in2(N__57955),
            .in3(N__65179),
            .lcout(\c0.n33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i213_LC_23_16_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i213_LC_23_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i213_LC_23_16_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i213_LC_23_16_3  (
            .in0(N__63225),
            .in1(N__69204),
            .in2(N__59499),
            .in3(N__67759),
            .lcout(\c0.data_in_frame_26_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66789),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1372_LC_23_16_4 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1372_LC_23_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1372_LC_23_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_3_lut_adj_1372_LC_23_16_4  (
            .in0(N__59489),
            .in1(N__64947),
            .in2(_gnd_net_),
            .in3(N__58390),
            .lcout(),
            .ltout(\c0.n6_adj_4292_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1379_LC_23_16_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1379_LC_23_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1379_LC_23_16_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1379_LC_23_16_5  (
            .in0(N__65062),
            .in1(N__58996),
            .in2(N__58384),
            .in3(N__58381),
            .lcout(\c0.n23073 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1277_LC_23_16_6 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1277_LC_23_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1277_LC_23_16_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1277_LC_23_16_6  (
            .in0(N__58342),
            .in1(N__58300),
            .in2(N__61209),
            .in3(N__62850),
            .lcout(\c0.n24_adj_4248 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1348_LC_23_17_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1348_LC_23_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1348_LC_23_17_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1348_LC_23_17_0  (
            .in0(_gnd_net_),
            .in1(N__62765),
            .in2(_gnd_net_),
            .in3(N__58256),
            .lcout(\c0.n21905 ),
            .ltout(\c0.n21905_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1349_LC_23_17_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1349_LC_23_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1349_LC_23_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1349_LC_23_17_1  (
            .in0(N__61667),
            .in1(N__62893),
            .in2(N__58294),
            .in3(N__64111),
            .lcout(\c0.n20288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1270_LC_23_17_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1270_LC_23_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1270_LC_23_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1270_LC_23_17_2  (
            .in0(N__65719),
            .in1(N__66049),
            .in2(_gnd_net_),
            .in3(N__58291),
            .lcout(\c0.n22399 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1739_LC_23_17_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1739_LC_23_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1739_LC_23_17_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_4_lut_adj_1739_LC_23_17_3  (
            .in0(N__58257),
            .in1(N__58279),
            .in2(N__59832),
            .in3(N__62702),
            .lcout(\c0.n22020 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i164_LC_23_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i164_LC_23_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i164_LC_23_17_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i164_LC_23_17_4  (
            .in0(N__64535),
            .in1(N__68086),
            .in2(N__58261),
            .in3(N__64853),
            .lcout(\c0.data_in_frame_20_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66799),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i196_LC_23_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i196_LC_23_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i196_LC_23_17_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i196_LC_23_17_5  (
            .in0(N__64852),
            .in1(N__66001),
            .in2(N__59006),
            .in3(N__67676),
            .lcout(\c0.data_in_frame_24_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66799),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1856_LC_23_17_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1856_LC_23_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1856_LC_23_17_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1856_LC_23_17_6  (
            .in0(N__61741),
            .in1(N__61666),
            .in2(N__62706),
            .in3(N__58541),
            .lcout(\c0.n22458 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i165_LC_23_17_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i165_LC_23_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i165_LC_23_17_7 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i165_LC_23_17_7  (
            .in0(N__62766),
            .in1(N__63178),
            .in2(N__68147),
            .in3(N__64536),
            .lcout(\c0.data_in_frame_20_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66799),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_4_lut_LC_23_18_0 .C_ON=1'b0;
    defparam \c0.i4_2_lut_4_lut_LC_23_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_4_lut_LC_23_18_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_2_lut_4_lut_LC_23_18_0  (
            .in0(N__59335),
            .in1(N__58446),
            .in2(N__63310),
            .in3(N__58458),
            .lcout(),
            .ltout(\c0.n18_adj_4249_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1279_LC_23_18_1 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1279_LC_23_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1279_LC_23_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1279_LC_23_18_1  (
            .in0(N__65364),
            .in1(N__58528),
            .in2(N__58516),
            .in3(N__58513),
            .lcout(\c0.n26_adj_4250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1272_LC_23_18_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1272_LC_23_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1272_LC_23_18_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1272_LC_23_18_2  (
            .in0(N__64054),
            .in1(N__58490),
            .in2(N__63416),
            .in3(N__61786),
            .lcout(\c0.n23072 ),
            .ltout(\c0.n23072_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1274_LC_23_18_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1274_LC_23_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1274_LC_23_18_3 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.i2_3_lut_adj_1274_LC_23_18_3  (
            .in0(N__58447),
            .in1(_gnd_net_),
            .in2(N__58432),
            .in3(N__63308),
            .lcout(\c0.n22364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1256_LC_23_18_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1256_LC_23_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1256_LC_23_18_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_1256_LC_23_18_4  (
            .in0(_gnd_net_),
            .in1(N__62707),
            .in2(_gnd_net_),
            .in3(N__61668),
            .lcout(\c0.n21124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1284_LC_23_18_5 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1284_LC_23_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1284_LC_23_18_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1284_LC_23_18_5  (
            .in0(N__58428),
            .in1(N__63316),
            .in2(N__65400),
            .in3(N__58396),
            .lcout(\c0.n21039 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i161_LC_23_18_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i161_LC_23_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i161_LC_23_18_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i161_LC_23_18_6  (
            .in0(N__59336),
            .in1(N__69560),
            .in2(N__68164),
            .in3(N__64560),
            .lcout(\c0.data_in_frame_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66808),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1356_LC_23_19_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1356_LC_23_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1356_LC_23_19_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i5_3_lut_adj_1356_LC_23_19_0  (
            .in0(N__58837),
            .in1(N__58774),
            .in2(_gnd_net_),
            .in3(N__58726),
            .lcout(\c0.n14_adj_4283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1352_LC_23_19_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1352_LC_23_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1352_LC_23_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1352_LC_23_19_1  (
            .in0(N__60490),
            .in1(N__61695),
            .in2(N__60277),
            .in3(N__58740),
            .lcout(),
            .ltout(\c0.n24_adj_4282_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1354_LC_23_19_2 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1354_LC_23_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1354_LC_23_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1354_LC_23_19_2  (
            .in0(N__59770),
            .in1(N__65206),
            .in2(N__58729),
            .in3(N__63238),
            .lcout(\c0.n22711 ),
            .ltout(\c0.n22711_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1209_LC_23_19_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1209_LC_23_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1209_LC_23_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1209_LC_23_19_3  (
            .in0(_gnd_net_),
            .in1(N__63560),
            .in2(N__58720),
            .in3(N__58712),
            .lcout(\c0.n21087 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1357_LC_23_19_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1357_LC_23_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1357_LC_23_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1357_LC_23_19_4  (
            .in0(N__63432),
            .in1(N__58696),
            .in2(N__58675),
            .in3(N__58651),
            .lcout(),
            .ltout(\c0.n15_adj_4284_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1359_LC_23_19_5 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1359_LC_23_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1359_LC_23_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1359_LC_23_19_5  (
            .in0(N__62599),
            .in1(N__63877),
            .in2(N__58660),
            .in3(N__58657),
            .lcout(\c0.n22373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1212_LC_23_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1212_LC_23_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1212_LC_23_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1212_LC_23_20_0  (
            .in0(_gnd_net_),
            .in1(N__69595),
            .in2(_gnd_net_),
            .in3(N__59031),
            .lcout(\c0.n22437 ),
            .ltout(\c0.n22437_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_adj_1730_LC_23_20_1 .C_ON=1'b0;
    defparam \c0.i21_4_lut_adj_1730_LC_23_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_adj_1730_LC_23_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i21_4_lut_adj_1730_LC_23_20_1  (
            .in0(N__58643),
            .in1(N__58618),
            .in2(N__58573),
            .in3(N__59044),
            .lcout(\c0.n50_adj_4487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1904_LC_23_20_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1904_LC_23_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1904_LC_23_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1904_LC_23_20_2  (
            .in0(N__63501),
            .in1(N__58560),
            .in2(N__63546),
            .in3(N__59065),
            .lcout(\c0.n20537 ),
            .ltout(\c0.n20537_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1723_LC_23_20_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1723_LC_23_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1723_LC_23_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1723_LC_23_20_3  (
            .in0(N__59104),
            .in1(N__59256),
            .in2(N__59095),
            .in3(N__59092),
            .lcout(\c0.n21890 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1563_LC_23_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1563_LC_23_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1563_LC_23_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1563_LC_23_20_4  (
            .in0(N__58953),
            .in1(N__65193),
            .in2(N__65053),
            .in3(N__59008),
            .lcout(\c0.n13320 ),
            .ltout(\c0.n13320_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_LC_23_20_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_LC_23_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_LC_23_20_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_LC_23_20_5  (
            .in0(N__59066),
            .in1(N__68712),
            .in2(N__59047),
            .in3(N__59043),
            .lcout(),
            .ltout(\c0.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1897_LC_23_20_6 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1897_LC_23_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1897_LC_23_20_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1897_LC_23_20_6  (
            .in0(N__64258),
            .in1(N__64224),
            .in2(N__59035),
            .in3(N__59032),
            .lcout(\c0.n22314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1210_LC_23_20_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1210_LC_23_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1210_LC_23_20_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1210_LC_23_20_7  (
            .in0(_gnd_net_),
            .in1(N__59007),
            .in2(_gnd_net_),
            .in3(N__58952),
            .lcout(\c0.n22142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1206_LC_23_21_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1206_LC_23_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1206_LC_23_21_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1206_LC_23_21_0  (
            .in0(N__58960),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59257),
            .lcout(\c0.n22337 ),
            .ltout(\c0.n22337_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1743_LC_23_21_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1743_LC_23_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1743_LC_23_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1743_LC_23_21_1  (
            .in0(N__58852),
            .in1(N__58918),
            .in2(N__58906),
            .in3(N__58903),
            .lcout(\c0.n21095 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1651_LC_23_21_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1651_LC_23_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1651_LC_23_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1651_LC_23_21_2  (
            .in0(N__59446),
            .in1(N__66066),
            .in2(N__68705),
            .in3(N__59409),
            .lcout(\c0.n6_adj_4418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1361_LC_23_21_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1361_LC_23_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1361_LC_23_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1361_LC_23_21_3  (
            .in0(N__59500),
            .in1(N__64911),
            .in2(N__64275),
            .in3(N__59470),
            .lcout(),
            .ltout(\c0.n10_adj_4285_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1373_LC_23_21_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1373_LC_23_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1373_LC_23_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_1373_LC_23_21_4  (
            .in0(_gnd_net_),
            .in1(N__62635),
            .in2(N__59464),
            .in3(N__65016),
            .lcout(\c0.n22995 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1741_LC_23_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1741_LC_23_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1741_LC_23_21_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1741_LC_23_21_5  (
            .in0(_gnd_net_),
            .in1(N__59445),
            .in2(_gnd_net_),
            .in3(N__68695),
            .lcout(\c0.n22054 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1740_LC_23_21_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1740_LC_23_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1740_LC_23_21_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1740_LC_23_21_6  (
            .in0(_gnd_net_),
            .in1(N__66067),
            .in2(_gnd_net_),
            .in3(N__59410),
            .lcout(\c0.n22434 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1203_LC_23_21_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1203_LC_23_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1203_LC_23_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1203_LC_23_21_7  (
            .in0(N__59352),
            .in1(N__61641),
            .in2(N__59317),
            .in3(N__59290),
            .lcout(\c0.n20596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i96_LC_23_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i96_LC_23_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i96_LC_23_22_2 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i96_LC_23_22_2  (
            .in0(N__68785),
            .in1(N__62508),
            .in2(N__67480),
            .in3(N__59226),
            .lcout(\c0.data_in_frame_11_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66854),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i180_LC_23_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i180_LC_23_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i180_LC_23_22_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i180_LC_23_22_3  (
            .in0(N__64885),
            .in1(N__61694),
            .in2(_gnd_net_),
            .in3(N__59212),
            .lcout(data_in_frame_22_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66854),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i174_LC_23_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i174_LC_23_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i174_LC_23_22_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i174_LC_23_22_4  (
            .in0(N__65357),
            .in1(N__66974),
            .in2(N__62121),
            .in3(N__68160),
            .lcout(\c0.data_in_frame_21_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66854),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_LC_23_22_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_LC_23_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_LC_23_22_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_LC_23_22_5  (
            .in0(N__63573),
            .in1(N__65356),
            .in2(N__59125),
            .in3(N__59976),
            .lcout(\c0.n22215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i156_LC_23_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i156_LC_23_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i156_LC_23_22_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i156_LC_23_22_6  (
            .in0(N__67471),
            .in1(N__68159),
            .in2(N__63917),
            .in3(N__64886),
            .lcout(\c0.data_in_frame_19_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66854),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i6_LC_23_22_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i6_LC_23_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i6_LC_23_22_7 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.rx.r_Rx_Byte_i6_LC_23_22_7  (
            .in0(N__65501),
            .in1(N__59965),
            .in2(N__59709),
            .in3(N__59939),
            .lcout(rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66854),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i4_LC_23_23_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i4_LC_23_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i4_LC_23_23_1 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.rx.r_Rx_Byte_i4_LC_23_23_1  (
            .in0(N__62975),
            .in1(N__59756),
            .in2(N__59715),
            .in3(N__59592),
            .lcout(rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66862),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i1_LC_23_23_2 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i1_LC_23_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i1_LC_23_23_2 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \c0.rx.r_Bit_Index_i1_LC_23_23_2  (
            .in0(N__59910),
            .in1(N__59864),
            .in2(N__59758),
            .in3(N__59899),
            .lcout(r_Bit_Index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66862),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1353_LC_23_23_4 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1353_LC_23_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1353_LC_23_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1353_LC_23_23_4  (
            .in0(N__67811),
            .in1(N__59833),
            .in2(N__62752),
            .in3(N__59787),
            .lcout(\c0.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i5_LC_23_23_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i5_LC_23_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i5_LC_23_23_6 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \c0.rx.r_Rx_Byte_i5_LC_23_23_6  (
            .in0(N__59757),
            .in1(N__59708),
            .in2(N__59593),
            .in3(N__66975),
            .lcout(rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66862),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i97_LC_24_9_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i97_LC_24_9_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i97_LC_24_9_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i97_LC_24_9_7  (
            .in0(N__64345),
            .in1(N__62378),
            .in2(N__59578),
            .in3(N__69502),
            .lcout(\c0.data_in_frame_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66708),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i200_LC_24_10_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i200_LC_24_10_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i200_LC_24_10_1 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i200_LC_24_10_1  (
            .in0(N__68980),
            .in1(N__66030),
            .in2(N__59522),
            .in3(N__67775),
            .lcout(\c0.data_in_frame_24_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66722),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i98_LC_24_10_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i98_LC_24_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i98_LC_24_10_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i98_LC_24_10_2  (
            .in0(N__64356),
            .in1(N__62525),
            .in2(N__60259),
            .in3(N__63861),
            .lcout(\c0.data_in_frame_12_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66722),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i99_LC_24_10_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i99_LC_24_10_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i99_LC_24_10_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i99_LC_24_10_3  (
            .in0(N__62522),
            .in1(N__64357),
            .in2(N__68442),
            .in3(N__60235),
            .lcout(\c0.data_in_frame_12_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66722),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i107_LC_24_10_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i107_LC_24_10_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i107_LC_24_10_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i107_LC_24_10_4  (
            .in0(N__61970),
            .in1(N__62524),
            .in2(N__60211),
            .in3(N__68433),
            .lcout(\c0.data_in_frame_13_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66722),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1786_LC_24_10_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1786_LC_24_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1786_LC_24_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1786_LC_24_10_5  (
            .in0(N__60207),
            .in1(N__61138),
            .in2(_gnd_net_),
            .in3(N__61107),
            .lcout(\c0.n22274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i106_LC_24_10_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i106_LC_24_10_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i106_LC_24_10_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i106_LC_24_10_6  (
            .in0(N__61969),
            .in1(N__62523),
            .in2(N__60195),
            .in3(N__63860),
            .lcout(\c0.data_in_frame_13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66722),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i89_LC_24_11_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i89_LC_24_11_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i89_LC_24_11_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i89_LC_24_11_1  (
            .in0(N__67408),
            .in1(N__69492),
            .in2(N__60150),
            .in3(N__62527),
            .lcout(\c0.data_in_frame_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66736),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1305_LC_24_11_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1305_LC_24_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1305_LC_24_11_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1305_LC_24_11_2  (
            .in0(_gnd_net_),
            .in1(N__60143),
            .in2(_gnd_net_),
            .in3(N__60512),
            .lcout(),
            .ltout(\c0.n13999_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1248_LC_24_11_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1248_LC_24_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1248_LC_24_11_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1248_LC_24_11_3  (
            .in0(N__60117),
            .in1(N__60102),
            .in2(N__60061),
            .in3(N__60058),
            .lcout(\c0.n13233 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i75_LC_24_11_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i75_LC_24_11_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i75_LC_24_11_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i75_LC_24_11_4  (
            .in0(N__62526),
            .in1(N__69880),
            .in2(N__68441),
            .in3(N__60003),
            .lcout(\c0.data_in_frame_9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66736),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1346_LC_24_11_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1346_LC_24_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1346_LC_24_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1346_LC_24_11_5  (
            .in0(N__60553),
            .in1(N__61542),
            .in2(N__61261),
            .in3(N__60535),
            .lcout(\c0.n21114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3286_2_lut_LC_24_11_6 .C_ON=1'b0;
    defparam \c0.i3286_2_lut_LC_24_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3286_2_lut_LC_24_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3286_2_lut_LC_24_11_6  (
            .in0(_gnd_net_),
            .in1(N__62671),
            .in2(_gnd_net_),
            .in3(N__61886),
            .lcout(\c0.n5965 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i90_LC_24_11_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i90_LC_24_11_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i90_LC_24_11_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i90_LC_24_11_7  (
            .in0(N__63793),
            .in1(N__67457),
            .in2(N__60519),
            .in3(N__62528),
            .lcout(\c0.data_in_frame_11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66736),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i188_LC_24_12_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i188_LC_24_12_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i188_LC_24_12_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i188_LC_24_12_1  (
            .in0(N__68157),
            .in1(N__68552),
            .in2(N__60482),
            .in3(N__64873),
            .lcout(\c0.data_in_frame_23_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66750),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i186_LC_24_12_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i186_LC_24_12_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i186_LC_24_12_2 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \c0.data_in_frame_0__i186_LC_24_12_2  (
            .in0(N__60333),
            .in1(N__63830),
            .in2(N__68590),
            .in3(N__68158),
            .lcout(\c0.data_in_frame_23_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66750),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1341_LC_24_12_3 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1341_LC_24_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1341_LC_24_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_1341_LC_24_12_3  (
            .in0(N__60451),
            .in1(N__60436),
            .in2(N__60421),
            .in3(N__60412),
            .lcout(\c0.n8_adj_4276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i105_LC_24_12_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i105_LC_24_12_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i105_LC_24_12_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i105_LC_24_12_4  (
            .in0(N__62544),
            .in1(N__62120),
            .in2(N__60398),
            .in3(N__69564),
            .lcout(\c0.data_in_frame_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66750),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i104_LC_24_12_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i104_LC_24_12_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i104_LC_24_12_5 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i104_LC_24_12_5  (
            .in0(N__68866),
            .in1(N__62545),
            .in2(N__64458),
            .in3(N__60356),
            .lcout(\c0.data_in_frame_12_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66750),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1281_LC_24_12_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1281_LC_24_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1281_LC_24_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1281_LC_24_12_6  (
            .in0(_gnd_net_),
            .in1(N__60329),
            .in2(_gnd_net_),
            .in3(N__60311),
            .lcout(\c0.n21995 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i59_LC_24_12_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i59_LC_24_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i59_LC_24_12_7 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i59_LC_24_12_7  (
            .in0(N__60863),
            .in1(N__68553),
            .in2(N__60997),
            .in3(N__68434),
            .lcout(\c0.data_in_frame_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66750),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i176_LC_24_13_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i176_LC_24_13_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i176_LC_24_13_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i176_LC_24_13_0  (
            .in0(N__62086),
            .in1(N__68148),
            .in2(N__61202),
            .in3(N__68909),
            .lcout(\c0.data_in_frame_21_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66765),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1859_LC_24_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1859_LC_24_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1859_LC_24_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1859_LC_24_13_1  (
            .in0(N__61887),
            .in1(N__62672),
            .in2(_gnd_net_),
            .in3(N__61176),
            .lcout(\c0.n22091 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1578_LC_24_13_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1578_LC_24_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1578_LC_24_13_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1578_LC_24_13_3  (
            .in0(_gnd_net_),
            .in1(N__61131),
            .in2(_gnd_net_),
            .in3(N__61111),
            .lcout(\c0.n13421 ),
            .ltout(\c0.n13421_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1287_LC_24_13_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1287_LC_24_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1287_LC_24_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1287_LC_24_13_4  (
            .in0(N__61044),
            .in1(N__60972),
            .in2(N__61027),
            .in3(N__61023),
            .lcout(\c0.n10_adj_4252 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1303_LC_24_13_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1303_LC_24_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1303_LC_24_13_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1303_LC_24_13_5  (
            .in0(N__60989),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60566),
            .lcout(\c0.n22343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1325_LC_24_13_6 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1325_LC_24_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1325_LC_24_13_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1325_LC_24_13_6  (
            .in0(N__61312),
            .in1(N__60958),
            .in2(N__60949),
            .in3(N__61448),
            .lcout(\c0.n16_adj_4268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i57_LC_24_13_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i57_LC_24_13_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i57_LC_24_13_7 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \c0.data_in_frame_0__i57_LC_24_13_7  (
            .in0(N__68545),
            .in1(N__60567),
            .in2(N__60893),
            .in3(N__69450),
            .lcout(\c0.data_in_frame_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66765),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i166_LC_24_14_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i166_LC_24_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i166_LC_24_14_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i166_LC_24_14_0  (
            .in0(N__68143),
            .in1(N__64534),
            .in2(N__63309),
            .in3(N__67104),
            .lcout(\c0.data_in_frame_20_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i130_LC_24_14_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i130_LC_24_14_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i130_LC_24_14_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i130_LC_24_14_1  (
            .in0(N__65992),
            .in1(N__68144),
            .in2(N__61525),
            .in3(N__63851),
            .lcout(\c0.data_in_frame_16_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i160_LC_24_14_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i160_LC_24_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i160_LC_24_14_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i160_LC_24_14_2  (
            .in0(N__68142),
            .in1(N__67453),
            .in2(N__63355),
            .in3(N__68971),
            .lcout(\c0.data_in_frame_19_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1299_LC_24_14_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1299_LC_24_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1299_LC_24_14_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1299_LC_24_14_3  (
            .in0(_gnd_net_),
            .in1(N__61343),
            .in2(_gnd_net_),
            .in3(N__61481),
            .lcout(\c0.n21975 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_LC_24_14_4 .C_ON=1'b0;
    defparam \c0.i5_2_lut_LC_24_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_LC_24_14_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i5_2_lut_LC_24_14_4  (
            .in0(_gnd_net_),
            .in1(N__61434),
            .in2(_gnd_net_),
            .in3(N__61390),
            .lcout(\c0.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i101_LC_24_14_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i101_LC_24_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i101_LC_24_14_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i101_LC_24_14_5  (
            .in0(N__64533),
            .in1(N__62556),
            .in2(N__61359),
            .in3(N__63161),
            .lcout(\c0.data_in_frame_12_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i108_LC_24_14_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i108_LC_24_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i108_LC_24_14_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i108_LC_24_14_6  (
            .in0(N__62555),
            .in1(N__62087),
            .in2(N__61330),
            .in3(N__64875),
            .lcout(\c0.data_in_frame_13_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1345_LC_24_14_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1345_LC_24_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1345_LC_24_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1345_LC_24_14_7  (
            .in0(_gnd_net_),
            .in1(N__62661),
            .in2(_gnd_net_),
            .in3(N__61294),
            .lcout(\c0.n14081 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i129_LC_24_15_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i129_LC_24_15_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i129_LC_24_15_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i129_LC_24_15_1  (
            .in0(N__65940),
            .in1(N__68145),
            .in2(N__61243),
            .in3(N__69566),
            .lcout(\c0.data_in_frame_16_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66790),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1197_LC_24_15_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1197_LC_24_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1197_LC_24_15_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1197_LC_24_15_2  (
            .in0(N__63295),
            .in1(N__62770),
            .in2(N__62751),
            .in3(N__62698),
            .lcout(\c0.n22105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i111_LC_24_15_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i111_LC_24_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i111_LC_24_15_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i111_LC_24_15_3  (
            .in0(N__65570),
            .in1(N__62503),
            .in2(N__62676),
            .in3(N__62181),
            .lcout(\c0.data_in_frame_13_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66790),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i214_LC_24_15_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i214_LC_24_15_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i214_LC_24_15_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i214_LC_24_15_4  (
            .in0(N__69151),
            .in1(N__67103),
            .in2(N__62630),
            .in3(N__67744),
            .lcout(\c0.data_in_frame_26_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66790),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i175_LC_24_15_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i175_LC_24_15_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i175_LC_24_15_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i175_LC_24_15_5  (
            .in0(N__65571),
            .in1(N__68146),
            .in2(N__62591),
            .in3(N__62182),
            .lcout(\c0.data_in_frame_21_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66790),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i112_LC_24_15_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i112_LC_24_15_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i112_LC_24_15_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i112_LC_24_15_6  (
            .in0(N__62502),
            .in1(N__68970),
            .in2(N__62203),
            .in3(N__61885),
            .lcout(\c0.data_in_frame_13_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66790),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_4_lut_LC_24_16_3 .C_ON=1'b0;
    defparam \c0.i7_3_lut_4_lut_LC_24_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_4_lut_LC_24_16_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_3_lut_4_lut_LC_24_16_3  (
            .in0(N__61852),
            .in1(N__61828),
            .in2(N__62901),
            .in3(N__64207),
            .lcout(\c0.n20_adj_4247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_1896_LC_24_16_4 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_1896_LC_24_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_1896_LC_24_16_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_1896_LC_24_16_4  (
            .in0(N__61774),
            .in1(N__61746),
            .in2(N__61708),
            .in3(N__61672),
            .lcout(\c0.n22007 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1257_LC_24_16_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1257_LC_24_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1257_LC_24_16_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1257_LC_24_16_5  (
            .in0(_gnd_net_),
            .in1(N__63351),
            .in2(_gnd_net_),
            .in3(N__61618),
            .lcout(\c0.n13768 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1276_LC_24_16_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1276_LC_24_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1276_LC_24_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1276_LC_24_16_7  (
            .in0(N__61578),
            .in1(N__61561),
            .in2(_gnd_net_),
            .in3(N__61546),
            .lcout(\c0.n14143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i154_LC_24_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i154_LC_24_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i154_LC_24_17_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i154_LC_24_17_1  (
            .in0(N__67469),
            .in1(N__68087),
            .in2(N__63417),
            .in3(N__63813),
            .lcout(\c0.data_in_frame_19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66809),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i198_LC_24_17_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i198_LC_24_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i198_LC_24_17_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i198_LC_24_17_2  (
            .in0(N__67673),
            .in1(N__65949),
            .in2(N__63539),
            .in3(N__67063),
            .lcout(\c0.data_in_frame_24_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66809),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1283_LC_24_17_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1283_LC_24_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1283_LC_24_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1283_LC_24_17_3  (
            .in0(N__63387),
            .in1(N__63364),
            .in2(N__63358),
            .in3(N__64123),
            .lcout(\c0.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1351_LC_24_17_5 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1351_LC_24_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1351_LC_24_17_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i11_4_lut_adj_1351_LC_24_17_5  (
            .in0(N__63304),
            .in1(N__62869),
            .in2(N__62827),
            .in3(N__63267),
            .lcout(\c0.n26_adj_4281 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i229_LC_24_17_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i229_LC_24_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i229_LC_24_17_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i229_LC_24_17_7  (
            .in0(N__64498),
            .in1(N__63106),
            .in2(N__64932),
            .in3(N__67674),
            .lcout(\c0.data_in_frame_28_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66809),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1496_LC_24_18_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1496_LC_24_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1496_LC_24_18_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1496_LC_24_18_0  (
            .in0(N__62902),
            .in1(N__64110),
            .in2(_gnd_net_),
            .in3(N__64219),
            .lcout(\c0.n22095 ),
            .ltout(\c0.n22095_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_LC_24_18_1 .C_ON=1'b0;
    defparam \c0.i12_4_lut_LC_24_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_LC_24_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_LC_24_18_1  (
            .in0(N__62863),
            .in1(N__66048),
            .in2(N__62857),
            .in3(N__62854),
            .lcout(\c0.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1883_LC_24_18_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1883_LC_24_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1883_LC_24_18_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1883_LC_24_18_3  (
            .in0(_gnd_net_),
            .in1(N__62826),
            .in2(_gnd_net_),
            .in3(N__63876),
            .lcout(\c0.n22267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1198_LC_24_18_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1198_LC_24_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1198_LC_24_18_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_1198_LC_24_18_4  (
            .in0(_gnd_net_),
            .in1(N__64244),
            .in2(_gnd_net_),
            .in3(N__64220),
            .lcout(\c0.n20406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_LC_24_18_6 .C_ON=1'b0;
    defparam \c0.i8_4_lut_LC_24_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_LC_24_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_LC_24_18_6  (
            .in0(N__64177),
            .in1(N__64156),
            .in2(N__64135),
            .in3(N__64122),
            .lcout(),
            .ltout(\c0.n21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1271_LC_24_18_7 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1271_LC_24_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1271_LC_24_18_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i11_4_lut_adj_1271_LC_24_18_7  (
            .in0(N__64109),
            .in1(N__64084),
            .in2(N__64072),
            .in3(N__64065),
            .lcout(\c0.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1218_LC_24_19_1 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1218_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1218_LC_24_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1218_LC_24_19_1  (
            .in0(N__64048),
            .in1(N__64036),
            .in2(N__63994),
            .in3(N__63979),
            .lcout(\c0.n23287 ),
            .ltout(\c0.n23287_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1355_LC_24_19_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1355_LC_24_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1355_LC_24_19_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1355_LC_24_19_2  (
            .in0(N__65304),
            .in1(N__65365),
            .in2(N__63922),
            .in3(N__63919),
            .lcout(\c0.n21921 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i194_LC_24_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i194_LC_24_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i194_LC_24_19_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i194_LC_24_19_3  (
            .in0(N__67791),
            .in1(N__66003),
            .in2(N__65060),
            .in3(N__63852),
            .lcout(\c0.data_in_frame_24_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66833),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i193_LC_24_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i193_LC_24_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i193_LC_24_19_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i193_LC_24_19_4  (
            .in0(N__66002),
            .in1(N__69451),
            .in2(N__63574),
            .in3(N__67792),
            .lcout(\c0.data_in_frame_24_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66833),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1564_LC_24_19_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1564_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1564_LC_24_19_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1564_LC_24_19_6  (
            .in0(N__65246),
            .in1(N__63538),
            .in2(N__63505),
            .in3(N__63485),
            .lcout(\c0.n22255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_LC_24_19_7 .C_ON=1'b0;
    defparam \c0.i8_3_lut_LC_24_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_LC_24_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i8_3_lut_LC_24_19_7  (
            .in0(N__65305),
            .in1(N__65265),
            .in2(_gnd_net_),
            .in3(N__65245),
            .lcout(\c0.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1205_LC_24_20_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1205_LC_24_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1205_LC_24_20_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_4_lut_adj_1205_LC_24_20_0  (
            .in0(N__65200),
            .in1(N__65154),
            .in2(N__65113),
            .in3(N__65080),
            .lcout(\c0.n22455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_adj_1365_LC_24_20_1 .C_ON=1'b0;
    defparam \c0.i3_3_lut_adj_1365_LC_24_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_adj_1365_LC_24_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_3_lut_adj_1365_LC_24_20_1  (
            .in0(N__65059),
            .in1(N__65020),
            .in2(_gnd_net_),
            .in3(N__64989),
            .lcout(),
            .ltout(\c0.n8_adj_4288_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1368_LC_24_20_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1368_LC_24_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1368_LC_24_20_2 .LUT_INIT=16'b1111111110010110;
    LogicCell40 \c0.i6_4_lut_adj_1368_LC_24_20_2  (
            .in0(N__64599),
            .in1(N__64963),
            .in2(N__64975),
            .in3(N__64900),
            .lcout(\c0.n24_adj_4289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1366_LC_24_20_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1366_LC_24_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1366_LC_24_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1366_LC_24_20_3  (
            .in0(N__64962),
            .in1(N__64951),
            .in2(N__64933),
            .in3(N__64912),
            .lcout(\c0.n22997 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i228_LC_24_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i228_LC_24_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i228_LC_24_20_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i228_LC_24_20_5  (
            .in0(N__64511),
            .in1(N__64864),
            .in2(N__64603),
            .in3(N__67794),
            .lcout(\c0.data_in_frame_28_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66845),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i232_LC_24_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i232_LC_24_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i232_LC_24_20_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i232_LC_24_20_6  (
            .in0(N__67793),
            .in1(N__64513),
            .in2(N__64587),
            .in3(N__68883),
            .lcout(\c0.data_in_frame_28_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66845),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i231_LC_24_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i231_LC_24_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i231_LC_24_20_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i231_LC_24_20_7  (
            .in0(N__64512),
            .in1(N__65574),
            .in2(N__64276),
            .in3(N__67795),
            .lcout(\c0.data_in_frame_28_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66845),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i224_LC_24_21_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i224_LC_24_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i224_LC_24_21_0 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i224_LC_24_21_0  (
            .in0(N__66124),
            .in1(N__68882),
            .in2(N__67479),
            .in3(N__67750),
            .lcout(\c0.data_in_frame_27_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i223_LC_24_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i223_LC_24_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i223_LC_24_21_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i223_LC_24_21_1  (
            .in0(N__67748),
            .in1(N__67462),
            .in2(N__66095),
            .in3(N__65503),
            .lcout(\c0.data_in_frame_27_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i217_LC_24_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i217_LC_24_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i217_LC_24_21_2 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i217_LC_24_21_2  (
            .in0(N__69561),
            .in1(N__66065),
            .in2(N__67478),
            .in3(N__67749),
            .lcout(\c0.data_in_frame_27_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3589_2_lut_LC_24_21_3 .C_ON=1'b0;
    defparam \c0.i3589_2_lut_LC_24_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3589_2_lut_LC_24_21_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3589_2_lut_LC_24_21_3  (
            .in0(_gnd_net_),
            .in1(N__65417),
            .in2(_gnd_net_),
            .in3(N__65378),
            .lcout(\c0.n6268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i136_LC_24_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i136_LC_24_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i136_LC_24_21_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i136_LC_24_21_4  (
            .in0(N__66031),
            .in1(N__68137),
            .in2(N__65750),
            .in3(N__68881),
            .lcout(\c0.data_in_frame_16_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i153_LC_24_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i153_LC_24_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i153_LC_24_21_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i153_LC_24_21_5  (
            .in0(N__68136),
            .in1(N__67461),
            .in2(N__65718),
            .in3(N__69562),
            .lcout(\c0.data_in_frame_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i151_LC_24_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i151_LC_24_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i151_LC_24_21_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i151_LC_24_21_6  (
            .in0(N__65502),
            .in1(N__69199),
            .in2(N__65424),
            .in3(N__68138),
            .lcout(\c0.data_in_frame_18_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i152_LC_24_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i152_LC_24_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i152_LC_24_21_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i152_LC_24_21_7  (
            .in0(N__68135),
            .in1(N__65379),
            .in2(N__69232),
            .in3(N__68876),
            .lcout(\c0.data_in_frame_18_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1360_LC_24_22_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1360_LC_24_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1360_LC_24_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1360_LC_24_22_1  (
            .in0(N__69584),
            .in1(N__69269),
            .in2(_gnd_net_),
            .in3(N__65355),
            .lcout(\c0.n22123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i208_LC_24_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i208_LC_24_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i208_LC_24_22_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i208_LC_24_22_2  (
            .in0(N__69879),
            .in1(N__68938),
            .in2(N__69594),
            .in3(N__67777),
            .lcout(\c0.data_in_frame_25_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66863),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i209_LC_24_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i209_LC_24_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i209_LC_24_22_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i209_LC_24_22_3  (
            .in0(N__67763),
            .in1(N__69198),
            .in2(N__69279),
            .in3(N__69452),
            .lcout(\c0.data_in_frame_26_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66863),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i216_LC_24_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i216_LC_24_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i216_LC_24_22_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i216_LC_24_22_4  (
            .in0(N__69197),
            .in1(N__68939),
            .in2(N__68713),
            .in3(N__67778),
            .lcout(\c0.data_in_frame_26_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66863),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i187_LC_24_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i187_LC_24_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i187_LC_24_22_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.data_in_frame_0__i187_LC_24_22_6  (
            .in0(N__68589),
            .in1(N__68435),
            .in2(N__67819),
            .in3(N__68165),
            .lcout(\c0.data_in_frame_23_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66863),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i222_LC_24_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i222_LC_24_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i222_LC_24_22_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i222_LC_24_22_7  (
            .in0(N__67764),
            .in1(N__67470),
            .in2(N__66912),
            .in3(N__67005),
            .lcout(\c0.data_in_frame_27_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__66863),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
