-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Aug 26 2019 00:03:51

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    PIN_9 : in std_logic;
    PIN_8 : in std_logic;
    PIN_7 : in std_logic;
    PIN_6 : in std_logic;
    PIN_5 : in std_logic;
    PIN_4 : in std_logic;
    PIN_3 : inout std_logic;
    PIN_24 : in std_logic;
    PIN_23 : in std_logic;
    PIN_22 : in std_logic;
    PIN_21 : in std_logic;
    PIN_20 : in std_logic;
    PIN_2 : in std_logic;
    PIN_19 : in std_logic;
    PIN_18 : in std_logic;
    PIN_17 : in std_logic;
    PIN_16 : in std_logic;
    PIN_15 : in std_logic;
    PIN_14 : in std_logic;
    PIN_13 : in std_logic;
    PIN_12 : in std_logic;
    PIN_11 : in std_logic;
    PIN_10 : in std_logic;
    PIN_1 : inout std_logic;
    LED : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__23697\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17070\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14964\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14142\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13751\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal n26 : std_logic;
signal \bfn_1_22_0_\ : std_logic;
signal n25 : std_logic;
signal n3851 : std_logic;
signal n24 : std_logic;
signal n3852 : std_logic;
signal n23 : std_logic;
signal n3853 : std_logic;
signal n22 : std_logic;
signal n3854 : std_logic;
signal n21 : std_logic;
signal n3855 : std_logic;
signal n20 : std_logic;
signal n3856 : std_logic;
signal n19 : std_logic;
signal n3857 : std_logic;
signal n3858 : std_logic;
signal n18 : std_logic;
signal \bfn_1_23_0_\ : std_logic;
signal n17 : std_logic;
signal n3859 : std_logic;
signal n16 : std_logic;
signal n3860 : std_logic;
signal n15 : std_logic;
signal n3861 : std_logic;
signal n14 : std_logic;
signal n3862 : std_logic;
signal n13 : std_logic;
signal n3863 : std_logic;
signal n12 : std_logic;
signal n3864 : std_logic;
signal n11 : std_logic;
signal n3865 : std_logic;
signal n3866 : std_logic;
signal n10 : std_logic;
signal \bfn_1_24_0_\ : std_logic;
signal n9 : std_logic;
signal n3867 : std_logic;
signal n8 : std_logic;
signal n3868 : std_logic;
signal n7 : std_logic;
signal n3869 : std_logic;
signal n6 : std_logic;
signal n3870 : std_logic;
signal n3871 : std_logic;
signal n3872 : std_logic;
signal n3873 : std_logic;
signal n3874 : std_logic;
signal \bfn_1_25_0_\ : std_logic;
signal n3875 : std_logic;
signal \c0.n4849_cascade_\ : std_logic;
signal \c0.n4568\ : std_logic;
signal \c0.n4582\ : std_logic;
signal \c0.n4591_cascade_\ : std_logic;
signal \c0.n28_cascade_\ : std_logic;
signal \c0.n22\ : std_logic;
signal \c0.data_in_frame_6_6\ : std_logic;
signal \c0.n4592\ : std_logic;
signal \c0.n25_cascade_\ : std_logic;
signal data_in_1_5 : std_logic;
signal \c0.n28_adj_868\ : std_logic;
signal \c0.n26\ : std_logic;
signal \c0.data_in_frame_7_3\ : std_logic;
signal \c0.n4601\ : std_logic;
signal \c0.data_in_frame_6_3\ : std_logic;
signal \c0.data_in_frame_7_6\ : std_logic;
signal \c0.n4831\ : std_logic;
signal \tx2_data_6_keep_cascade_\ : std_logic;
signal \r_Tx_Data_6_adj_958\ : std_logic;
signal \c0.data_in_frame_6_4\ : std_logic;
signal \c0.data_in_frame_7_2\ : std_logic;
signal \c0.n4604_cascade_\ : std_logic;
signal \c0.data_in_frame_6_7\ : std_logic;
signal \c0.n4583\ : std_logic;
signal \c0.data_in_frame_7_7\ : std_logic;
signal \c0.data_in_frame_7_4\ : std_logic;
signal \c0.n4555\ : std_logic;
signal tx2_data_7_keep : std_logic;
signal \r_Tx_Data_5_adj_959\ : std_logic;
signal n4624 : std_logic;
signal \c0.n4801_cascade_\ : std_logic;
signal \tx2_data_1_keep_cascade_\ : std_logic;
signal \r_Tx_Data_1_adj_963\ : std_logic;
signal \r_Tx_Data_7_adj_957\ : std_logic;
signal n4625 : std_logic;
signal \c0.n4540\ : std_logic;
signal \c0.n4606\ : std_logic;
signal \c0.n4552\ : std_logic;
signal \c0.n4553_cascade_\ : std_logic;
signal tx2_data_5_keep : std_logic;
signal data_in_0_5 : std_logic;
signal data_in_1_0 : std_logic;
signal data_in_5_6 : std_logic;
signal \c0.n4594\ : std_logic;
signal \c0.n4825\ : std_logic;
signal \c0.n4813\ : std_logic;
signal \tx2_data_3_keep_cascade_\ : std_logic;
signal \r_Tx_Data_3_adj_961\ : std_logic;
signal \c0.n4600\ : std_logic;
signal data_in_0_6 : std_logic;
signal data_in_1_3 : std_logic;
signal data_in_0_0 : std_logic;
signal \c0.n30\ : std_logic;
signal \c0.n25_adj_870_cascade_\ : std_logic;
signal \c0.n3933\ : std_logic;
signal \c0.n1197_cascade_\ : std_logic;
signal \c0.data_in_frame_6_0\ : std_logic;
signal data_in_3_5 : std_logic;
signal \c0.data_in_frame_7_0\ : std_logic;
signal data_in_2_6 : std_logic;
signal rx_data_2 : std_logic;
signal \PIN_2_c\ : std_logic;
signal data_in_1_6 : std_logic;
signal \c0.n26_adj_869\ : std_logic;
signal data_in_2_0 : std_logic;
signal \c0.n27\ : std_logic;
signal \c0.rx.r_Rx_Data_R\ : std_logic;
signal data_in_1_4 : std_logic;
signal data_in_1_7 : std_logic;
signal n11_adj_941 : std_logic;
signal \n4638_cascade_\ : std_logic;
signal tx2_done : std_logic;
signal \c0.n4598\ : std_logic;
signal \c0.n4807\ : std_logic;
signal \tx2_data_2_keep_cascade_\ : std_logic;
signal \r_Tx_Data_2_adj_962\ : std_logic;
signal n9_adj_939 : std_logic;
signal \n4512_cascade_\ : std_logic;
signal \c0.n4546\ : std_logic;
signal \c0.n4603\ : std_logic;
signal n1611 : std_logic;
signal \n2326_cascade_\ : std_logic;
signal n4514 : std_logic;
signal n4512 : std_logic;
signal n4523 : std_logic;
signal \n4522_cascade_\ : std_logic;
signal n4777 : std_logic;
signal \r_Bit_Index_1\ : std_logic;
signal \r_Bit_Index_0_adj_956\ : std_logic;
signal \r_Bit_Index_2_adj_955\ : std_logic;
signal \c0.data_in_field_22\ : std_logic;
signal \c0.n4556\ : std_logic;
signal \c0.n10_adj_874_cascade_\ : std_logic;
signal \c0.n4567\ : std_logic;
signal data_in_0_7 : std_logic;
signal \c0.n4541\ : std_logic;
signal \c0.n4544\ : std_logic;
signal \c0.data_in_field_6\ : std_logic;
signal \c0.n1284\ : std_logic;
signal \c0.n4408_cascade_\ : std_logic;
signal \c0.n4468\ : std_logic;
signal data_in_2_3 : std_logic;
signal data_in_3_2 : std_logic;
signal data_in_2_5 : std_logic;
signal \c0.n1271_cascade_\ : std_logic;
signal \c0.n4429_cascade_\ : std_logic;
signal \c0.n4429\ : std_logic;
signal \c0.data_in_field_46\ : std_logic;
signal \c0.n6_adj_877\ : std_logic;
signal \c0.data_in_field_5\ : std_logic;
signal \c0.n4450\ : std_logic;
signal data_in_0_4 : std_logic;
signal \c0.data_in_field_31\ : std_logic;
signal \c0.n1261_cascade_\ : std_logic;
signal \c0.n4411\ : std_logic;
signal \c0.n4411_cascade_\ : std_logic;
signal \c0.data_in_frame_6_5\ : std_logic;
signal \c0.n4595\ : std_logic;
signal \c0.n1340_cascade_\ : std_logic;
signal \c0.data_in_field_16\ : std_logic;
signal \c0.data_in_field_33\ : std_logic;
signal data_in_2_2 : std_logic;
signal \c0.data_in_field_18\ : std_logic;
signal data_in_2_1 : std_logic;
signal \c0.data_in_field_17\ : std_logic;
signal \c0.data_in_field_15\ : std_logic;
signal \c0.data_in_field_27\ : std_logic;
signal \c0.n4547\ : std_logic;
signal data_in_0_3 : std_logic;
signal \c0.data_in_frame_7_5\ : std_logic;
signal \c0.data_in_field_34\ : std_logic;
signal \c0.data_in_field_3\ : std_logic;
signal \c0.data_in_field_19\ : std_logic;
signal \c0.n10\ : std_logic;
signal \c0.data_in_field_29\ : std_logic;
signal rx_data_3 : std_logic;
signal data_in_0_1 : std_logic;
signal data_in_5_5 : std_logic;
signal data_in_4_5 : std_logic;
signal \c0.rx.n4873_cascade_\ : std_logic;
signal data_in_3_7 : std_logic;
signal data_in_4_1 : std_logic;
signal data_in_3_1 : std_logic;
signal \bfn_4_21_0_\ : std_logic;
signal n1710 : std_logic;
signal \c0.tx2.n3891\ : std_logic;
signal \c0.tx2.n3892\ : std_logic;
signal \c0.tx2.n3893\ : std_logic;
signal \c0.tx2.n3894\ : std_logic;
signal n1698 : std_logic;
signal \c0.tx2.n3895\ : std_logic;
signal \c0.tx2.n3896\ : std_logic;
signal \c0.tx2.n3897\ : std_logic;
signal \c0.tx2.n3898\ : std_logic;
signal \bfn_4_22_0_\ : std_logic;
signal n1689 : std_logic;
signal n1704 : std_logic;
signal n1707 : std_logic;
signal n1768 : std_logic;
signal \c0.tx2.r_Clock_Count_0\ : std_logic;
signal \c0.tx2.r_Clock_Count_2\ : std_logic;
signal \c0.tx2.r_Clock_Count_5\ : std_logic;
signal \c0.tx2.r_Clock_Count_1\ : std_logic;
signal \c0.tx2.r_Clock_Count_3\ : std_logic;
signal \c0.tx2.n5_cascade_\ : std_logic;
signal n1701 : std_logic;
signal \c0.tx2.r_Clock_Count_4\ : std_logic;
signal n1692 : std_logic;
signal \c0.tx2.r_Clock_Count_7\ : std_logic;
signal \r_SM_Main_2_N_759_1_cascade_\ : std_logic;
signal \c0.tx2.r_Clock_Count_8\ : std_logic;
signal \c0.tx2.n2902\ : std_logic;
signal n4_adj_965 : std_logic;
signal \c0.n4543\ : std_logic;
signal blink_counter_22 : std_logic;
signal blink_counter_24 : std_logic;
signal blink_counter_21 : std_logic;
signal blink_counter_23 : std_logic;
signal \c0.n4580\ : std_logic;
signal \c0.n4571\ : std_logic;
signal \c0.n4855_cascade_\ : std_logic;
signal \tx2_data_0_keep_cascade_\ : std_logic;
signal \r_Tx_Data_0_adj_964\ : std_logic;
signal \c0.data_in_field_32\ : std_logic;
signal \c0.n4579\ : std_logic;
signal \c0.n4819\ : std_logic;
signal \c0.n4549_cascade_\ : std_logic;
signal n1030 : std_logic;
signal \tx2_data_4_keep_cascade_\ : std_logic;
signal \r_Tx_Data_4_adj_960\ : std_logic;
signal \c0.n4597\ : std_logic;
signal \c0.data_in_field_20\ : std_logic;
signal \c0.n4550\ : std_logic;
signal \c0.tx2.n23\ : std_logic;
signal \n865_cascade_\ : std_logic;
signal \r_SM_Main_2_N_759_1\ : std_logic;
signal \n4366_cascade_\ : std_logic;
signal data_in_4_2 : std_logic;
signal \c0.data_in_field_11\ : std_logic;
signal \c0.n8_adj_879_cascade_\ : std_logic;
signal \c0.n4451_cascade_\ : std_logic;
signal \c0.n8_adj_880\ : std_logic;
signal \c0.n10_adj_876\ : std_logic;
signal \c0.n4469\ : std_logic;
signal \c0.n1357_cascade_\ : std_logic;
signal \c0.n4399\ : std_logic;
signal \c0.n17\ : std_logic;
signal \c0.n4430\ : std_logic;
signal \c0.n15_adj_885\ : std_logic;
signal \c0.n16_adj_884\ : std_logic;
signal \c0.n17_adj_889_cascade_\ : std_logic;
signal \c0.n4387_cascade_\ : std_logic;
signal data_in_4_7 : std_logic;
signal data_in_5_7 : std_logic;
signal \c0.n1296\ : std_logic;
signal \c0.n11_adj_888\ : std_logic;
signal data_in_2_7 : std_logic;
signal data_in_1_1 : std_logic;
signal \c0.n8_adj_871_cascade_\ : std_logic;
signal \c0.n12\ : std_logic;
signal \c0.n1418\ : std_logic;
signal \c0.data_in_field_4\ : std_logic;
signal \c0.n1418_cascade_\ : std_logic;
signal \c0.n4474_cascade_\ : std_logic;
signal data_in_4_6 : std_logic;
signal \c0.n4396\ : std_logic;
signal \c0.data_in_field_21\ : std_logic;
signal \c0.n4396_cascade_\ : std_logic;
signal \c0.data_in_field_7\ : std_logic;
signal \c0.data_in_field_0\ : std_logic;
signal \c0.data_in_field_8\ : std_logic;
signal \c0.n4570\ : std_logic;
signal \c0.data_in_field_39\ : std_logic;
signal \c0.data_in_field_38\ : std_logic;
signal data_in_6_4 : std_logic;
signal data_in_4_4 : std_logic;
signal \c0.n8_adj_872\ : std_logic;
signal data_in_0_2 : std_logic;
signal \c0.data_in_field_2\ : std_logic;
signal \c0.data_in_frame_7_1\ : std_logic;
signal \c0.n4607\ : std_logic;
signal data_in_3_6 : std_logic;
signal \c0.data_in_frame_6_1\ : std_logic;
signal data_in_5_4 : std_logic;
signal \c0.data_in_field_44\ : std_logic;
signal data_in_3_4 : std_logic;
signal data_in_2_4 : std_logic;
signal rx_data_5 : std_logic;
signal rx_data_7 : std_logic;
signal \r_SM_Main_0_adj_954\ : std_logic;
signal \r_SM_Main_1_adj_953\ : std_logic;
signal n4780 : std_logic;
signal \r_SM_Main_2_adj_952\ : std_logic;
signal \n3_cascade_\ : std_logic;
signal rx_data_6 : std_logic;
signal \c0.rx.n4876\ : std_logic;
signal tx_enable : std_logic;
signal data_in_7_5 : std_logic;
signal data_in_6_5 : std_logic;
signal n4519 : std_logic;
signal n4520 : std_logic;
signal blink_counter_25 : std_logic;
signal \LED_c\ : std_logic;
signal \bfn_5_24_0_\ : std_logic;
signal \c0.n3921\ : std_logic;
signal \c0.n3922\ : std_logic;
signal \c0.n1675\ : std_logic;
signal \c0.n688\ : std_logic;
signal tx2_active : std_logic;
signal \c0.n2643\ : std_logic;
signal \c0.n2643_cascade_\ : std_logic;
signal \c0.tx2_transmit\ : std_logic;
signal \c0.n21\ : std_logic;
signal \c0.n22_adj_881\ : std_logic;
signal \c0.n30_adj_892_cascade_\ : std_logic;
signal \c0.n25_adj_893\ : std_logic;
signal \c0.n2637\ : std_logic;
signal \c0.n1261\ : std_logic;
signal \c0.data_in_field_45\ : std_logic;
signal \c0.n14\ : std_logic;
signal \c0.n12_adj_873\ : std_logic;
signal \c0.n16_cascade_\ : std_logic;
signal \c0.n15\ : std_logic;
signal \c0.n24\ : std_logic;
signal \c0.n4388\ : std_logic;
signal \c0.n4445\ : std_logic;
signal \c0.n26_adj_890\ : std_logic;
signal \c0.data_in_frame_6_2\ : std_logic;
signal \c0.n1280\ : std_logic;
signal \c0.n4390\ : std_logic;
signal \c0.data_in_field_47\ : std_logic;
signal \c0.n4391\ : std_logic;
signal \c0.data_in_field_1\ : std_logic;
signal \c0.data_in_field_14\ : std_logic;
signal \c0.n4474\ : std_logic;
signal \c0.n12_adj_887\ : std_logic;
signal data_in_7_7 : std_logic;
signal data_in_6_7 : std_logic;
signal \c0.data_in_field_35\ : std_logic;
signal \c0.data_in_field_36\ : std_logic;
signal \c0.n11\ : std_logic;
signal \c0.data_in_field_43\ : std_logic;
signal \c0.data_in_field_26\ : std_logic;
signal \c0.n4415_cascade_\ : std_logic;
signal \c0.data_in_field_9\ : std_logic;
signal \c0.n23\ : std_logic;
signal \c0.data_in_field_30\ : std_logic;
signal \c0.n4927\ : std_logic;
signal \c0.n1267\ : std_logic;
signal \c0.n4421\ : std_logic;
signal \c0.data_in_field_23\ : std_logic;
signal \c0.data_in_field_37\ : std_logic;
signal \c0.n8_adj_883\ : std_logic;
signal \c0.data_in_field_25\ : std_logic;
signal \c0.n1290\ : std_logic;
signal \c0.n4441\ : std_logic;
signal \c0.data_in_field_28\ : std_logic;
signal \c0.data_in_field_42\ : std_logic;
signal \c0.data_in_field_13\ : std_logic;
signal \c0.n4414\ : std_logic;
signal data_in_7_3 : std_logic;
signal data_in_7_6 : std_logic;
signal tx2_o_adj_949 : std_logic;
signal tx2_enable : std_logic;
signal \c0.data_in_field_12\ : std_logic;
signal \c0.data_in_field_40\ : std_logic;
signal data_in_6_6 : std_logic;
signal \c0.data_in_field_41\ : std_logic;
signal \c0.n12_adj_878\ : std_logic;
signal rx_data_4 : std_logic;
signal data_in_7_4 : std_logic;
signal data_in_3_0 : std_logic;
signal \c0.data_in_field_24\ : std_logic;
signal data_in_1_2 : std_logic;
signal \c0.n1197\ : std_logic;
signal \c0.FRAME_MATCHER_wait_for_transmission\ : std_logic;
signal \c0.data_in_field_10\ : std_logic;
signal n2651 : std_logic;
signal data_in_5_0 : std_logic;
signal data_in_4_0 : std_logic;
signal data_in_4_3 : std_logic;
signal data_in_3_3 : std_logic;
signal data_in_5_2 : std_logic;
signal n1222 : std_logic;
signal \n1222_cascade_\ : std_logic;
signal rx_data_0 : std_logic;
signal n4_adj_950 : std_logic;
signal n4 : std_logic;
signal \c0.rx.n2269\ : std_logic;
signal \c0.rx.n2269_cascade_\ : std_logic;
signal n1227 : std_logic;
signal \n1227_cascade_\ : std_logic;
signal \bfn_5_32_0_\ : std_logic;
signal \c0.rx.n3884\ : std_logic;
signal \c0.rx.n3885\ : std_logic;
signal \c0.rx.n3886\ : std_logic;
signal \c0.rx.n3887\ : std_logic;
signal \c0.rx.n3888\ : std_logic;
signal \c0.rx.n3889\ : std_logic;
signal \c0.rx.n3890\ : std_logic;
signal n1695 : std_logic;
signal n6_adj_940 : std_logic;
signal \c0.tx2.r_Clock_Count_6\ : std_logic;
signal \bfn_6_25_0_\ : std_logic;
signal \c0.n3906\ : std_logic;
signal \c0.n3907\ : std_logic;
signal \c0.n3908\ : std_logic;
signal \c0.n3909\ : std_logic;
signal \c0.n3910\ : std_logic;
signal \c0.n3911\ : std_logic;
signal \c0.n3912\ : std_logic;
signal \c0.n3913\ : std_logic;
signal \bfn_6_26_0_\ : std_logic;
signal \c0.n3914\ : std_logic;
signal \c0.n3915\ : std_logic;
signal \c0.n3916\ : std_logic;
signal \c0.n3917\ : std_logic;
signal \c0.n3918\ : std_logic;
signal \c0.n3919\ : std_logic;
signal \c0.n3920\ : std_logic;
signal \c0.byte_transmit_counter2_2\ : std_logic;
signal \c0.byte_transmit_counter2_1\ : std_logic;
signal \c0.byte_transmit_counter2_0\ : std_logic;
signal \c0.FRAME_MATCHER_wait_for_transmission_N_423\ : std_logic;
signal \c0.data_9\ : std_logic;
signal \c0.n4619_cascade_\ : std_logic;
signal \c0.data_1\ : std_logic;
signal data_in_7_2 : std_logic;
signal data_in_6_2 : std_logic;
signal \c0.n4517_cascade_\ : std_logic;
signal \c0.n4867_cascade_\ : std_logic;
signal \tx_data_2_keep_cascade_\ : std_logic;
signal \c0.n4564\ : std_logic;
signal \c0.n4408\ : std_logic;
signal \c0.n1271\ : std_logic;
signal \c0.n4409\ : std_logic;
signal \c0.rx.n232_cascade_\ : std_logic;
signal \c0.n4516\ : std_logic;
signal \c0.rx.n1464_cascade_\ : std_logic;
signal n1527 : std_logic;
signal \n1527_cascade_\ : std_logic;
signal n2142 : std_logic;
signal data_in_7_0 : std_logic;
signal data_in_6_0 : std_logic;
signal \c0.rx.n232\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_816_2_cascade_\ : std_logic;
signal \c0.rx.n4678\ : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal n4_adj_943 : std_logic;
signal n223 : std_logic;
signal \c0.rx.n214\ : std_logic;
signal \r_Clock_Count_3\ : std_logic;
signal \c0.rx.n214_cascade_\ : std_logic;
signal \c0.rx.n4_cascade_\ : std_logic;
signal \r_Bit_Index_2\ : std_logic;
signal \c0.rx.r_Bit_Index_1\ : std_logic;
signal n4_adj_951 : std_logic;
signal \c0.rx.n4679\ : std_logic;
signal \c0.rx.r_Clock_Count_1\ : std_logic;
signal n219 : std_logic;
signal \r_Clock_Count_7\ : std_logic;
signal \c0.rx.n4677\ : std_logic;
signal n226 : std_logic;
signal \n573_cascade_\ : std_logic;
signal \r_Clock_Count_0\ : std_logic;
signal n222 : std_logic;
signal \r_Clock_Count_4\ : std_logic;
signal \c0.rx.n4641_cascade_\ : std_logic;
signal \c0.rx.n8\ : std_logic;
signal \c0.rx.n4\ : std_logic;
signal \c0.rx.n7\ : std_logic;
signal \c0.rx.n4093_cascade_\ : std_logic;
signal \c0.rx.n2246\ : std_logic;
signal n221 : std_logic;
signal \r_Clock_Count_5\ : std_logic;
signal \c0.n4783_cascade_\ : std_logic;
signal \c0.n4526\ : std_logic;
signal \tx_data_3_keep_cascade_\ : std_logic;
signal \c0.n4622\ : std_logic;
signal \c0.n4621\ : std_logic;
signal \c0.n4525\ : std_logic;
signal data_in_6_3 : std_logic;
signal data_in_5_3 : std_logic;
signal \c0.n4768_cascade_\ : std_logic;
signal \tx_data_7_keep_cascade_\ : std_logic;
signal \c0.n4843_cascade_\ : std_logic;
signal \tx_data_1_keep_cascade_\ : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal \c0.n4585\ : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal \c0.n4861_cascade_\ : std_logic;
signal \tx_data_0_keep_cascade_\ : std_logic;
signal \c0.n4586\ : std_logic;
signal \c0.n4573\ : std_logic;
signal \c0.n4789\ : std_logic;
signal \tx_data_4_keep_cascade_\ : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal \c0.n4576\ : std_logic;
signal \c0.tx.n4589\ : std_logic;
signal \c0.tx.n4588\ : std_logic;
signal \tx_data_5_keep_cascade_\ : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal \c0.tx.n1588\ : std_logic;
signal \c0.tx.n4715_cascade_\ : std_logic;
signal rx_data_1 : std_logic;
signal data_in_7_1 : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal \r_Tx_Data_0\ : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal \c0.tx.n4558\ : std_logic;
signal \c0.tx.n4559_cascade_\ : std_logic;
signal \c0.tx.n4837\ : std_logic;
signal tx_o : std_logic;
signal rx_data_ready_keep : std_logic;
signal data_in_6_1 : std_logic;
signal data_in_5_1 : std_logic;
signal n224 : std_logic;
signal \r_Clock_Count_2\ : std_logic;
signal \c0.n4528\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_816_2\ : std_logic;
signal \c0.rx.n1024\ : std_logic;
signal \c0.tx.o_Tx_Serial_N_790\ : std_logic;
signal \c0.tx.n12\ : std_logic;
signal \c0.rx.n6_cascade_\ : std_logic;
signal \c0.rx.n357\ : std_logic;
signal \c0.rx.n4093\ : std_logic;
signal \c0.rx.n4378\ : std_logic;
signal \c0.rx.n13_cascade_\ : std_logic;
signal \c0.rx.n6\ : std_logic;
signal n1554 : std_logic;
signal n220 : std_logic;
signal n573 : std_logic;
signal \n1554_cascade_\ : std_logic;
signal \r_Clock_Count_6\ : std_logic;
signal \c0.rx.n2179\ : std_logic;
signal \c0.rx.r_SM_Main_0\ : std_logic;
signal \r_Rx_Data\ : std_logic;
signal \c0.rx.r_SM_Main_2\ : std_logic;
signal \c0.rx.n4666_cascade_\ : std_logic;
signal \c0.rx.n4667\ : std_logic;
signal \c0.rx.r_SM_Main_1\ : std_logic;
signal \bfn_9_25_0_\ : std_logic;
signal \c0.n3899\ : std_logic;
signal \c0.n3900\ : std_logic;
signal \c0.n3901\ : std_logic;
signal \c0.n3902\ : std_logic;
signal \c0.n3903\ : std_logic;
signal \c0.n3904\ : std_logic;
signal \c0.n3905\ : std_logic;
signal data_out_6_1 : std_logic;
signal \c0.data_15\ : std_logic;
signal \c0.n4888\ : std_logic;
signal \c0.n2429\ : std_logic;
signal \c0.data_6\ : std_logic;
signal \c0.data_7\ : std_logic;
signal \c0.data_14\ : std_logic;
signal data_out_7_3 : std_logic;
signal \c0.data_8\ : std_logic;
signal \n8_adj_932_cascade_\ : std_logic;
signal data_out_7_2 : std_logic;
signal data_out_7_1 : std_logic;
signal \c0.n4574\ : std_logic;
signal \c0.data_10\ : std_logic;
signal data_out_field_19 : std_logic;
signal n8_adj_936 : std_logic;
signal data_out_6_2 : std_logic;
signal \c0.n4565\ : std_logic;
signal \n11_adj_967_cascade_\ : std_logic;
signal data_out_7_4 : std_logic;
signal data_out_field_11 : std_logic;
signal \c0.n6_cascade_\ : std_logic;
signal data_out_field_24 : std_logic;
signal \c0.n4456_cascade_\ : std_logic;
signal \c0.data_0\ : std_logic;
signal data_out_field_17 : std_logic;
signal \c0.n4562\ : std_logic;
signal \c0.data_out_field_47_N_682_41\ : std_logic;
signal \c0.data_out_field_47_N_682_34\ : std_logic;
signal \c0.n1384_cascade_\ : std_logic;
signal \c0.data_out_field_47_N_682_32\ : std_logic;
signal data_out_field_3 : std_logic;
signal data_out_field_4 : std_logic;
signal \c0.n4529\ : std_logic;
signal n7_adj_937 : std_logic;
signal \c0.delay_counter_6\ : std_logic;
signal \c0.delay_counter_0\ : std_logic;
signal \c0.delay_counter_2\ : std_logic;
signal \c0.delay_counter_4\ : std_logic;
signal \c0.delay_counter_5\ : std_logic;
signal \c0.delay_counter_1\ : std_logic;
signal \c0.delay_counter_7\ : std_logic;
signal \c0.delay_counter_3\ : std_logic;
signal \c0.n13\ : std_logic;
signal \c0.n14_adj_902_cascade_\ : std_logic;
signal \c0.data_4\ : std_logic;
signal \n3580_cascade_\ : std_logic;
signal \c0.data_11\ : std_logic;
signal \c0.data_3\ : std_logic;
signal n7_adj_933 : std_logic;
signal \c0.n4885\ : std_logic;
signal \c0.data_5\ : std_logic;
signal \c0.n6_adj_904_cascade_\ : std_logic;
signal \n7_adj_938_cascade_\ : std_logic;
signal data_out_6_3 : std_logic;
signal \c0.n4380\ : std_logic;
signal \c0.data_out_field_47_N_682_33\ : std_logic;
signal \c0.n4393\ : std_logic;
signal n12_adj_966 : std_logic;
signal \n1677_cascade_\ : std_logic;
signal data_out_6_7 : std_logic;
signal n7_adj_935 : std_logic;
signal \n8_adj_934_cascade_\ : std_logic;
signal data_out_7_7 : std_logic;
signal \c0.n1333\ : std_logic;
signal \c0.n4447_cascade_\ : std_logic;
signal n9_adj_972 : std_logic;
signal \c0.n4795\ : std_logic;
signal n11_adj_945 : std_logic;
signal n4_adj_970 : std_logic;
signal data_out_field_16 : std_logic;
signal \c0.n4447\ : std_logic;
signal \n7_adj_969_cascade_\ : std_logic;
signal \c0.tx.r_Bit_Index_2\ : std_logic;
signal \c0.tx.r_Bit_Index_1\ : std_logic;
signal \c0.tx.r_Bit_Index_0\ : std_logic;
signal data_out_6_5 : std_logic;
signal \c0.n4616\ : std_logic;
signal data_out_field_25 : std_logic;
signal \c0.data_out_field_47_N_682_40\ : std_logic;
signal \c0.n4561\ : std_logic;
signal \c0.data_2\ : std_logic;
signal \c0.n4771_cascade_\ : std_logic;
signal \c0.n4774_cascade_\ : std_logic;
signal tx_data_6_keep : std_logic;
signal n10_adj_971 : std_logic;
signal \c0.data_12\ : std_logic;
signal data_out_field_7 : std_logic;
signal data_out_field_6 : std_logic;
signal \n1246_cascade_\ : std_logic;
signal data_out_field_22 : std_logic;
signal \bfn_11_27_0_\ : std_logic;
signal \c0.n3844\ : std_logic;
signal \c0.byte_transmit_counter_2\ : std_logic;
signal \c0.n3845\ : std_logic;
signal \c0.byte_transmit_counter_3\ : std_logic;
signal \c0.tx_transmit_N_274_3\ : std_logic;
signal \c0.n3846\ : std_logic;
signal \c0.byte_transmit_counter_4\ : std_logic;
signal \c0.tx_transmit_N_274_4\ : std_logic;
signal \c0.n3847\ : std_logic;
signal \c0.byte_transmit_counter_5\ : std_logic;
signal \c0.tx_transmit_N_274_5\ : std_logic;
signal \c0.n3848\ : std_logic;
signal \c0.byte_transmit_counter_6\ : std_logic;
signal \c0.tx_transmit_N_274_6\ : std_logic;
signal \c0.n3849\ : std_logic;
signal \c0.byte_transmit_counter_7\ : std_logic;
signal \c0.n3850\ : std_logic;
signal \c0.tx_transmit_N_274_7\ : std_logic;
signal \c0.data_out_field_47_N_682_35\ : std_logic;
signal n10_adj_947 : std_logic;
signal \n9_adj_948_cascade_\ : std_logic;
signal data_out_field_27 : std_logic;
signal n4_adj_942 : std_logic;
signal \c0.n4531\ : std_logic;
signal n8_adj_968 : std_logic;
signal data_out_7_0 : std_logic;
signal data_out_6_0 : std_logic;
signal \c0.n4577\ : std_logic;
signal n1255 : std_logic;
signal data_out_6_4 : std_logic;
signal data_out_field_5 : std_logic;
signal data_out_field_18 : std_logic;
signal data_out_field_20 : std_logic;
signal data_out_field_12 : std_logic;
signal \c0.n4432_cascade_\ : std_logic;
signal \c0.n4417\ : std_logic;
signal \c0.n4483\ : std_logic;
signal \c0.n10_adj_900_cascade_\ : std_logic;
signal n4438 : std_logic;
signal \c0.n4489\ : std_logic;
signal \c0.n4532\ : std_logic;
signal n1677 : std_logic;
signal \c0.n4465\ : std_logic;
signal \c0.data_out_7_5\ : std_logic;
signal \c0.data_out_field_47_N_682_45\ : std_logic;
signal \c0.n4615\ : std_logic;
signal data_out_6_6 : std_logic;
signal data_out_7_6 : std_logic;
signal \c0.n4879_cascade_\ : std_logic;
signal \c0.data_out_field_47_N_682_46\ : std_logic;
signal \c0.n4882\ : std_logic;
signal data_out_field_13 : std_logic;
signal data_out_field_28 : std_logic;
signal \c0.data_out_field_47_N_682_44\ : std_logic;
signal \c0.data_out_field_47_N_682_36\ : std_logic;
signal \c0.n4618\ : std_logic;
signal data_out_field_21 : std_logic;
signal n1246 : std_logic;
signal n4663 : std_logic;
signal \c0.byte_transmit_counter_1\ : std_logic;
signal data_out_field_31 : std_logic;
signal \c0.byte_transmit_counter_0\ : std_logic;
signal \c0.n4765\ : std_logic;
signal data_out_field_14 : std_logic;
signal \c0.data_out_field_47_N_682_42\ : std_logic;
signal n4423 : std_logic;
signal n4462 : std_logic;
signal data_out_field_26 : std_logic;
signal n4655 : std_logic;
signal data_out_field_2 : std_logic;
signal data_out_field_43 : std_logic;
signal data_out_field_15 : std_logic;
signal data_out_field_30 : std_logic;
signal \c0.tx.n1514\ : std_logic;
signal data_out_field_38 : std_logic;
signal data_out_field_9 : std_logic;
signal \c0.data_out_field_47_N_682_39\ : std_logic;
signal n4426 : std_logic;
signal \n4426_cascade_\ : std_logic;
signal data_out_field_10 : std_logic;
signal n4659 : std_logic;
signal \c0.data_13\ : std_logic;
signal \c0.data_out_field_47_N_682_37\ : std_logic;
signal n3580 : std_logic;
signal n7_adj_938 : std_logic;
signal data_out_field_1 : std_logic;
signal data_out_field_29 : std_logic;
signal \c0.n4453\ : std_logic;
signal \c0.n1312\ : std_logic;
signal \c0.n1306_cascade_\ : std_logic;
signal \c0.data_out_field_47_N_682_47\ : std_logic;
signal n4454 : std_logic;
signal \c0.tx_active_prev\ : std_logic;
signal \c0.n50\ : std_logic;
signal \c0.tx.n2908_cascade_\ : std_logic;
signal \c0.tx.n1457_cascade_\ : std_logic;
signal \c0.tx_active\ : std_logic;
signal data_out_field_8 : std_logic;
signal data_out_field_23 : std_logic;
signal n1325 : std_logic;
signal n1025 : std_logic;
signal \c0.tx.n752\ : std_logic;
signal \c0.tx_transmit\ : std_logic;
signal data_out_field_0 : std_logic;
signal \c0.n1421\ : std_logic;
signal \c0.n1306\ : std_logic;
signal \c0.tx.n6\ : std_logic;
signal \c0.tx.n5_cascade_\ : std_logic;
signal \c0.tx.n17_cascade_\ : std_logic;
signal \c0.n1378\ : std_logic;
signal \c0.n4477\ : std_logic;
signal n4480 : std_logic;
signal \c0.n4456\ : std_logic;
signal n12_adj_944 : std_logic;
signal \n4_adj_946_cascade_\ : std_logic;
signal n88 : std_logic;
signal tx_done : std_logic;
signal \c0.tx.n84\ : std_logic;
signal \c0.tx.n3643\ : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal n4375 : std_logic;
signal \c0.tx.n25_cascade_\ : std_logic;
signal \c0.tx.n17\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal \CLK_c\ : std_logic;
signal \c0.tx.r_Clock_Count_0\ : std_logic;
signal \c0.tx.n1979\ : std_logic;
signal \bfn_14_27_0_\ : std_logic;
signal \c0.tx.r_Clock_Count_1\ : std_logic;
signal \c0.tx.n1754\ : std_logic;
signal \c0.tx.n3876\ : std_logic;
signal \c0.tx.r_Clock_Count_2\ : std_logic;
signal \c0.tx.n1751\ : std_logic;
signal \c0.tx.n3877\ : std_logic;
signal \c0.tx.r_Clock_Count_3\ : std_logic;
signal \c0.tx.n1748\ : std_logic;
signal \c0.tx.n3878\ : std_logic;
signal \c0.tx.r_Clock_Count_4\ : std_logic;
signal \c0.tx.n1745\ : std_logic;
signal \c0.tx.n3879\ : std_logic;
signal \c0.tx.r_Clock_Count_5\ : std_logic;
signal \c0.tx.n1742\ : std_logic;
signal \c0.tx.n3880\ : std_logic;
signal \c0.tx.r_Clock_Count_6\ : std_logic;
signal \c0.tx.n1739\ : std_logic;
signal \c0.tx.n3881\ : std_logic;
signal \c0.tx.r_Clock_Count_7\ : std_logic;
signal \c0.tx.n1736\ : std_logic;
signal \c0.tx.n3882\ : std_logic;
signal \c0.tx.n3883\ : std_logic;
signal \c0.tx.r_Clock_Count_8\ : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal \bfn_14_28_0_\ : std_logic;
signal \c0.tx.n1733\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \LED_wire\ : std_logic;
signal \PIN_2_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    LED <= \LED_wire\;
    \PIN_2_wire\ <= PIN_2;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23697\,
            DIN => \N__23696\,
            DOUT => \N__23695\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23697\,
            PADOUT => \N__23696\,
            PADIN => \N__23695\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12218\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23688\,
            DIN => \N__23687\,
            DOUT => \N__23686\,
            PACKAGEPIN => \PIN_2_wire\
        );

    \PIN_2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23688\,
            PADOUT => \N__23687\,
            PADIN => \N__23686\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_2_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23679\,
            DIN => \N__23678\,
            DOUT => \N__23677\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23679\,
            PADOUT => \N__23678\,
            PADIN => \N__23677\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \tx2_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23670\,
            DIN => \N__23669\,
            DOUT => \N__23668\,
            PACKAGEPIN => PIN_3
        );

    \tx2_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23670\,
            PADOUT => \N__23669\,
            PADIN => \N__23668\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14060\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__14033\
        );

    \tx_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23661\,
            DIN => \N__23660\,
            DOUT => \N__23659\,
            PACKAGEPIN => PIN_1
        );

    \tx_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23661\,
            PADOUT => \N__23660\,
            PADIN => \N__23659\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__17162\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__12317\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23652\,
            DIN => \N__23651\,
            DOUT => \N__23650\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23652\,
            PADOUT => \N__23651\,
            PADIN => \N__23650\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__5783\ : InMux
    port map (
            O => \N__23633\,
            I => \N__23628\
        );

    \I__5782\ : InMux
    port map (
            O => \N__23632\,
            I => \N__23625\
        );

    \I__5781\ : InMux
    port map (
            O => \N__23631\,
            I => \N__23622\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__23628\,
            I => \c0.tx.r_Clock_Count_4\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__23625\,
            I => \c0.tx.r_Clock_Count_4\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__23622\,
            I => \c0.tx.r_Clock_Count_4\
        );

    \I__5777\ : InMux
    port map (
            O => \N__23615\,
            I => \N__23612\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__23612\,
            I => \c0.tx.n1745\
        );

    \I__5775\ : InMux
    port map (
            O => \N__23609\,
            I => \c0.tx.n3879\
        );

    \I__5774\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23601\
        );

    \I__5773\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23598\
        );

    \I__5772\ : InMux
    port map (
            O => \N__23604\,
            I => \N__23595\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__23601\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__23598\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__23595\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__5768\ : CascadeMux
    port map (
            O => \N__23588\,
            I => \N__23585\
        );

    \I__5767\ : InMux
    port map (
            O => \N__23585\,
            I => \N__23582\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__23582\,
            I => \c0.tx.n1742\
        );

    \I__5765\ : InMux
    port map (
            O => \N__23579\,
            I => \c0.tx.n3880\
        );

    \I__5764\ : InMux
    port map (
            O => \N__23576\,
            I => \N__23571\
        );

    \I__5763\ : InMux
    port map (
            O => \N__23575\,
            I => \N__23568\
        );

    \I__5762\ : InMux
    port map (
            O => \N__23574\,
            I => \N__23565\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__23571\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__23568\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__23565\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__5758\ : InMux
    port map (
            O => \N__23558\,
            I => \N__23555\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__23555\,
            I => \c0.tx.n1739\
        );

    \I__5756\ : InMux
    port map (
            O => \N__23552\,
            I => \c0.tx.n3881\
        );

    \I__5755\ : InMux
    port map (
            O => \N__23549\,
            I => \N__23544\
        );

    \I__5754\ : InMux
    port map (
            O => \N__23548\,
            I => \N__23541\
        );

    \I__5753\ : InMux
    port map (
            O => \N__23547\,
            I => \N__23538\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__23544\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__23541\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__23538\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__5749\ : InMux
    port map (
            O => \N__23531\,
            I => \N__23528\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__23528\,
            I => \c0.tx.n1736\
        );

    \I__5747\ : InMux
    port map (
            O => \N__23525\,
            I => \c0.tx.n3882\
        );

    \I__5746\ : InMux
    port map (
            O => \N__23522\,
            I => \N__23517\
        );

    \I__5745\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23514\
        );

    \I__5744\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23511\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__23517\,
            I => \N__23508\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__23514\,
            I => \c0.tx.r_Clock_Count_8\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__23511\,
            I => \c0.tx.r_Clock_Count_8\
        );

    \I__5740\ : Odrv4
    port map (
            O => \N__23508\,
            I => \c0.tx.r_Clock_Count_8\
        );

    \I__5739\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23498\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__23498\,
            I => \N__23495\
        );

    \I__5737\ : Span4Mux_s2_v
    port map (
            O => \N__23495\,
            I => \N__23490\
        );

    \I__5736\ : CascadeMux
    port map (
            O => \N__23494\,
            I => \N__23487\
        );

    \I__5735\ : CascadeMux
    port map (
            O => \N__23493\,
            I => \N__23460\
        );

    \I__5734\ : Span4Mux_h
    port map (
            O => \N__23490\,
            I => \N__23457\
        );

    \I__5733\ : InMux
    port map (
            O => \N__23487\,
            I => \N__23454\
        );

    \I__5732\ : CascadeMux
    port map (
            O => \N__23486\,
            I => \N__23450\
        );

    \I__5731\ : CascadeMux
    port map (
            O => \N__23485\,
            I => \N__23447\
        );

    \I__5730\ : CascadeMux
    port map (
            O => \N__23484\,
            I => \N__23444\
        );

    \I__5729\ : CascadeMux
    port map (
            O => \N__23483\,
            I => \N__23441\
        );

    \I__5728\ : CascadeMux
    port map (
            O => \N__23482\,
            I => \N__23438\
        );

    \I__5727\ : CascadeMux
    port map (
            O => \N__23481\,
            I => \N__23435\
        );

    \I__5726\ : CascadeMux
    port map (
            O => \N__23480\,
            I => \N__23432\
        );

    \I__5725\ : CascadeMux
    port map (
            O => \N__23479\,
            I => \N__23429\
        );

    \I__5724\ : InMux
    port map (
            O => \N__23478\,
            I => \N__23422\
        );

    \I__5723\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23422\
        );

    \I__5722\ : InMux
    port map (
            O => \N__23476\,
            I => \N__23422\
        );

    \I__5721\ : InMux
    port map (
            O => \N__23475\,
            I => \N__23419\
        );

    \I__5720\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23416\
        );

    \I__5719\ : InMux
    port map (
            O => \N__23473\,
            I => \N__23413\
        );

    \I__5718\ : InMux
    port map (
            O => \N__23472\,
            I => \N__23408\
        );

    \I__5717\ : InMux
    port map (
            O => \N__23471\,
            I => \N__23408\
        );

    \I__5716\ : InMux
    port map (
            O => \N__23470\,
            I => \N__23405\
        );

    \I__5715\ : InMux
    port map (
            O => \N__23469\,
            I => \N__23396\
        );

    \I__5714\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23396\
        );

    \I__5713\ : InMux
    port map (
            O => \N__23467\,
            I => \N__23396\
        );

    \I__5712\ : InMux
    port map (
            O => \N__23466\,
            I => \N__23396\
        );

    \I__5711\ : InMux
    port map (
            O => \N__23465\,
            I => \N__23387\
        );

    \I__5710\ : InMux
    port map (
            O => \N__23464\,
            I => \N__23387\
        );

    \I__5709\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23387\
        );

    \I__5708\ : InMux
    port map (
            O => \N__23460\,
            I => \N__23387\
        );

    \I__5707\ : Span4Mux_v
    port map (
            O => \N__23457\,
            I => \N__23384\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__23454\,
            I => \N__23381\
        );

    \I__5705\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23378\
        );

    \I__5704\ : InMux
    port map (
            O => \N__23450\,
            I => \N__23369\
        );

    \I__5703\ : InMux
    port map (
            O => \N__23447\,
            I => \N__23369\
        );

    \I__5702\ : InMux
    port map (
            O => \N__23444\,
            I => \N__23369\
        );

    \I__5701\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23369\
        );

    \I__5700\ : InMux
    port map (
            O => \N__23438\,
            I => \N__23360\
        );

    \I__5699\ : InMux
    port map (
            O => \N__23435\,
            I => \N__23360\
        );

    \I__5698\ : InMux
    port map (
            O => \N__23432\,
            I => \N__23360\
        );

    \I__5697\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23360\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__23422\,
            I => \N__23349\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__23419\,
            I => \N__23349\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__23416\,
            I => \N__23349\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__23413\,
            I => \N__23349\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__23408\,
            I => \N__23349\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__23405\,
            I => \r_SM_Main_2\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__23396\,
            I => \r_SM_Main_2\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__23387\,
            I => \r_SM_Main_2\
        );

    \I__5688\ : Odrv4
    port map (
            O => \N__23384\,
            I => \r_SM_Main_2\
        );

    \I__5687\ : Odrv4
    port map (
            O => \N__23381\,
            I => \r_SM_Main_2\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__23378\,
            I => \r_SM_Main_2\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__23369\,
            I => \r_SM_Main_2\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__23360\,
            I => \r_SM_Main_2\
        );

    \I__5683\ : Odrv4
    port map (
            O => \N__23349\,
            I => \r_SM_Main_2\
        );

    \I__5682\ : InMux
    port map (
            O => \N__23330\,
            I => \bfn_14_28_0_\
        );

    \I__5681\ : InMux
    port map (
            O => \N__23327\,
            I => \N__23324\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__23324\,
            I => \c0.tx.n1733\
        );

    \I__5679\ : CascadeMux
    port map (
            O => \N__23321\,
            I => \n4_adj_946_cascade_\
        );

    \I__5678\ : CascadeMux
    port map (
            O => \N__23318\,
            I => \N__23310\
        );

    \I__5677\ : InMux
    port map (
            O => \N__23317\,
            I => \N__23299\
        );

    \I__5676\ : InMux
    port map (
            O => \N__23316\,
            I => \N__23299\
        );

    \I__5675\ : InMux
    port map (
            O => \N__23315\,
            I => \N__23299\
        );

    \I__5674\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23288\
        );

    \I__5673\ : InMux
    port map (
            O => \N__23313\,
            I => \N__23288\
        );

    \I__5672\ : InMux
    port map (
            O => \N__23310\,
            I => \N__23288\
        );

    \I__5671\ : InMux
    port map (
            O => \N__23309\,
            I => \N__23288\
        );

    \I__5670\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23288\
        );

    \I__5669\ : CascadeMux
    port map (
            O => \N__23307\,
            I => \N__23285\
        );

    \I__5668\ : InMux
    port map (
            O => \N__23306\,
            I => \N__23282\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__23299\,
            I => \N__23279\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__23288\,
            I => \N__23276\
        );

    \I__5665\ : InMux
    port map (
            O => \N__23285\,
            I => \N__23273\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__23282\,
            I => n88
        );

    \I__5663\ : Odrv4
    port map (
            O => \N__23279\,
            I => n88
        );

    \I__5662\ : Odrv4
    port map (
            O => \N__23276\,
            I => n88
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__23273\,
            I => n88
        );

    \I__5660\ : CascadeMux
    port map (
            O => \N__23264\,
            I => \N__23260\
        );

    \I__5659\ : InMux
    port map (
            O => \N__23263\,
            I => \N__23257\
        );

    \I__5658\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23254\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__23257\,
            I => tx_done
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__23254\,
            I => tx_done
        );

    \I__5655\ : InMux
    port map (
            O => \N__23249\,
            I => \N__23246\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__23246\,
            I => \N__23241\
        );

    \I__5653\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23238\
        );

    \I__5652\ : InMux
    port map (
            O => \N__23244\,
            I => \N__23235\
        );

    \I__5651\ : Span4Mux_v
    port map (
            O => \N__23241\,
            I => \N__23232\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__23238\,
            I => \N__23229\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__23235\,
            I => \N__23226\
        );

    \I__5648\ : Span4Mux_h
    port map (
            O => \N__23232\,
            I => \N__23221\
        );

    \I__5647\ : Span4Mux_h
    port map (
            O => \N__23229\,
            I => \N__23221\
        );

    \I__5646\ : Span4Mux_h
    port map (
            O => \N__23226\,
            I => \N__23218\
        );

    \I__5645\ : Odrv4
    port map (
            O => \N__23221\,
            I => \c0.tx.n84\
        );

    \I__5644\ : Odrv4
    port map (
            O => \N__23218\,
            I => \c0.tx.n84\
        );

    \I__5643\ : InMux
    port map (
            O => \N__23213\,
            I => \N__23210\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__23210\,
            I => \c0.tx.n3643\
        );

    \I__5641\ : InMux
    port map (
            O => \N__23207\,
            I => \N__23202\
        );

    \I__5640\ : InMux
    port map (
            O => \N__23206\,
            I => \N__23197\
        );

    \I__5639\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23194\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__23202\,
            I => \N__23190\
        );

    \I__5637\ : CascadeMux
    port map (
            O => \N__23201\,
            I => \N__23186\
        );

    \I__5636\ : CascadeMux
    port map (
            O => \N__23200\,
            I => \N__23183\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__23197\,
            I => \N__23179\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__23194\,
            I => \N__23176\
        );

    \I__5633\ : CascadeMux
    port map (
            O => \N__23193\,
            I => \N__23173\
        );

    \I__5632\ : Span4Mux_v
    port map (
            O => \N__23190\,
            I => \N__23169\
        );

    \I__5631\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23166\
        );

    \I__5630\ : InMux
    port map (
            O => \N__23186\,
            I => \N__23163\
        );

    \I__5629\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23155\
        );

    \I__5628\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23155\
        );

    \I__5627\ : Span4Mux_s3_v
    port map (
            O => \N__23179\,
            I => \N__23150\
        );

    \I__5626\ : Span4Mux_v
    port map (
            O => \N__23176\,
            I => \N__23150\
        );

    \I__5625\ : InMux
    port map (
            O => \N__23173\,
            I => \N__23145\
        );

    \I__5624\ : InMux
    port map (
            O => \N__23172\,
            I => \N__23145\
        );

    \I__5623\ : Span4Mux_h
    port map (
            O => \N__23169\,
            I => \N__23142\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__23166\,
            I => \N__23137\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__23163\,
            I => \N__23137\
        );

    \I__5620\ : InMux
    port map (
            O => \N__23162\,
            I => \N__23130\
        );

    \I__5619\ : InMux
    port map (
            O => \N__23161\,
            I => \N__23130\
        );

    \I__5618\ : InMux
    port map (
            O => \N__23160\,
            I => \N__23130\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__23155\,
            I => \N__23125\
        );

    \I__5616\ : Span4Mux_h
    port map (
            O => \N__23150\,
            I => \N__23125\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__23145\,
            I => \r_SM_Main_1\
        );

    \I__5614\ : Odrv4
    port map (
            O => \N__23142\,
            I => \r_SM_Main_1\
        );

    \I__5613\ : Odrv4
    port map (
            O => \N__23137\,
            I => \r_SM_Main_1\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__23130\,
            I => \r_SM_Main_1\
        );

    \I__5611\ : Odrv4
    port map (
            O => \N__23125\,
            I => \r_SM_Main_1\
        );

    \I__5610\ : InMux
    port map (
            O => \N__23114\,
            I => \N__23108\
        );

    \I__5609\ : InMux
    port map (
            O => \N__23113\,
            I => \N__23108\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__23108\,
            I => n4375
        );

    \I__5607\ : CascadeMux
    port map (
            O => \N__23105\,
            I => \c0.tx.n25_cascade_\
        );

    \I__5606\ : CascadeMux
    port map (
            O => \N__23102\,
            I => \N__23093\
        );

    \I__5605\ : CascadeMux
    port map (
            O => \N__23101\,
            I => \N__23090\
        );

    \I__5604\ : CascadeMux
    port map (
            O => \N__23100\,
            I => \N__23087\
        );

    \I__5603\ : CascadeMux
    port map (
            O => \N__23099\,
            I => \N__23084\
        );

    \I__5602\ : CascadeMux
    port map (
            O => \N__23098\,
            I => \N__23081\
        );

    \I__5601\ : InMux
    port map (
            O => \N__23097\,
            I => \N__23073\
        );

    \I__5600\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23073\
        );

    \I__5599\ : InMux
    port map (
            O => \N__23093\,
            I => \N__23062\
        );

    \I__5598\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23062\
        );

    \I__5597\ : InMux
    port map (
            O => \N__23087\,
            I => \N__23062\
        );

    \I__5596\ : InMux
    port map (
            O => \N__23084\,
            I => \N__23057\
        );

    \I__5595\ : InMux
    port map (
            O => \N__23081\,
            I => \N__23057\
        );

    \I__5594\ : InMux
    port map (
            O => \N__23080\,
            I => \N__23054\
        );

    \I__5593\ : InMux
    port map (
            O => \N__23079\,
            I => \N__23049\
        );

    \I__5592\ : InMux
    port map (
            O => \N__23078\,
            I => \N__23049\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__23073\,
            I => \N__23046\
        );

    \I__5590\ : InMux
    port map (
            O => \N__23072\,
            I => \N__23043\
        );

    \I__5589\ : InMux
    port map (
            O => \N__23071\,
            I => \N__23038\
        );

    \I__5588\ : InMux
    port map (
            O => \N__23070\,
            I => \N__23038\
        );

    \I__5587\ : InMux
    port map (
            O => \N__23069\,
            I => \N__23035\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__23062\,
            I => \c0.tx.n17\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__23057\,
            I => \c0.tx.n17\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__23054\,
            I => \c0.tx.n17\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__23049\,
            I => \c0.tx.n17\
        );

    \I__5582\ : Odrv4
    port map (
            O => \N__23046\,
            I => \c0.tx.n17\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__23043\,
            I => \c0.tx.n17\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__23038\,
            I => \c0.tx.n17\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__23035\,
            I => \c0.tx.n17\
        );

    \I__5578\ : InMux
    port map (
            O => \N__23018\,
            I => \N__23015\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__23015\,
            I => \N__23010\
        );

    \I__5576\ : InMux
    port map (
            O => \N__23014\,
            I => \N__23007\
        );

    \I__5575\ : InMux
    port map (
            O => \N__23013\,
            I => \N__23004\
        );

    \I__5574\ : Span4Mux_h
    port map (
            O => \N__23010\,
            I => \N__22997\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__23007\,
            I => \N__22994\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__23004\,
            I => \N__22988\
        );

    \I__5571\ : InMux
    port map (
            O => \N__23003\,
            I => \N__22979\
        );

    \I__5570\ : InMux
    port map (
            O => \N__23002\,
            I => \N__22979\
        );

    \I__5569\ : InMux
    port map (
            O => \N__23001\,
            I => \N__22979\
        );

    \I__5568\ : InMux
    port map (
            O => \N__23000\,
            I => \N__22979\
        );

    \I__5567\ : Span4Mux_h
    port map (
            O => \N__22997\,
            I => \N__22974\
        );

    \I__5566\ : Span4Mux_h
    port map (
            O => \N__22994\,
            I => \N__22974\
        );

    \I__5565\ : InMux
    port map (
            O => \N__22993\,
            I => \N__22967\
        );

    \I__5564\ : InMux
    port map (
            O => \N__22992\,
            I => \N__22967\
        );

    \I__5563\ : InMux
    port map (
            O => \N__22991\,
            I => \N__22967\
        );

    \I__5562\ : Odrv12
    port map (
            O => \N__22988\,
            I => \r_SM_Main_0\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__22979\,
            I => \r_SM_Main_0\
        );

    \I__5560\ : Odrv4
    port map (
            O => \N__22974\,
            I => \r_SM_Main_0\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__22967\,
            I => \r_SM_Main_0\
        );

    \I__5558\ : ClkMux
    port map (
            O => \N__22958\,
            I => \N__22679\
        );

    \I__5557\ : ClkMux
    port map (
            O => \N__22957\,
            I => \N__22679\
        );

    \I__5556\ : ClkMux
    port map (
            O => \N__22956\,
            I => \N__22679\
        );

    \I__5555\ : ClkMux
    port map (
            O => \N__22955\,
            I => \N__22679\
        );

    \I__5554\ : ClkMux
    port map (
            O => \N__22954\,
            I => \N__22679\
        );

    \I__5553\ : ClkMux
    port map (
            O => \N__22953\,
            I => \N__22679\
        );

    \I__5552\ : ClkMux
    port map (
            O => \N__22952\,
            I => \N__22679\
        );

    \I__5551\ : ClkMux
    port map (
            O => \N__22951\,
            I => \N__22679\
        );

    \I__5550\ : ClkMux
    port map (
            O => \N__22950\,
            I => \N__22679\
        );

    \I__5549\ : ClkMux
    port map (
            O => \N__22949\,
            I => \N__22679\
        );

    \I__5548\ : ClkMux
    port map (
            O => \N__22948\,
            I => \N__22679\
        );

    \I__5547\ : ClkMux
    port map (
            O => \N__22947\,
            I => \N__22679\
        );

    \I__5546\ : ClkMux
    port map (
            O => \N__22946\,
            I => \N__22679\
        );

    \I__5545\ : ClkMux
    port map (
            O => \N__22945\,
            I => \N__22679\
        );

    \I__5544\ : ClkMux
    port map (
            O => \N__22944\,
            I => \N__22679\
        );

    \I__5543\ : ClkMux
    port map (
            O => \N__22943\,
            I => \N__22679\
        );

    \I__5542\ : ClkMux
    port map (
            O => \N__22942\,
            I => \N__22679\
        );

    \I__5541\ : ClkMux
    port map (
            O => \N__22941\,
            I => \N__22679\
        );

    \I__5540\ : ClkMux
    port map (
            O => \N__22940\,
            I => \N__22679\
        );

    \I__5539\ : ClkMux
    port map (
            O => \N__22939\,
            I => \N__22679\
        );

    \I__5538\ : ClkMux
    port map (
            O => \N__22938\,
            I => \N__22679\
        );

    \I__5537\ : ClkMux
    port map (
            O => \N__22937\,
            I => \N__22679\
        );

    \I__5536\ : ClkMux
    port map (
            O => \N__22936\,
            I => \N__22679\
        );

    \I__5535\ : ClkMux
    port map (
            O => \N__22935\,
            I => \N__22679\
        );

    \I__5534\ : ClkMux
    port map (
            O => \N__22934\,
            I => \N__22679\
        );

    \I__5533\ : ClkMux
    port map (
            O => \N__22933\,
            I => \N__22679\
        );

    \I__5532\ : ClkMux
    port map (
            O => \N__22932\,
            I => \N__22679\
        );

    \I__5531\ : ClkMux
    port map (
            O => \N__22931\,
            I => \N__22679\
        );

    \I__5530\ : ClkMux
    port map (
            O => \N__22930\,
            I => \N__22679\
        );

    \I__5529\ : ClkMux
    port map (
            O => \N__22929\,
            I => \N__22679\
        );

    \I__5528\ : ClkMux
    port map (
            O => \N__22928\,
            I => \N__22679\
        );

    \I__5527\ : ClkMux
    port map (
            O => \N__22927\,
            I => \N__22679\
        );

    \I__5526\ : ClkMux
    port map (
            O => \N__22926\,
            I => \N__22679\
        );

    \I__5525\ : ClkMux
    port map (
            O => \N__22925\,
            I => \N__22679\
        );

    \I__5524\ : ClkMux
    port map (
            O => \N__22924\,
            I => \N__22679\
        );

    \I__5523\ : ClkMux
    port map (
            O => \N__22923\,
            I => \N__22679\
        );

    \I__5522\ : ClkMux
    port map (
            O => \N__22922\,
            I => \N__22679\
        );

    \I__5521\ : ClkMux
    port map (
            O => \N__22921\,
            I => \N__22679\
        );

    \I__5520\ : ClkMux
    port map (
            O => \N__22920\,
            I => \N__22679\
        );

    \I__5519\ : ClkMux
    port map (
            O => \N__22919\,
            I => \N__22679\
        );

    \I__5518\ : ClkMux
    port map (
            O => \N__22918\,
            I => \N__22679\
        );

    \I__5517\ : ClkMux
    port map (
            O => \N__22917\,
            I => \N__22679\
        );

    \I__5516\ : ClkMux
    port map (
            O => \N__22916\,
            I => \N__22679\
        );

    \I__5515\ : ClkMux
    port map (
            O => \N__22915\,
            I => \N__22679\
        );

    \I__5514\ : ClkMux
    port map (
            O => \N__22914\,
            I => \N__22679\
        );

    \I__5513\ : ClkMux
    port map (
            O => \N__22913\,
            I => \N__22679\
        );

    \I__5512\ : ClkMux
    port map (
            O => \N__22912\,
            I => \N__22679\
        );

    \I__5511\ : ClkMux
    port map (
            O => \N__22911\,
            I => \N__22679\
        );

    \I__5510\ : ClkMux
    port map (
            O => \N__22910\,
            I => \N__22679\
        );

    \I__5509\ : ClkMux
    port map (
            O => \N__22909\,
            I => \N__22679\
        );

    \I__5508\ : ClkMux
    port map (
            O => \N__22908\,
            I => \N__22679\
        );

    \I__5507\ : ClkMux
    port map (
            O => \N__22907\,
            I => \N__22679\
        );

    \I__5506\ : ClkMux
    port map (
            O => \N__22906\,
            I => \N__22679\
        );

    \I__5505\ : ClkMux
    port map (
            O => \N__22905\,
            I => \N__22679\
        );

    \I__5504\ : ClkMux
    port map (
            O => \N__22904\,
            I => \N__22679\
        );

    \I__5503\ : ClkMux
    port map (
            O => \N__22903\,
            I => \N__22679\
        );

    \I__5502\ : ClkMux
    port map (
            O => \N__22902\,
            I => \N__22679\
        );

    \I__5501\ : ClkMux
    port map (
            O => \N__22901\,
            I => \N__22679\
        );

    \I__5500\ : ClkMux
    port map (
            O => \N__22900\,
            I => \N__22679\
        );

    \I__5499\ : ClkMux
    port map (
            O => \N__22899\,
            I => \N__22679\
        );

    \I__5498\ : ClkMux
    port map (
            O => \N__22898\,
            I => \N__22679\
        );

    \I__5497\ : ClkMux
    port map (
            O => \N__22897\,
            I => \N__22679\
        );

    \I__5496\ : ClkMux
    port map (
            O => \N__22896\,
            I => \N__22679\
        );

    \I__5495\ : ClkMux
    port map (
            O => \N__22895\,
            I => \N__22679\
        );

    \I__5494\ : ClkMux
    port map (
            O => \N__22894\,
            I => \N__22679\
        );

    \I__5493\ : ClkMux
    port map (
            O => \N__22893\,
            I => \N__22679\
        );

    \I__5492\ : ClkMux
    port map (
            O => \N__22892\,
            I => \N__22679\
        );

    \I__5491\ : ClkMux
    port map (
            O => \N__22891\,
            I => \N__22679\
        );

    \I__5490\ : ClkMux
    port map (
            O => \N__22890\,
            I => \N__22679\
        );

    \I__5489\ : ClkMux
    port map (
            O => \N__22889\,
            I => \N__22679\
        );

    \I__5488\ : ClkMux
    port map (
            O => \N__22888\,
            I => \N__22679\
        );

    \I__5487\ : ClkMux
    port map (
            O => \N__22887\,
            I => \N__22679\
        );

    \I__5486\ : ClkMux
    port map (
            O => \N__22886\,
            I => \N__22679\
        );

    \I__5485\ : ClkMux
    port map (
            O => \N__22885\,
            I => \N__22679\
        );

    \I__5484\ : ClkMux
    port map (
            O => \N__22884\,
            I => \N__22679\
        );

    \I__5483\ : ClkMux
    port map (
            O => \N__22883\,
            I => \N__22679\
        );

    \I__5482\ : ClkMux
    port map (
            O => \N__22882\,
            I => \N__22679\
        );

    \I__5481\ : ClkMux
    port map (
            O => \N__22881\,
            I => \N__22679\
        );

    \I__5480\ : ClkMux
    port map (
            O => \N__22880\,
            I => \N__22679\
        );

    \I__5479\ : ClkMux
    port map (
            O => \N__22879\,
            I => \N__22679\
        );

    \I__5478\ : ClkMux
    port map (
            O => \N__22878\,
            I => \N__22679\
        );

    \I__5477\ : ClkMux
    port map (
            O => \N__22877\,
            I => \N__22679\
        );

    \I__5476\ : ClkMux
    port map (
            O => \N__22876\,
            I => \N__22679\
        );

    \I__5475\ : ClkMux
    port map (
            O => \N__22875\,
            I => \N__22679\
        );

    \I__5474\ : ClkMux
    port map (
            O => \N__22874\,
            I => \N__22679\
        );

    \I__5473\ : ClkMux
    port map (
            O => \N__22873\,
            I => \N__22679\
        );

    \I__5472\ : ClkMux
    port map (
            O => \N__22872\,
            I => \N__22679\
        );

    \I__5471\ : ClkMux
    port map (
            O => \N__22871\,
            I => \N__22679\
        );

    \I__5470\ : ClkMux
    port map (
            O => \N__22870\,
            I => \N__22679\
        );

    \I__5469\ : ClkMux
    port map (
            O => \N__22869\,
            I => \N__22679\
        );

    \I__5468\ : ClkMux
    port map (
            O => \N__22868\,
            I => \N__22679\
        );

    \I__5467\ : ClkMux
    port map (
            O => \N__22867\,
            I => \N__22679\
        );

    \I__5466\ : ClkMux
    port map (
            O => \N__22866\,
            I => \N__22679\
        );

    \I__5465\ : GlobalMux
    port map (
            O => \N__22679\,
            I => \N__22676\
        );

    \I__5464\ : gio2CtrlBuf
    port map (
            O => \N__22676\,
            I => \CLK_c\
        );

    \I__5463\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22669\
        );

    \I__5462\ : InMux
    port map (
            O => \N__22672\,
            I => \N__22666\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__22669\,
            I => \c0.tx.r_Clock_Count_0\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__22666\,
            I => \c0.tx.r_Clock_Count_0\
        );

    \I__5459\ : InMux
    port map (
            O => \N__22661\,
            I => \N__22658\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__22658\,
            I => \c0.tx.n1979\
        );

    \I__5457\ : InMux
    port map (
            O => \N__22655\,
            I => \bfn_14_27_0_\
        );

    \I__5456\ : InMux
    port map (
            O => \N__22652\,
            I => \N__22647\
        );

    \I__5455\ : InMux
    port map (
            O => \N__22651\,
            I => \N__22644\
        );

    \I__5454\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22641\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__22647\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__22644\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__22641\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__5450\ : InMux
    port map (
            O => \N__22634\,
            I => \N__22631\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__22631\,
            I => \c0.tx.n1754\
        );

    \I__5448\ : InMux
    port map (
            O => \N__22628\,
            I => \c0.tx.n3876\
        );

    \I__5447\ : CascadeMux
    port map (
            O => \N__22625\,
            I => \N__22620\
        );

    \I__5446\ : InMux
    port map (
            O => \N__22624\,
            I => \N__22617\
        );

    \I__5445\ : InMux
    port map (
            O => \N__22623\,
            I => \N__22614\
        );

    \I__5444\ : InMux
    port map (
            O => \N__22620\,
            I => \N__22611\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__22617\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__22614\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__22611\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__5440\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22601\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__22601\,
            I => \c0.tx.n1751\
        );

    \I__5438\ : InMux
    port map (
            O => \N__22598\,
            I => \c0.tx.n3877\
        );

    \I__5437\ : InMux
    port map (
            O => \N__22595\,
            I => \N__22590\
        );

    \I__5436\ : InMux
    port map (
            O => \N__22594\,
            I => \N__22587\
        );

    \I__5435\ : InMux
    port map (
            O => \N__22593\,
            I => \N__22584\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__22590\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__22587\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__22584\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__5431\ : InMux
    port map (
            O => \N__22577\,
            I => \N__22574\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__22574\,
            I => \c0.tx.n1748\
        );

    \I__5429\ : InMux
    port map (
            O => \N__22571\,
            I => \c0.tx.n3878\
        );

    \I__5428\ : InMux
    port map (
            O => \N__22568\,
            I => \N__22565\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__22565\,
            I => \c0.tx.n6\
        );

    \I__5426\ : CascadeMux
    port map (
            O => \N__22562\,
            I => \c0.tx.n5_cascade_\
        );

    \I__5425\ : CascadeMux
    port map (
            O => \N__22559\,
            I => \c0.tx.n17_cascade_\
        );

    \I__5424\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22553\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__22553\,
            I => \N__22550\
        );

    \I__5422\ : Odrv4
    port map (
            O => \N__22550\,
            I => \c0.n1378\
        );

    \I__5421\ : InMux
    port map (
            O => \N__22547\,
            I => \N__22544\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__22544\,
            I => \N__22541\
        );

    \I__5419\ : Span4Mux_h
    port map (
            O => \N__22541\,
            I => \N__22537\
        );

    \I__5418\ : InMux
    port map (
            O => \N__22540\,
            I => \N__22534\
        );

    \I__5417\ : Odrv4
    port map (
            O => \N__22537\,
            I => \c0.n4477\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__22534\,
            I => \c0.n4477\
        );

    \I__5415\ : CascadeMux
    port map (
            O => \N__22529\,
            I => \N__22526\
        );

    \I__5414\ : InMux
    port map (
            O => \N__22526\,
            I => \N__22522\
        );

    \I__5413\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22519\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__22522\,
            I => \N__22516\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__22519\,
            I => \N__22513\
        );

    \I__5410\ : Span4Mux_h
    port map (
            O => \N__22516\,
            I => \N__22510\
        );

    \I__5409\ : Span4Mux_h
    port map (
            O => \N__22513\,
            I => \N__22507\
        );

    \I__5408\ : Odrv4
    port map (
            O => \N__22510\,
            I => n4480
        );

    \I__5407\ : Odrv4
    port map (
            O => \N__22507\,
            I => n4480
        );

    \I__5406\ : InMux
    port map (
            O => \N__22502\,
            I => \N__22499\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__22499\,
            I => \N__22496\
        );

    \I__5404\ : Span4Mux_h
    port map (
            O => \N__22496\,
            I => \N__22493\
        );

    \I__5403\ : Odrv4
    port map (
            O => \N__22493\,
            I => \c0.n4456\
        );

    \I__5402\ : InMux
    port map (
            O => \N__22490\,
            I => \N__22487\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__22487\,
            I => \N__22484\
        );

    \I__5400\ : Odrv12
    port map (
            O => \N__22484\,
            I => n12_adj_944
        );

    \I__5399\ : CascadeMux
    port map (
            O => \N__22481\,
            I => \N__22478\
        );

    \I__5398\ : InMux
    port map (
            O => \N__22478\,
            I => \N__22472\
        );

    \I__5397\ : InMux
    port map (
            O => \N__22477\,
            I => \N__22472\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__22472\,
            I => \N__22468\
        );

    \I__5395\ : InMux
    port map (
            O => \N__22471\,
            I => \N__22465\
        );

    \I__5394\ : Span4Mux_v
    port map (
            O => \N__22468\,
            I => \N__22460\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__22465\,
            I => \N__22460\
        );

    \I__5392\ : Span4Mux_h
    port map (
            O => \N__22460\,
            I => \N__22454\
        );

    \I__5391\ : InMux
    port map (
            O => \N__22459\,
            I => \N__22451\
        );

    \I__5390\ : InMux
    port map (
            O => \N__22458\,
            I => \N__22446\
        );

    \I__5389\ : InMux
    port map (
            O => \N__22457\,
            I => \N__22446\
        );

    \I__5388\ : Odrv4
    port map (
            O => \N__22454\,
            I => \c0.tx_transmit\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__22451\,
            I => \c0.tx_transmit\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__22446\,
            I => \c0.tx_transmit\
        );

    \I__5385\ : InMux
    port map (
            O => \N__22439\,
            I => \N__22435\
        );

    \I__5384\ : InMux
    port map (
            O => \N__22438\,
            I => \N__22432\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__22435\,
            I => \N__22428\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__22432\,
            I => \N__22424\
        );

    \I__5381\ : InMux
    port map (
            O => \N__22431\,
            I => \N__22421\
        );

    \I__5380\ : Span4Mux_v
    port map (
            O => \N__22428\,
            I => \N__22418\
        );

    \I__5379\ : InMux
    port map (
            O => \N__22427\,
            I => \N__22415\
        );

    \I__5378\ : Span4Mux_v
    port map (
            O => \N__22424\,
            I => \N__22412\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__22421\,
            I => \N__22409\
        );

    \I__5376\ : Span4Mux_h
    port map (
            O => \N__22418\,
            I => \N__22406\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__22415\,
            I => \N__22401\
        );

    \I__5374\ : Span4Mux_h
    port map (
            O => \N__22412\,
            I => \N__22401\
        );

    \I__5373\ : Span4Mux_v
    port map (
            O => \N__22409\,
            I => \N__22398\
        );

    \I__5372\ : Odrv4
    port map (
            O => \N__22406\,
            I => data_out_field_0
        );

    \I__5371\ : Odrv4
    port map (
            O => \N__22401\,
            I => data_out_field_0
        );

    \I__5370\ : Odrv4
    port map (
            O => \N__22398\,
            I => data_out_field_0
        );

    \I__5369\ : InMux
    port map (
            O => \N__22391\,
            I => \N__22387\
        );

    \I__5368\ : InMux
    port map (
            O => \N__22390\,
            I => \N__22384\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__22387\,
            I => \c0.n1421\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__22384\,
            I => \c0.n1421\
        );

    \I__5365\ : InMux
    port map (
            O => \N__22379\,
            I => \N__22376\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__22376\,
            I => \c0.n1306\
        );

    \I__5363\ : InMux
    port map (
            O => \N__22373\,
            I => \N__22370\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__22370\,
            I => \N__22366\
        );

    \I__5361\ : InMux
    port map (
            O => \N__22369\,
            I => \N__22363\
        );

    \I__5360\ : Span4Mux_h
    port map (
            O => \N__22366\,
            I => \N__22360\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__22363\,
            I => \c0.n4453\
        );

    \I__5358\ : Odrv4
    port map (
            O => \N__22360\,
            I => \c0.n4453\
        );

    \I__5357\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22352\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__22352\,
            I => \N__22349\
        );

    \I__5355\ : Span4Mux_h
    port map (
            O => \N__22349\,
            I => \N__22345\
        );

    \I__5354\ : InMux
    port map (
            O => \N__22348\,
            I => \N__22342\
        );

    \I__5353\ : Odrv4
    port map (
            O => \N__22345\,
            I => \c0.n1312\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__22342\,
            I => \c0.n1312\
        );

    \I__5351\ : CascadeMux
    port map (
            O => \N__22337\,
            I => \c0.n1306_cascade_\
        );

    \I__5350\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__22331\,
            I => \N__22326\
        );

    \I__5348\ : InMux
    port map (
            O => \N__22330\,
            I => \N__22319\
        );

    \I__5347\ : InMux
    port map (
            O => \N__22329\,
            I => \N__22319\
        );

    \I__5346\ : Span4Mux_v
    port map (
            O => \N__22326\,
            I => \N__22316\
        );

    \I__5345\ : InMux
    port map (
            O => \N__22325\,
            I => \N__22311\
        );

    \I__5344\ : InMux
    port map (
            O => \N__22324\,
            I => \N__22311\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__22319\,
            I => \N__22308\
        );

    \I__5342\ : Odrv4
    port map (
            O => \N__22316\,
            I => \c0.data_out_field_47_N_682_47\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__22311\,
            I => \c0.data_out_field_47_N_682_47\
        );

    \I__5340\ : Odrv4
    port map (
            O => \N__22308\,
            I => \c0.data_out_field_47_N_682_47\
        );

    \I__5339\ : CascadeMux
    port map (
            O => \N__22301\,
            I => \N__22298\
        );

    \I__5338\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22295\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__22295\,
            I => \N__22292\
        );

    \I__5336\ : Odrv12
    port map (
            O => \N__22292\,
            I => n4454
        );

    \I__5335\ : InMux
    port map (
            O => \N__22289\,
            I => \N__22286\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__22286\,
            I => \c0.tx_active_prev\
        );

    \I__5333\ : InMux
    port map (
            O => \N__22283\,
            I => \N__22280\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__22280\,
            I => \c0.n50\
        );

    \I__5331\ : CascadeMux
    port map (
            O => \N__22277\,
            I => \c0.tx.n2908_cascade_\
        );

    \I__5330\ : CascadeMux
    port map (
            O => \N__22274\,
            I => \c0.tx.n1457_cascade_\
        );

    \I__5329\ : InMux
    port map (
            O => \N__22271\,
            I => \N__22266\
        );

    \I__5328\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22261\
        );

    \I__5327\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22261\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__22266\,
            I => \N__22258\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__22261\,
            I => \N__22255\
        );

    \I__5324\ : Span4Mux_v
    port map (
            O => \N__22258\,
            I => \N__22249\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__22255\,
            I => \N__22246\
        );

    \I__5322\ : InMux
    port map (
            O => \N__22254\,
            I => \N__22239\
        );

    \I__5321\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22239\
        );

    \I__5320\ : InMux
    port map (
            O => \N__22252\,
            I => \N__22239\
        );

    \I__5319\ : Odrv4
    port map (
            O => \N__22249\,
            I => \c0.tx_active\
        );

    \I__5318\ : Odrv4
    port map (
            O => \N__22246\,
            I => \c0.tx_active\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__22239\,
            I => \c0.tx_active\
        );

    \I__5316\ : InMux
    port map (
            O => \N__22232\,
            I => \N__22228\
        );

    \I__5315\ : InMux
    port map (
            O => \N__22231\,
            I => \N__22225\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__22228\,
            I => \N__22222\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__22225\,
            I => \N__22218\
        );

    \I__5312\ : Span4Mux_v
    port map (
            O => \N__22222\,
            I => \N__22215\
        );

    \I__5311\ : InMux
    port map (
            O => \N__22221\,
            I => \N__22211\
        );

    \I__5310\ : Span4Mux_h
    port map (
            O => \N__22218\,
            I => \N__22208\
        );

    \I__5309\ : Span4Mux_h
    port map (
            O => \N__22215\,
            I => \N__22205\
        );

    \I__5308\ : InMux
    port map (
            O => \N__22214\,
            I => \N__22202\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__22211\,
            I => data_out_field_8
        );

    \I__5306\ : Odrv4
    port map (
            O => \N__22208\,
            I => data_out_field_8
        );

    \I__5305\ : Odrv4
    port map (
            O => \N__22205\,
            I => data_out_field_8
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__22202\,
            I => data_out_field_8
        );

    \I__5303\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22188\
        );

    \I__5302\ : InMux
    port map (
            O => \N__22192\,
            I => \N__22184\
        );

    \I__5301\ : InMux
    port map (
            O => \N__22191\,
            I => \N__22181\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__22188\,
            I => \N__22178\
        );

    \I__5299\ : InMux
    port map (
            O => \N__22187\,
            I => \N__22175\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__22184\,
            I => data_out_field_23
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__22181\,
            I => data_out_field_23
        );

    \I__5296\ : Odrv4
    port map (
            O => \N__22178\,
            I => data_out_field_23
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__22175\,
            I => data_out_field_23
        );

    \I__5294\ : InMux
    port map (
            O => \N__22166\,
            I => \N__22163\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__22163\,
            I => \N__22159\
        );

    \I__5292\ : InMux
    port map (
            O => \N__22162\,
            I => \N__22156\
        );

    \I__5291\ : Odrv4
    port map (
            O => \N__22159\,
            I => n1325
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__22156\,
            I => n1325
        );

    \I__5289\ : InMux
    port map (
            O => \N__22151\,
            I => \N__22147\
        );

    \I__5288\ : InMux
    port map (
            O => \N__22150\,
            I => \N__22144\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__22147\,
            I => \N__22138\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__22144\,
            I => \N__22135\
        );

    \I__5285\ : InMux
    port map (
            O => \N__22143\,
            I => \N__22132\
        );

    \I__5284\ : InMux
    port map (
            O => \N__22142\,
            I => \N__22127\
        );

    \I__5283\ : InMux
    port map (
            O => \N__22141\,
            I => \N__22127\
        );

    \I__5282\ : Span4Mux_v
    port map (
            O => \N__22138\,
            I => \N__22120\
        );

    \I__5281\ : Span4Mux_h
    port map (
            O => \N__22135\,
            I => \N__22120\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__22132\,
            I => \N__22120\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__22127\,
            I => \N__22117\
        );

    \I__5278\ : Span4Mux_v
    port map (
            O => \N__22120\,
            I => \N__22109\
        );

    \I__5277\ : Span4Mux_v
    port map (
            O => \N__22117\,
            I => \N__22109\
        );

    \I__5276\ : InMux
    port map (
            O => \N__22116\,
            I => \N__22106\
        );

    \I__5275\ : InMux
    port map (
            O => \N__22115\,
            I => \N__22101\
        );

    \I__5274\ : InMux
    port map (
            O => \N__22114\,
            I => \N__22101\
        );

    \I__5273\ : Span4Mux_h
    port map (
            O => \N__22109\,
            I => \N__22098\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__22106\,
            I => \N__22093\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__22101\,
            I => \N__22093\
        );

    \I__5270\ : Odrv4
    port map (
            O => \N__22098\,
            I => n1025
        );

    \I__5269\ : Odrv12
    port map (
            O => \N__22093\,
            I => n1025
        );

    \I__5268\ : InMux
    port map (
            O => \N__22088\,
            I => \N__22085\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__22085\,
            I => \c0.tx.n752\
        );

    \I__5266\ : InMux
    port map (
            O => \N__22082\,
            I => \N__22078\
        );

    \I__5265\ : InMux
    port map (
            O => \N__22081\,
            I => \N__22075\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__22078\,
            I => \N__22072\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__22075\,
            I => n4423
        );

    \I__5262\ : Odrv4
    port map (
            O => \N__22072\,
            I => n4423
        );

    \I__5261\ : CascadeMux
    port map (
            O => \N__22067\,
            I => \N__22064\
        );

    \I__5260\ : InMux
    port map (
            O => \N__22064\,
            I => \N__22060\
        );

    \I__5259\ : InMux
    port map (
            O => \N__22063\,
            I => \N__22057\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__22060\,
            I => \N__22054\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__22057\,
            I => \N__22051\
        );

    \I__5256\ : Span4Mux_h
    port map (
            O => \N__22054\,
            I => \N__22048\
        );

    \I__5255\ : Odrv4
    port map (
            O => \N__22051\,
            I => n4462
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__22048\,
            I => n4462
        );

    \I__5253\ : InMux
    port map (
            O => \N__22043\,
            I => \N__22039\
        );

    \I__5252\ : InMux
    port map (
            O => \N__22042\,
            I => \N__22035\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__22039\,
            I => \N__22032\
        );

    \I__5250\ : InMux
    port map (
            O => \N__22038\,
            I => \N__22028\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__22035\,
            I => \N__22023\
        );

    \I__5248\ : Span4Mux_v
    port map (
            O => \N__22032\,
            I => \N__22023\
        );

    \I__5247\ : InMux
    port map (
            O => \N__22031\,
            I => \N__22020\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__22028\,
            I => \N__22017\
        );

    \I__5245\ : Odrv4
    port map (
            O => \N__22023\,
            I => data_out_field_26
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__22020\,
            I => data_out_field_26
        );

    \I__5243\ : Odrv12
    port map (
            O => \N__22017\,
            I => data_out_field_26
        );

    \I__5242\ : CascadeMux
    port map (
            O => \N__22010\,
            I => \N__22007\
        );

    \I__5241\ : InMux
    port map (
            O => \N__22007\,
            I => \N__22004\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__22004\,
            I => n4655
        );

    \I__5239\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21997\
        );

    \I__5238\ : CascadeMux
    port map (
            O => \N__22000\,
            I => \N__21993\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__21997\,
            I => \N__21987\
        );

    \I__5236\ : InMux
    port map (
            O => \N__21996\,
            I => \N__21982\
        );

    \I__5235\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21982\
        );

    \I__5234\ : InMux
    port map (
            O => \N__21992\,
            I => \N__21979\
        );

    \I__5233\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21976\
        );

    \I__5232\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21973\
        );

    \I__5231\ : Span12Mux_s10_h
    port map (
            O => \N__21987\,
            I => \N__21970\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__21982\,
            I => data_out_field_2
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__21979\,
            I => data_out_field_2
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__21976\,
            I => data_out_field_2
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__21973\,
            I => data_out_field_2
        );

    \I__5226\ : Odrv12
    port map (
            O => \N__21970\,
            I => data_out_field_2
        );

    \I__5225\ : InMux
    port map (
            O => \N__21959\,
            I => \N__21951\
        );

    \I__5224\ : InMux
    port map (
            O => \N__21958\,
            I => \N__21951\
        );

    \I__5223\ : InMux
    port map (
            O => \N__21957\,
            I => \N__21948\
        );

    \I__5222\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21945\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__21951\,
            I => \N__21940\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__21948\,
            I => \N__21940\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__21945\,
            I => data_out_field_43
        );

    \I__5218\ : Odrv12
    port map (
            O => \N__21940\,
            I => data_out_field_43
        );

    \I__5217\ : CascadeMux
    port map (
            O => \N__21935\,
            I => \N__21932\
        );

    \I__5216\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21928\
        );

    \I__5215\ : CascadeMux
    port map (
            O => \N__21931\,
            I => \N__21925\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__21928\,
            I => \N__21922\
        );

    \I__5213\ : InMux
    port map (
            O => \N__21925\,
            I => \N__21919\
        );

    \I__5212\ : Span4Mux_h
    port map (
            O => \N__21922\,
            I => \N__21912\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__21919\,
            I => \N__21912\
        );

    \I__5210\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21909\
        );

    \I__5209\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21906\
        );

    \I__5208\ : Span4Mux_h
    port map (
            O => \N__21912\,
            I => \N__21903\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__21909\,
            I => \N__21900\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__21906\,
            I => data_out_field_15
        );

    \I__5205\ : Odrv4
    port map (
            O => \N__21903\,
            I => data_out_field_15
        );

    \I__5204\ : Odrv4
    port map (
            O => \N__21900\,
            I => data_out_field_15
        );

    \I__5203\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21886\
        );

    \I__5202\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21879\
        );

    \I__5201\ : InMux
    port map (
            O => \N__21891\,
            I => \N__21879\
        );

    \I__5200\ : InMux
    port map (
            O => \N__21890\,
            I => \N__21879\
        );

    \I__5199\ : InMux
    port map (
            O => \N__21889\,
            I => \N__21876\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__21886\,
            I => \N__21873\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__21879\,
            I => \N__21867\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__21876\,
            I => \N__21867\
        );

    \I__5195\ : Span4Mux_h
    port map (
            O => \N__21873\,
            I => \N__21864\
        );

    \I__5194\ : InMux
    port map (
            O => \N__21872\,
            I => \N__21861\
        );

    \I__5193\ : Odrv4
    port map (
            O => \N__21867\,
            I => data_out_field_30
        );

    \I__5192\ : Odrv4
    port map (
            O => \N__21864\,
            I => data_out_field_30
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__21861\,
            I => data_out_field_30
        );

    \I__5190\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21847\
        );

    \I__5189\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21847\
        );

    \I__5188\ : InMux
    port map (
            O => \N__21852\,
            I => \N__21844\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__21847\,
            I => \N__21841\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__21844\,
            I => \N__21838\
        );

    \I__5185\ : Span4Mux_h
    port map (
            O => \N__21841\,
            I => \N__21835\
        );

    \I__5184\ : Span4Mux_h
    port map (
            O => \N__21838\,
            I => \N__21832\
        );

    \I__5183\ : Span4Mux_h
    port map (
            O => \N__21835\,
            I => \N__21829\
        );

    \I__5182\ : Odrv4
    port map (
            O => \N__21832\,
            I => \c0.tx.n1514\
        );

    \I__5181\ : Odrv4
    port map (
            O => \N__21829\,
            I => \c0.tx.n1514\
        );

    \I__5180\ : InMux
    port map (
            O => \N__21824\,
            I => \N__21819\
        );

    \I__5179\ : InMux
    port map (
            O => \N__21823\,
            I => \N__21816\
        );

    \I__5178\ : InMux
    port map (
            O => \N__21822\,
            I => \N__21811\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__21819\,
            I => \N__21808\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__21816\,
            I => \N__21805\
        );

    \I__5175\ : InMux
    port map (
            O => \N__21815\,
            I => \N__21802\
        );

    \I__5174\ : InMux
    port map (
            O => \N__21814\,
            I => \N__21799\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__21811\,
            I => \N__21796\
        );

    \I__5172\ : Span4Mux_h
    port map (
            O => \N__21808\,
            I => \N__21793\
        );

    \I__5171\ : Span4Mux_h
    port map (
            O => \N__21805\,
            I => \N__21788\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__21802\,
            I => \N__21788\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__21799\,
            I => data_out_field_38
        );

    \I__5168\ : Odrv12
    port map (
            O => \N__21796\,
            I => data_out_field_38
        );

    \I__5167\ : Odrv4
    port map (
            O => \N__21793\,
            I => data_out_field_38
        );

    \I__5166\ : Odrv4
    port map (
            O => \N__21788\,
            I => data_out_field_38
        );

    \I__5165\ : CascadeMux
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__5164\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21772\
        );

    \I__5163\ : InMux
    port map (
            O => \N__21775\,
            I => \N__21769\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__21772\,
            I => \N__21764\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__21769\,
            I => \N__21761\
        );

    \I__5160\ : InMux
    port map (
            O => \N__21768\,
            I => \N__21758\
        );

    \I__5159\ : InMux
    port map (
            O => \N__21767\,
            I => \N__21755\
        );

    \I__5158\ : Span4Mux_h
    port map (
            O => \N__21764\,
            I => \N__21752\
        );

    \I__5157\ : Span4Mux_v
    port map (
            O => \N__21761\,
            I => \N__21749\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__21758\,
            I => data_out_field_9
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__21755\,
            I => data_out_field_9
        );

    \I__5154\ : Odrv4
    port map (
            O => \N__21752\,
            I => data_out_field_9
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__21749\,
            I => data_out_field_9
        );

    \I__5152\ : CascadeMux
    port map (
            O => \N__21740\,
            I => \N__21737\
        );

    \I__5151\ : InMux
    port map (
            O => \N__21737\,
            I => \N__21732\
        );

    \I__5150\ : InMux
    port map (
            O => \N__21736\,
            I => \N__21729\
        );

    \I__5149\ : CascadeMux
    port map (
            O => \N__21735\,
            I => \N__21725\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__21732\,
            I => \N__21721\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__21729\,
            I => \N__21718\
        );

    \I__5146\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21715\
        );

    \I__5145\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21710\
        );

    \I__5144\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21710\
        );

    \I__5143\ : Span4Mux_v
    port map (
            O => \N__21721\,
            I => \N__21707\
        );

    \I__5142\ : Span4Mux_h
    port map (
            O => \N__21718\,
            I => \N__21704\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__21715\,
            I => \N__21701\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__21710\,
            I => \c0.data_out_field_47_N_682_39\
        );

    \I__5139\ : Odrv4
    port map (
            O => \N__21707\,
            I => \c0.data_out_field_47_N_682_39\
        );

    \I__5138\ : Odrv4
    port map (
            O => \N__21704\,
            I => \c0.data_out_field_47_N_682_39\
        );

    \I__5137\ : Odrv12
    port map (
            O => \N__21701\,
            I => \c0.data_out_field_47_N_682_39\
        );

    \I__5136\ : InMux
    port map (
            O => \N__21692\,
            I => \N__21689\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__21689\,
            I => \N__21686\
        );

    \I__5134\ : Odrv12
    port map (
            O => \N__21686\,
            I => n4426
        );

    \I__5133\ : CascadeMux
    port map (
            O => \N__21683\,
            I => \n4426_cascade_\
        );

    \I__5132\ : InMux
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__21677\,
            I => \N__21673\
        );

    \I__5130\ : InMux
    port map (
            O => \N__21676\,
            I => \N__21668\
        );

    \I__5129\ : Span4Mux_v
    port map (
            O => \N__21673\,
            I => \N__21665\
        );

    \I__5128\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21662\
        );

    \I__5127\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21659\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__21668\,
            I => \N__21656\
        );

    \I__5125\ : Span4Mux_h
    port map (
            O => \N__21665\,
            I => \N__21651\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__21662\,
            I => \N__21651\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__21659\,
            I => data_out_field_10
        );

    \I__5122\ : Odrv4
    port map (
            O => \N__21656\,
            I => data_out_field_10
        );

    \I__5121\ : Odrv4
    port map (
            O => \N__21651\,
            I => data_out_field_10
        );

    \I__5120\ : InMux
    port map (
            O => \N__21644\,
            I => \N__21641\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__21641\,
            I => \N__21638\
        );

    \I__5118\ : Span4Mux_h
    port map (
            O => \N__21638\,
            I => \N__21635\
        );

    \I__5117\ : Odrv4
    port map (
            O => \N__21635\,
            I => n4659
        );

    \I__5116\ : CascadeMux
    port map (
            O => \N__21632\,
            I => \N__21629\
        );

    \I__5115\ : InMux
    port map (
            O => \N__21629\,
            I => \N__21626\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__21626\,
            I => \N__21623\
        );

    \I__5113\ : Span4Mux_v
    port map (
            O => \N__21623\,
            I => \N__21620\
        );

    \I__5112\ : Span4Mux_h
    port map (
            O => \N__21620\,
            I => \N__21616\
        );

    \I__5111\ : InMux
    port map (
            O => \N__21619\,
            I => \N__21613\
        );

    \I__5110\ : Odrv4
    port map (
            O => \N__21616\,
            I => \c0.data_13\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__21613\,
            I => \c0.data_13\
        );

    \I__5108\ : InMux
    port map (
            O => \N__21608\,
            I => \N__21603\
        );

    \I__5107\ : InMux
    port map (
            O => \N__21607\,
            I => \N__21597\
        );

    \I__5106\ : InMux
    port map (
            O => \N__21606\,
            I => \N__21597\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__21603\,
            I => \N__21594\
        );

    \I__5104\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21591\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__21597\,
            I => \c0.data_out_field_47_N_682_37\
        );

    \I__5102\ : Odrv4
    port map (
            O => \N__21594\,
            I => \c0.data_out_field_47_N_682_37\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__21591\,
            I => \c0.data_out_field_47_N_682_37\
        );

    \I__5100\ : CascadeMux
    port map (
            O => \N__21584\,
            I => \N__21580\
        );

    \I__5099\ : InMux
    port map (
            O => \N__21583\,
            I => \N__21565\
        );

    \I__5098\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21565\
        );

    \I__5097\ : InMux
    port map (
            O => \N__21579\,
            I => \N__21565\
        );

    \I__5096\ : InMux
    port map (
            O => \N__21578\,
            I => \N__21565\
        );

    \I__5095\ : InMux
    port map (
            O => \N__21577\,
            I => \N__21565\
        );

    \I__5094\ : InMux
    port map (
            O => \N__21576\,
            I => \N__21556\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__21565\,
            I => \N__21551\
        );

    \I__5092\ : InMux
    port map (
            O => \N__21564\,
            I => \N__21546\
        );

    \I__5091\ : InMux
    port map (
            O => \N__21563\,
            I => \N__21546\
        );

    \I__5090\ : InMux
    port map (
            O => \N__21562\,
            I => \N__21533\
        );

    \I__5089\ : InMux
    port map (
            O => \N__21561\,
            I => \N__21530\
        );

    \I__5088\ : InMux
    port map (
            O => \N__21560\,
            I => \N__21527\
        );

    \I__5087\ : InMux
    port map (
            O => \N__21559\,
            I => \N__21515\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__21556\,
            I => \N__21512\
        );

    \I__5085\ : InMux
    port map (
            O => \N__21555\,
            I => \N__21509\
        );

    \I__5084\ : InMux
    port map (
            O => \N__21554\,
            I => \N__21506\
        );

    \I__5083\ : Span4Mux_v
    port map (
            O => \N__21551\,
            I => \N__21501\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__21546\,
            I => \N__21501\
        );

    \I__5081\ : InMux
    port map (
            O => \N__21545\,
            I => \N__21490\
        );

    \I__5080\ : InMux
    port map (
            O => \N__21544\,
            I => \N__21490\
        );

    \I__5079\ : InMux
    port map (
            O => \N__21543\,
            I => \N__21490\
        );

    \I__5078\ : InMux
    port map (
            O => \N__21542\,
            I => \N__21490\
        );

    \I__5077\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21490\
        );

    \I__5076\ : InMux
    port map (
            O => \N__21540\,
            I => \N__21487\
        );

    \I__5075\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21476\
        );

    \I__5074\ : InMux
    port map (
            O => \N__21538\,
            I => \N__21476\
        );

    \I__5073\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21476\
        );

    \I__5072\ : InMux
    port map (
            O => \N__21536\,
            I => \N__21476\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__21533\,
            I => \N__21473\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__21530\,
            I => \N__21470\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__21527\,
            I => \N__21467\
        );

    \I__5068\ : CascadeMux
    port map (
            O => \N__21526\,
            I => \N__21459\
        );

    \I__5067\ : InMux
    port map (
            O => \N__21525\,
            I => \N__21456\
        );

    \I__5066\ : InMux
    port map (
            O => \N__21524\,
            I => \N__21453\
        );

    \I__5065\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21450\
        );

    \I__5064\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21430\
        );

    \I__5063\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21421\
        );

    \I__5062\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21421\
        );

    \I__5061\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21421\
        );

    \I__5060\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21421\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__21515\,
            I => \N__21414\
        );

    \I__5058\ : Span4Mux_h
    port map (
            O => \N__21512\,
            I => \N__21414\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__21509\,
            I => \N__21414\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__21506\,
            I => \N__21411\
        );

    \I__5055\ : Span4Mux_h
    port map (
            O => \N__21501\,
            I => \N__21406\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__21490\,
            I => \N__21406\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__21487\,
            I => \N__21403\
        );

    \I__5052\ : InMux
    port map (
            O => \N__21486\,
            I => \N__21398\
        );

    \I__5051\ : InMux
    port map (
            O => \N__21485\,
            I => \N__21398\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__21476\,
            I => \N__21389\
        );

    \I__5049\ : Span4Mux_v
    port map (
            O => \N__21473\,
            I => \N__21389\
        );

    \I__5048\ : Span4Mux_v
    port map (
            O => \N__21470\,
            I => \N__21389\
        );

    \I__5047\ : Span4Mux_v
    port map (
            O => \N__21467\,
            I => \N__21389\
        );

    \I__5046\ : InMux
    port map (
            O => \N__21466\,
            I => \N__21384\
        );

    \I__5045\ : InMux
    port map (
            O => \N__21465\,
            I => \N__21384\
        );

    \I__5044\ : InMux
    port map (
            O => \N__21464\,
            I => \N__21375\
        );

    \I__5043\ : InMux
    port map (
            O => \N__21463\,
            I => \N__21375\
        );

    \I__5042\ : InMux
    port map (
            O => \N__21462\,
            I => \N__21375\
        );

    \I__5041\ : InMux
    port map (
            O => \N__21459\,
            I => \N__21375\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__21456\,
            I => \N__21372\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__21453\,
            I => \N__21369\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__21450\,
            I => \N__21366\
        );

    \I__5037\ : InMux
    port map (
            O => \N__21449\,
            I => \N__21361\
        );

    \I__5036\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21361\
        );

    \I__5035\ : InMux
    port map (
            O => \N__21447\,
            I => \N__21358\
        );

    \I__5034\ : InMux
    port map (
            O => \N__21446\,
            I => \N__21355\
        );

    \I__5033\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21352\
        );

    \I__5032\ : InMux
    port map (
            O => \N__21444\,
            I => \N__21349\
        );

    \I__5031\ : InMux
    port map (
            O => \N__21443\,
            I => \N__21338\
        );

    \I__5030\ : InMux
    port map (
            O => \N__21442\,
            I => \N__21338\
        );

    \I__5029\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21338\
        );

    \I__5028\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21338\
        );

    \I__5027\ : InMux
    port map (
            O => \N__21439\,
            I => \N__21338\
        );

    \I__5026\ : InMux
    port map (
            O => \N__21438\,
            I => \N__21327\
        );

    \I__5025\ : InMux
    port map (
            O => \N__21437\,
            I => \N__21327\
        );

    \I__5024\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21327\
        );

    \I__5023\ : InMux
    port map (
            O => \N__21435\,
            I => \N__21327\
        );

    \I__5022\ : InMux
    port map (
            O => \N__21434\,
            I => \N__21327\
        );

    \I__5021\ : InMux
    port map (
            O => \N__21433\,
            I => \N__21324\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__21430\,
            I => \N__21321\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__21421\,
            I => \N__21318\
        );

    \I__5018\ : Span4Mux_v
    port map (
            O => \N__21414\,
            I => \N__21315\
        );

    \I__5017\ : Span4Mux_v
    port map (
            O => \N__21411\,
            I => \N__21312\
        );

    \I__5016\ : Span4Mux_h
    port map (
            O => \N__21406\,
            I => \N__21307\
        );

    \I__5015\ : Span4Mux_h
    port map (
            O => \N__21403\,
            I => \N__21307\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__21398\,
            I => \N__21302\
        );

    \I__5013\ : Span4Mux_h
    port map (
            O => \N__21389\,
            I => \N__21302\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__21384\,
            I => \N__21289\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__21375\,
            I => \N__21289\
        );

    \I__5010\ : Span4Mux_h
    port map (
            O => \N__21372\,
            I => \N__21289\
        );

    \I__5009\ : Span4Mux_v
    port map (
            O => \N__21369\,
            I => \N__21289\
        );

    \I__5008\ : Span4Mux_v
    port map (
            O => \N__21366\,
            I => \N__21289\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__21361\,
            I => \N__21289\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__21358\,
            I => n3580
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__21355\,
            I => n3580
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__21352\,
            I => n3580
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__21349\,
            I => n3580
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__21338\,
            I => n3580
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__21327\,
            I => n3580
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__21324\,
            I => n3580
        );

    \I__4999\ : Odrv4
    port map (
            O => \N__21321\,
            I => n3580
        );

    \I__4998\ : Odrv12
    port map (
            O => \N__21318\,
            I => n3580
        );

    \I__4997\ : Odrv4
    port map (
            O => \N__21315\,
            I => n3580
        );

    \I__4996\ : Odrv4
    port map (
            O => \N__21312\,
            I => n3580
        );

    \I__4995\ : Odrv4
    port map (
            O => \N__21307\,
            I => n3580
        );

    \I__4994\ : Odrv4
    port map (
            O => \N__21302\,
            I => n3580
        );

    \I__4993\ : Odrv4
    port map (
            O => \N__21289\,
            I => n3580
        );

    \I__4992\ : InMux
    port map (
            O => \N__21260\,
            I => \N__21252\
        );

    \I__4991\ : InMux
    port map (
            O => \N__21259\,
            I => \N__21243\
        );

    \I__4990\ : InMux
    port map (
            O => \N__21258\,
            I => \N__21239\
        );

    \I__4989\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21235\
        );

    \I__4988\ : InMux
    port map (
            O => \N__21256\,
            I => \N__21229\
        );

    \I__4987\ : InMux
    port map (
            O => \N__21255\,
            I => \N__21229\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__21252\,
            I => \N__21226\
        );

    \I__4985\ : InMux
    port map (
            O => \N__21251\,
            I => \N__21221\
        );

    \I__4984\ : InMux
    port map (
            O => \N__21250\,
            I => \N__21221\
        );

    \I__4983\ : InMux
    port map (
            O => \N__21249\,
            I => \N__21216\
        );

    \I__4982\ : InMux
    port map (
            O => \N__21248\,
            I => \N__21208\
        );

    \I__4981\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21208\
        );

    \I__4980\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21205\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__21243\,
            I => \N__21202\
        );

    \I__4978\ : InMux
    port map (
            O => \N__21242\,
            I => \N__21199\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__21239\,
            I => \N__21196\
        );

    \I__4976\ : InMux
    port map (
            O => \N__21238\,
            I => \N__21193\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__21235\,
            I => \N__21190\
        );

    \I__4974\ : InMux
    port map (
            O => \N__21234\,
            I => \N__21187\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__21229\,
            I => \N__21173\
        );

    \I__4972\ : Span4Mux_h
    port map (
            O => \N__21226\,
            I => \N__21170\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__21221\,
            I => \N__21167\
        );

    \I__4970\ : InMux
    port map (
            O => \N__21220\,
            I => \N__21162\
        );

    \I__4969\ : InMux
    port map (
            O => \N__21219\,
            I => \N__21162\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__21216\,
            I => \N__21159\
        );

    \I__4967\ : InMux
    port map (
            O => \N__21215\,
            I => \N__21154\
        );

    \I__4966\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21154\
        );

    \I__4965\ : InMux
    port map (
            O => \N__21213\,
            I => \N__21128\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__21208\,
            I => \N__21125\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__21205\,
            I => \N__21114\
        );

    \I__4962\ : Span4Mux_h
    port map (
            O => \N__21202\,
            I => \N__21114\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__21199\,
            I => \N__21114\
        );

    \I__4960\ : Span4Mux_v
    port map (
            O => \N__21196\,
            I => \N__21114\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__21193\,
            I => \N__21114\
        );

    \I__4958\ : Span4Mux_h
    port map (
            O => \N__21190\,
            I => \N__21109\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__21187\,
            I => \N__21109\
        );

    \I__4956\ : InMux
    port map (
            O => \N__21186\,
            I => \N__21098\
        );

    \I__4955\ : InMux
    port map (
            O => \N__21185\,
            I => \N__21098\
        );

    \I__4954\ : InMux
    port map (
            O => \N__21184\,
            I => \N__21098\
        );

    \I__4953\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21098\
        );

    \I__4952\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21098\
        );

    \I__4951\ : InMux
    port map (
            O => \N__21181\,
            I => \N__21093\
        );

    \I__4950\ : InMux
    port map (
            O => \N__21180\,
            I => \N__21093\
        );

    \I__4949\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21084\
        );

    \I__4948\ : InMux
    port map (
            O => \N__21178\,
            I => \N__21084\
        );

    \I__4947\ : InMux
    port map (
            O => \N__21177\,
            I => \N__21084\
        );

    \I__4946\ : InMux
    port map (
            O => \N__21176\,
            I => \N__21084\
        );

    \I__4945\ : Span4Mux_h
    port map (
            O => \N__21173\,
            I => \N__21075\
        );

    \I__4944\ : Span4Mux_v
    port map (
            O => \N__21170\,
            I => \N__21075\
        );

    \I__4943\ : Span4Mux_v
    port map (
            O => \N__21167\,
            I => \N__21075\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__21162\,
            I => \N__21075\
        );

    \I__4941\ : Span4Mux_h
    port map (
            O => \N__21159\,
            I => \N__21070\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__21154\,
            I => \N__21070\
        );

    \I__4939\ : InMux
    port map (
            O => \N__21153\,
            I => \N__21059\
        );

    \I__4938\ : InMux
    port map (
            O => \N__21152\,
            I => \N__21059\
        );

    \I__4937\ : InMux
    port map (
            O => \N__21151\,
            I => \N__21059\
        );

    \I__4936\ : InMux
    port map (
            O => \N__21150\,
            I => \N__21059\
        );

    \I__4935\ : InMux
    port map (
            O => \N__21149\,
            I => \N__21059\
        );

    \I__4934\ : InMux
    port map (
            O => \N__21148\,
            I => \N__21048\
        );

    \I__4933\ : InMux
    port map (
            O => \N__21147\,
            I => \N__21048\
        );

    \I__4932\ : InMux
    port map (
            O => \N__21146\,
            I => \N__21048\
        );

    \I__4931\ : InMux
    port map (
            O => \N__21145\,
            I => \N__21048\
        );

    \I__4930\ : InMux
    port map (
            O => \N__21144\,
            I => \N__21048\
        );

    \I__4929\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21041\
        );

    \I__4928\ : InMux
    port map (
            O => \N__21142\,
            I => \N__21041\
        );

    \I__4927\ : InMux
    port map (
            O => \N__21141\,
            I => \N__21041\
        );

    \I__4926\ : InMux
    port map (
            O => \N__21140\,
            I => \N__21032\
        );

    \I__4925\ : InMux
    port map (
            O => \N__21139\,
            I => \N__21032\
        );

    \I__4924\ : InMux
    port map (
            O => \N__21138\,
            I => \N__21032\
        );

    \I__4923\ : InMux
    port map (
            O => \N__21137\,
            I => \N__21032\
        );

    \I__4922\ : InMux
    port map (
            O => \N__21136\,
            I => \N__21019\
        );

    \I__4921\ : InMux
    port map (
            O => \N__21135\,
            I => \N__21019\
        );

    \I__4920\ : InMux
    port map (
            O => \N__21134\,
            I => \N__21019\
        );

    \I__4919\ : InMux
    port map (
            O => \N__21133\,
            I => \N__21019\
        );

    \I__4918\ : InMux
    port map (
            O => \N__21132\,
            I => \N__21019\
        );

    \I__4917\ : InMux
    port map (
            O => \N__21131\,
            I => \N__21019\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__21128\,
            I => n7_adj_938
        );

    \I__4915\ : Odrv4
    port map (
            O => \N__21125\,
            I => n7_adj_938
        );

    \I__4914\ : Odrv4
    port map (
            O => \N__21114\,
            I => n7_adj_938
        );

    \I__4913\ : Odrv4
    port map (
            O => \N__21109\,
            I => n7_adj_938
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__21098\,
            I => n7_adj_938
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__21093\,
            I => n7_adj_938
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__21084\,
            I => n7_adj_938
        );

    \I__4909\ : Odrv4
    port map (
            O => \N__21075\,
            I => n7_adj_938
        );

    \I__4908\ : Odrv4
    port map (
            O => \N__21070\,
            I => n7_adj_938
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__21059\,
            I => n7_adj_938
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__21048\,
            I => n7_adj_938
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__21041\,
            I => n7_adj_938
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__21032\,
            I => n7_adj_938
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__21019\,
            I => n7_adj_938
        );

    \I__4902\ : CascadeMux
    port map (
            O => \N__20990\,
            I => \N__20986\
        );

    \I__4901\ : InMux
    port map (
            O => \N__20989\,
            I => \N__20981\
        );

    \I__4900\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20978\
        );

    \I__4899\ : InMux
    port map (
            O => \N__20985\,
            I => \N__20975\
        );

    \I__4898\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20972\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__20981\,
            I => \N__20969\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__20978\,
            I => \N__20966\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__20975\,
            I => \N__20963\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__20972\,
            I => data_out_field_1
        );

    \I__4893\ : Odrv4
    port map (
            O => \N__20969\,
            I => data_out_field_1
        );

    \I__4892\ : Odrv4
    port map (
            O => \N__20966\,
            I => data_out_field_1
        );

    \I__4891\ : Odrv4
    port map (
            O => \N__20963\,
            I => data_out_field_1
        );

    \I__4890\ : InMux
    port map (
            O => \N__20954\,
            I => \N__20951\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__20951\,
            I => \N__20947\
        );

    \I__4888\ : InMux
    port map (
            O => \N__20950\,
            I => \N__20943\
        );

    \I__4887\ : Span4Mux_v
    port map (
            O => \N__20947\,
            I => \N__20940\
        );

    \I__4886\ : InMux
    port map (
            O => \N__20946\,
            I => \N__20937\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__20943\,
            I => data_out_field_29
        );

    \I__4884\ : Odrv4
    port map (
            O => \N__20940\,
            I => data_out_field_29
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__20937\,
            I => data_out_field_29
        );

    \I__4882\ : InMux
    port map (
            O => \N__20930\,
            I => \N__20927\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__20927\,
            I => \c0.n4882\
        );

    \I__4880\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20917\
        );

    \I__4879\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20917\
        );

    \I__4878\ : InMux
    port map (
            O => \N__20922\,
            I => \N__20914\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__20917\,
            I => \N__20910\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__20914\,
            I => \N__20907\
        );

    \I__4875\ : InMux
    port map (
            O => \N__20913\,
            I => \N__20904\
        );

    \I__4874\ : Span4Mux_v
    port map (
            O => \N__20910\,
            I => \N__20901\
        );

    \I__4873\ : Span4Mux_h
    port map (
            O => \N__20907\,
            I => \N__20898\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__20904\,
            I => data_out_field_13
        );

    \I__4871\ : Odrv4
    port map (
            O => \N__20901\,
            I => data_out_field_13
        );

    \I__4870\ : Odrv4
    port map (
            O => \N__20898\,
            I => data_out_field_13
        );

    \I__4869\ : InMux
    port map (
            O => \N__20891\,
            I => \N__20887\
        );

    \I__4868\ : InMux
    port map (
            O => \N__20890\,
            I => \N__20884\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__20887\,
            I => \N__20879\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__20884\,
            I => \N__20876\
        );

    \I__4865\ : InMux
    port map (
            O => \N__20883\,
            I => \N__20873\
        );

    \I__4864\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20870\
        );

    \I__4863\ : Span4Mux_s3_v
    port map (
            O => \N__20879\,
            I => \N__20865\
        );

    \I__4862\ : Span4Mux_h
    port map (
            O => \N__20876\,
            I => \N__20865\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__20873\,
            I => data_out_field_28
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__20870\,
            I => data_out_field_28
        );

    \I__4859\ : Odrv4
    port map (
            O => \N__20865\,
            I => data_out_field_28
        );

    \I__4858\ : InMux
    port map (
            O => \N__20858\,
            I => \N__20853\
        );

    \I__4857\ : InMux
    port map (
            O => \N__20857\,
            I => \N__20850\
        );

    \I__4856\ : InMux
    port map (
            O => \N__20856\,
            I => \N__20846\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__20853\,
            I => \N__20842\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__20850\,
            I => \N__20839\
        );

    \I__4853\ : InMux
    port map (
            O => \N__20849\,
            I => \N__20836\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__20846\,
            I => \N__20833\
        );

    \I__4851\ : InMux
    port map (
            O => \N__20845\,
            I => \N__20830\
        );

    \I__4850\ : Span4Mux_v
    port map (
            O => \N__20842\,
            I => \N__20825\
        );

    \I__4849\ : Span4Mux_h
    port map (
            O => \N__20839\,
            I => \N__20825\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__20836\,
            I => \c0.data_out_field_47_N_682_44\
        );

    \I__4847\ : Odrv4
    port map (
            O => \N__20833\,
            I => \c0.data_out_field_47_N_682_44\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__20830\,
            I => \c0.data_out_field_47_N_682_44\
        );

    \I__4845\ : Odrv4
    port map (
            O => \N__20825\,
            I => \c0.data_out_field_47_N_682_44\
        );

    \I__4844\ : InMux
    port map (
            O => \N__20816\,
            I => \N__20813\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__20813\,
            I => \N__20810\
        );

    \I__4842\ : Span4Mux_h
    port map (
            O => \N__20810\,
            I => \N__20803\
        );

    \I__4841\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20800\
        );

    \I__4840\ : InMux
    port map (
            O => \N__20808\,
            I => \N__20797\
        );

    \I__4839\ : InMux
    port map (
            O => \N__20807\,
            I => \N__20792\
        );

    \I__4838\ : InMux
    port map (
            O => \N__20806\,
            I => \N__20792\
        );

    \I__4837\ : Odrv4
    port map (
            O => \N__20803\,
            I => \c0.data_out_field_47_N_682_36\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__20800\,
            I => \c0.data_out_field_47_N_682_36\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__20797\,
            I => \c0.data_out_field_47_N_682_36\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__20792\,
            I => \c0.data_out_field_47_N_682_36\
        );

    \I__4833\ : InMux
    port map (
            O => \N__20783\,
            I => \N__20780\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__20780\,
            I => \N__20777\
        );

    \I__4831\ : Span4Mux_h
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__4830\ : Span4Mux_h
    port map (
            O => \N__20774\,
            I => \N__20771\
        );

    \I__4829\ : Odrv4
    port map (
            O => \N__20771\,
            I => \c0.n4618\
        );

    \I__4828\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20765\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__20765\,
            I => \N__20761\
        );

    \I__4826\ : CascadeMux
    port map (
            O => \N__20764\,
            I => \N__20756\
        );

    \I__4825\ : Span4Mux_v
    port map (
            O => \N__20761\,
            I => \N__20752\
        );

    \I__4824\ : InMux
    port map (
            O => \N__20760\,
            I => \N__20749\
        );

    \I__4823\ : InMux
    port map (
            O => \N__20759\,
            I => \N__20742\
        );

    \I__4822\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20742\
        );

    \I__4821\ : InMux
    port map (
            O => \N__20755\,
            I => \N__20742\
        );

    \I__4820\ : Odrv4
    port map (
            O => \N__20752\,
            I => data_out_field_21
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__20749\,
            I => data_out_field_21
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__20742\,
            I => data_out_field_21
        );

    \I__4817\ : CascadeMux
    port map (
            O => \N__20735\,
            I => \N__20732\
        );

    \I__4816\ : InMux
    port map (
            O => \N__20732\,
            I => \N__20729\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__20729\,
            I => \N__20726\
        );

    \I__4814\ : Odrv4
    port map (
            O => \N__20726\,
            I => n1246
        );

    \I__4813\ : CascadeMux
    port map (
            O => \N__20723\,
            I => \N__20720\
        );

    \I__4812\ : InMux
    port map (
            O => \N__20720\,
            I => \N__20717\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__20717\,
            I => \N__20714\
        );

    \I__4810\ : Span4Mux_h
    port map (
            O => \N__20714\,
            I => \N__20711\
        );

    \I__4809\ : Odrv4
    port map (
            O => \N__20711\,
            I => n4663
        );

    \I__4808\ : InMux
    port map (
            O => \N__20708\,
            I => \N__20702\
        );

    \I__4807\ : InMux
    port map (
            O => \N__20707\,
            I => \N__20698\
        );

    \I__4806\ : InMux
    port map (
            O => \N__20706\,
            I => \N__20695\
        );

    \I__4805\ : InMux
    port map (
            O => \N__20705\,
            I => \N__20690\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__20702\,
            I => \N__20686\
        );

    \I__4803\ : InMux
    port map (
            O => \N__20701\,
            I => \N__20683\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__20698\,
            I => \N__20676\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__20695\,
            I => \N__20673\
        );

    \I__4800\ : InMux
    port map (
            O => \N__20694\,
            I => \N__20670\
        );

    \I__4799\ : InMux
    port map (
            O => \N__20693\,
            I => \N__20667\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__20690\,
            I => \N__20664\
        );

    \I__4797\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20661\
        );

    \I__4796\ : Span4Mux_v
    port map (
            O => \N__20686\,
            I => \N__20655\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__20683\,
            I => \N__20655\
        );

    \I__4794\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20650\
        );

    \I__4793\ : InMux
    port map (
            O => \N__20681\,
            I => \N__20650\
        );

    \I__4792\ : InMux
    port map (
            O => \N__20680\,
            I => \N__20645\
        );

    \I__4791\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20645\
        );

    \I__4790\ : Span4Mux_v
    port map (
            O => \N__20676\,
            I => \N__20640\
        );

    \I__4789\ : Span12Mux_s5_v
    port map (
            O => \N__20673\,
            I => \N__20633\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__20670\,
            I => \N__20633\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__20667\,
            I => \N__20633\
        );

    \I__4786\ : Span4Mux_h
    port map (
            O => \N__20664\,
            I => \N__20628\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__20661\,
            I => \N__20628\
        );

    \I__4784\ : InMux
    port map (
            O => \N__20660\,
            I => \N__20625\
        );

    \I__4783\ : Span4Mux_h
    port map (
            O => \N__20655\,
            I => \N__20620\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__20650\,
            I => \N__20620\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__20645\,
            I => \N__20617\
        );

    \I__4780\ : InMux
    port map (
            O => \N__20644\,
            I => \N__20614\
        );

    \I__4779\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20611\
        );

    \I__4778\ : Odrv4
    port map (
            O => \N__20640\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__4777\ : Odrv12
    port map (
            O => \N__20633\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__20628\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__20625\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__20620\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__4773\ : Odrv4
    port map (
            O => \N__20617\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__20614\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__20611\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__4770\ : CascadeMux
    port map (
            O => \N__20594\,
            I => \N__20591\
        );

    \I__4769\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20587\
        );

    \I__4768\ : CascadeMux
    port map (
            O => \N__20590\,
            I => \N__20584\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__20587\,
            I => \N__20580\
        );

    \I__4766\ : InMux
    port map (
            O => \N__20584\,
            I => \N__20575\
        );

    \I__4765\ : InMux
    port map (
            O => \N__20583\,
            I => \N__20572\
        );

    \I__4764\ : Span4Mux_h
    port map (
            O => \N__20580\,
            I => \N__20569\
        );

    \I__4763\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20564\
        );

    \I__4762\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20564\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__20575\,
            I => data_out_field_31
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__20572\,
            I => data_out_field_31
        );

    \I__4759\ : Odrv4
    port map (
            O => \N__20569\,
            I => data_out_field_31
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__20564\,
            I => data_out_field_31
        );

    \I__4757\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20543\
        );

    \I__4756\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20540\
        );

    \I__4755\ : InMux
    port map (
            O => \N__20553\,
            I => \N__20535\
        );

    \I__4754\ : InMux
    port map (
            O => \N__20552\,
            I => \N__20535\
        );

    \I__4753\ : InMux
    port map (
            O => \N__20551\,
            I => \N__20532\
        );

    \I__4752\ : InMux
    port map (
            O => \N__20550\,
            I => \N__20527\
        );

    \I__4751\ : InMux
    port map (
            O => \N__20549\,
            I => \N__20527\
        );

    \I__4750\ : InMux
    port map (
            O => \N__20548\,
            I => \N__20520\
        );

    \I__4749\ : InMux
    port map (
            O => \N__20547\,
            I => \N__20520\
        );

    \I__4748\ : InMux
    port map (
            O => \N__20546\,
            I => \N__20520\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__20543\,
            I => \N__20513\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__20540\,
            I => \N__20502\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__20535\,
            I => \N__20502\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__20532\,
            I => \N__20502\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__20527\,
            I => \N__20502\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__20520\,
            I => \N__20502\
        );

    \I__4741\ : InMux
    port map (
            O => \N__20519\,
            I => \N__20497\
        );

    \I__4740\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20497\
        );

    \I__4739\ : CascadeMux
    port map (
            O => \N__20517\,
            I => \N__20490\
        );

    \I__4738\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20487\
        );

    \I__4737\ : Span4Mux_s3_v
    port map (
            O => \N__20513\,
            I => \N__20480\
        );

    \I__4736\ : Span4Mux_v
    port map (
            O => \N__20502\,
            I => \N__20480\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__20497\,
            I => \N__20480\
        );

    \I__4734\ : InMux
    port map (
            O => \N__20496\,
            I => \N__20472\
        );

    \I__4733\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20472\
        );

    \I__4732\ : InMux
    port map (
            O => \N__20494\,
            I => \N__20467\
        );

    \I__4731\ : InMux
    port map (
            O => \N__20493\,
            I => \N__20467\
        );

    \I__4730\ : InMux
    port map (
            O => \N__20490\,
            I => \N__20462\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__20487\,
            I => \N__20457\
        );

    \I__4728\ : Span4Mux_h
    port map (
            O => \N__20480\,
            I => \N__20457\
        );

    \I__4727\ : InMux
    port map (
            O => \N__20479\,
            I => \N__20454\
        );

    \I__4726\ : InMux
    port map (
            O => \N__20478\,
            I => \N__20448\
        );

    \I__4725\ : InMux
    port map (
            O => \N__20477\,
            I => \N__20445\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__20472\,
            I => \N__20442\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__20467\,
            I => \N__20439\
        );

    \I__4722\ : InMux
    port map (
            O => \N__20466\,
            I => \N__20433\
        );

    \I__4721\ : InMux
    port map (
            O => \N__20465\,
            I => \N__20433\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__20462\,
            I => \N__20430\
        );

    \I__4719\ : Span4Mux_h
    port map (
            O => \N__20457\,
            I => \N__20425\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__20454\,
            I => \N__20425\
        );

    \I__4717\ : CascadeMux
    port map (
            O => \N__20453\,
            I => \N__20420\
        );

    \I__4716\ : InMux
    port map (
            O => \N__20452\,
            I => \N__20415\
        );

    \I__4715\ : InMux
    port map (
            O => \N__20451\,
            I => \N__20415\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__20448\,
            I => \N__20412\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__20445\,
            I => \N__20409\
        );

    \I__4712\ : Span4Mux_v
    port map (
            O => \N__20442\,
            I => \N__20404\
        );

    \I__4711\ : Span4Mux_v
    port map (
            O => \N__20439\,
            I => \N__20404\
        );

    \I__4710\ : InMux
    port map (
            O => \N__20438\,
            I => \N__20401\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__20433\,
            I => \N__20394\
        );

    \I__4708\ : Span4Mux_h
    port map (
            O => \N__20430\,
            I => \N__20394\
        );

    \I__4707\ : Span4Mux_s3_v
    port map (
            O => \N__20425\,
            I => \N__20394\
        );

    \I__4706\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20389\
        );

    \I__4705\ : InMux
    port map (
            O => \N__20423\,
            I => \N__20389\
        );

    \I__4704\ : InMux
    port map (
            O => \N__20420\,
            I => \N__20386\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__20415\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__4702\ : Odrv4
    port map (
            O => \N__20412\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__4701\ : Odrv4
    port map (
            O => \N__20409\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__20404\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__20401\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__4698\ : Odrv4
    port map (
            O => \N__20394\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__20389\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__20386\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__4695\ : InMux
    port map (
            O => \N__20369\,
            I => \N__20366\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__20366\,
            I => \N__20363\
        );

    \I__4693\ : Odrv12
    port map (
            O => \N__20363\,
            I => \c0.n4765\
        );

    \I__4692\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20355\
        );

    \I__4691\ : InMux
    port map (
            O => \N__20359\,
            I => \N__20350\
        );

    \I__4690\ : InMux
    port map (
            O => \N__20358\,
            I => \N__20350\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__20355\,
            I => data_out_field_14
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__20350\,
            I => data_out_field_14
        );

    \I__4687\ : CascadeMux
    port map (
            O => \N__20345\,
            I => \N__20342\
        );

    \I__4686\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20338\
        );

    \I__4685\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20335\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__20338\,
            I => \N__20332\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__20335\,
            I => \N__20329\
        );

    \I__4682\ : Span4Mux_s3_v
    port map (
            O => \N__20332\,
            I => \N__20322\
        );

    \I__4681\ : Span4Mux_h
    port map (
            O => \N__20329\,
            I => \N__20322\
        );

    \I__4680\ : InMux
    port map (
            O => \N__20328\,
            I => \N__20319\
        );

    \I__4679\ : InMux
    port map (
            O => \N__20327\,
            I => \N__20316\
        );

    \I__4678\ : Span4Mux_v
    port map (
            O => \N__20322\,
            I => \N__20313\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__20319\,
            I => \c0.data_out_field_47_N_682_42\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__20316\,
            I => \c0.data_out_field_47_N_682_42\
        );

    \I__4675\ : Odrv4
    port map (
            O => \N__20313\,
            I => \c0.data_out_field_47_N_682_42\
        );

    \I__4674\ : CascadeMux
    port map (
            O => \N__20306\,
            I => \N__20303\
        );

    \I__4673\ : InMux
    port map (
            O => \N__20303\,
            I => \N__20300\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__20300\,
            I => \N__20296\
        );

    \I__4671\ : InMux
    port map (
            O => \N__20299\,
            I => \N__20293\
        );

    \I__4670\ : Odrv4
    port map (
            O => \N__20296\,
            I => n1255
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__20293\,
            I => n1255
        );

    \I__4668\ : InMux
    port map (
            O => \N__20288\,
            I => \N__20285\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__20285\,
            I => \N__20281\
        );

    \I__4666\ : InMux
    port map (
            O => \N__20284\,
            I => \N__20278\
        );

    \I__4665\ : Span4Mux_h
    port map (
            O => \N__20281\,
            I => \N__20275\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__20278\,
            I => \N__20272\
        );

    \I__4663\ : Span4Mux_h
    port map (
            O => \N__20275\,
            I => \N__20269\
        );

    \I__4662\ : Odrv4
    port map (
            O => \N__20272\,
            I => data_out_6_4
        );

    \I__4661\ : Odrv4
    port map (
            O => \N__20269\,
            I => data_out_6_4
        );

    \I__4660\ : CascadeMux
    port map (
            O => \N__20264\,
            I => \N__20259\
        );

    \I__4659\ : InMux
    port map (
            O => \N__20263\,
            I => \N__20252\
        );

    \I__4658\ : InMux
    port map (
            O => \N__20262\,
            I => \N__20252\
        );

    \I__4657\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20247\
        );

    \I__4656\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20247\
        );

    \I__4655\ : InMux
    port map (
            O => \N__20257\,
            I => \N__20244\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__20252\,
            I => data_out_field_5
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__20247\,
            I => data_out_field_5
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__20244\,
            I => data_out_field_5
        );

    \I__4651\ : CascadeMux
    port map (
            O => \N__20237\,
            I => \N__20231\
        );

    \I__4650\ : InMux
    port map (
            O => \N__20236\,
            I => \N__20228\
        );

    \I__4649\ : InMux
    port map (
            O => \N__20235\,
            I => \N__20225\
        );

    \I__4648\ : InMux
    port map (
            O => \N__20234\,
            I => \N__20221\
        );

    \I__4647\ : InMux
    port map (
            O => \N__20231\,
            I => \N__20218\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__20228\,
            I => \N__20215\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__20225\,
            I => \N__20212\
        );

    \I__4644\ : InMux
    port map (
            O => \N__20224\,
            I => \N__20209\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__20221\,
            I => data_out_field_18
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__20218\,
            I => data_out_field_18
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__20215\,
            I => data_out_field_18
        );

    \I__4640\ : Odrv4
    port map (
            O => \N__20212\,
            I => data_out_field_18
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__20209\,
            I => data_out_field_18
        );

    \I__4638\ : InMux
    port map (
            O => \N__20198\,
            I => \N__20195\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__20195\,
            I => \N__20189\
        );

    \I__4636\ : InMux
    port map (
            O => \N__20194\,
            I => \N__20186\
        );

    \I__4635\ : InMux
    port map (
            O => \N__20193\,
            I => \N__20182\
        );

    \I__4634\ : InMux
    port map (
            O => \N__20192\,
            I => \N__20179\
        );

    \I__4633\ : Span4Mux_h
    port map (
            O => \N__20189\,
            I => \N__20174\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__20186\,
            I => \N__20174\
        );

    \I__4631\ : InMux
    port map (
            O => \N__20185\,
            I => \N__20171\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__20182\,
            I => data_out_field_20
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__20179\,
            I => data_out_field_20
        );

    \I__4628\ : Odrv4
    port map (
            O => \N__20174\,
            I => data_out_field_20
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__20171\,
            I => data_out_field_20
        );

    \I__4626\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20158\
        );

    \I__4625\ : InMux
    port map (
            O => \N__20161\,
            I => \N__20155\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__20158\,
            I => \N__20152\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__20155\,
            I => \N__20147\
        );

    \I__4622\ : Span4Mux_h
    port map (
            O => \N__20152\,
            I => \N__20144\
        );

    \I__4621\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20139\
        );

    \I__4620\ : InMux
    port map (
            O => \N__20150\,
            I => \N__20139\
        );

    \I__4619\ : Span4Mux_h
    port map (
            O => \N__20147\,
            I => \N__20136\
        );

    \I__4618\ : Odrv4
    port map (
            O => \N__20144\,
            I => data_out_field_12
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__20139\,
            I => data_out_field_12
        );

    \I__4616\ : Odrv4
    port map (
            O => \N__20136\,
            I => data_out_field_12
        );

    \I__4615\ : CascadeMux
    port map (
            O => \N__20129\,
            I => \c0.n4432_cascade_\
        );

    \I__4614\ : InMux
    port map (
            O => \N__20126\,
            I => \N__20123\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__20123\,
            I => \c0.n4417\
        );

    \I__4612\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20117\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__20117\,
            I => \N__20114\
        );

    \I__4610\ : Odrv4
    port map (
            O => \N__20114\,
            I => \c0.n4483\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__20111\,
            I => \c0.n10_adj_900_cascade_\
        );

    \I__4608\ : InMux
    port map (
            O => \N__20108\,
            I => \N__20104\
        );

    \I__4607\ : InMux
    port map (
            O => \N__20107\,
            I => \N__20101\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__20104\,
            I => \N__20096\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__20101\,
            I => \N__20096\
        );

    \I__4604\ : Odrv4
    port map (
            O => \N__20096\,
            I => n4438
        );

    \I__4603\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20087\
        );

    \I__4602\ : InMux
    port map (
            O => \N__20092\,
            I => \N__20087\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__20087\,
            I => \c0.n4489\
        );

    \I__4600\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20081\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__20081\,
            I => \N__20078\
        );

    \I__4598\ : Odrv12
    port map (
            O => \N__20078\,
            I => \c0.n4532\
        );

    \I__4597\ : CascadeMux
    port map (
            O => \N__20075\,
            I => \N__20071\
        );

    \I__4596\ : CascadeMux
    port map (
            O => \N__20074\,
            I => \N__20067\
        );

    \I__4595\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20064\
        );

    \I__4594\ : InMux
    port map (
            O => \N__20070\,
            I => \N__20050\
        );

    \I__4593\ : InMux
    port map (
            O => \N__20067\,
            I => \N__20047\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__20064\,
            I => \N__20044\
        );

    \I__4591\ : InMux
    port map (
            O => \N__20063\,
            I => \N__20041\
        );

    \I__4590\ : InMux
    port map (
            O => \N__20062\,
            I => \N__20038\
        );

    \I__4589\ : InMux
    port map (
            O => \N__20061\,
            I => \N__20035\
        );

    \I__4588\ : InMux
    port map (
            O => \N__20060\,
            I => \N__20030\
        );

    \I__4587\ : InMux
    port map (
            O => \N__20059\,
            I => \N__20030\
        );

    \I__4586\ : InMux
    port map (
            O => \N__20058\,
            I => \N__20025\
        );

    \I__4585\ : InMux
    port map (
            O => \N__20057\,
            I => \N__20025\
        );

    \I__4584\ : InMux
    port map (
            O => \N__20056\,
            I => \N__20022\
        );

    \I__4583\ : InMux
    port map (
            O => \N__20055\,
            I => \N__20019\
        );

    \I__4582\ : InMux
    port map (
            O => \N__20054\,
            I => \N__20014\
        );

    \I__4581\ : InMux
    port map (
            O => \N__20053\,
            I => \N__20014\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__20050\,
            I => n1677
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__20047\,
            I => n1677
        );

    \I__4578\ : Odrv4
    port map (
            O => \N__20044\,
            I => n1677
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__20041\,
            I => n1677
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__20038\,
            I => n1677
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__20035\,
            I => n1677
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__20030\,
            I => n1677
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__20025\,
            I => n1677
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__20022\,
            I => n1677
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__20019\,
            I => n1677
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__20014\,
            I => n1677
        );

    \I__4569\ : InMux
    port map (
            O => \N__19991\,
            I => \N__19988\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__19988\,
            I => \N__19985\
        );

    \I__4567\ : Span4Mux_h
    port map (
            O => \N__19985\,
            I => \N__19979\
        );

    \I__4566\ : InMux
    port map (
            O => \N__19984\,
            I => \N__19972\
        );

    \I__4565\ : InMux
    port map (
            O => \N__19983\,
            I => \N__19972\
        );

    \I__4564\ : InMux
    port map (
            O => \N__19982\,
            I => \N__19972\
        );

    \I__4563\ : Odrv4
    port map (
            O => \N__19979\,
            I => \c0.n4465\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__19972\,
            I => \c0.n4465\
        );

    \I__4561\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19963\
        );

    \I__4560\ : InMux
    port map (
            O => \N__19966\,
            I => \N__19960\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__19963\,
            I => \c0.data_out_7_5\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__19960\,
            I => \c0.data_out_7_5\
        );

    \I__4557\ : CascadeMux
    port map (
            O => \N__19955\,
            I => \N__19950\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__19954\,
            I => \N__19947\
        );

    \I__4555\ : InMux
    port map (
            O => \N__19953\,
            I => \N__19940\
        );

    \I__4554\ : InMux
    port map (
            O => \N__19950\,
            I => \N__19940\
        );

    \I__4553\ : InMux
    port map (
            O => \N__19947\,
            I => \N__19935\
        );

    \I__4552\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19935\
        );

    \I__4551\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19932\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__19940\,
            I => \N__19927\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__19935\,
            I => \N__19927\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__19932\,
            I => \c0.data_out_field_47_N_682_45\
        );

    \I__4547\ : Odrv4
    port map (
            O => \N__19927\,
            I => \c0.data_out_field_47_N_682_45\
        );

    \I__4546\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19919\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__19919\,
            I => \c0.n4615\
        );

    \I__4544\ : InMux
    port map (
            O => \N__19916\,
            I => \N__19912\
        );

    \I__4543\ : InMux
    port map (
            O => \N__19915\,
            I => \N__19909\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__19912\,
            I => data_out_6_6
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__19909\,
            I => data_out_6_6
        );

    \I__4540\ : InMux
    port map (
            O => \N__19904\,
            I => \N__19900\
        );

    \I__4539\ : InMux
    port map (
            O => \N__19903\,
            I => \N__19897\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__19900\,
            I => \N__19894\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__19897\,
            I => data_out_7_6
        );

    \I__4536\ : Odrv4
    port map (
            O => \N__19894\,
            I => data_out_7_6
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__19889\,
            I => \c0.n4879_cascade_\
        );

    \I__4534\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19882\
        );

    \I__4533\ : InMux
    port map (
            O => \N__19885\,
            I => \N__19879\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__19882\,
            I => \N__19873\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__19879\,
            I => \N__19870\
        );

    \I__4530\ : InMux
    port map (
            O => \N__19878\,
            I => \N__19867\
        );

    \I__4529\ : InMux
    port map (
            O => \N__19877\,
            I => \N__19864\
        );

    \I__4528\ : InMux
    port map (
            O => \N__19876\,
            I => \N__19861\
        );

    \I__4527\ : Span4Mux_s3_v
    port map (
            O => \N__19873\,
            I => \N__19854\
        );

    \I__4526\ : Span4Mux_h
    port map (
            O => \N__19870\,
            I => \N__19854\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__19867\,
            I => \N__19854\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__19864\,
            I => \c0.data_out_field_47_N_682_46\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__19861\,
            I => \c0.data_out_field_47_N_682_46\
        );

    \I__4522\ : Odrv4
    port map (
            O => \N__19854\,
            I => \c0.data_out_field_47_N_682_46\
        );

    \I__4521\ : InMux
    port map (
            O => \N__19847\,
            I => \N__19844\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__19844\,
            I => \N__19841\
        );

    \I__4519\ : Span4Mux_h
    port map (
            O => \N__19841\,
            I => \N__19838\
        );

    \I__4518\ : Span4Mux_h
    port map (
            O => \N__19838\,
            I => \N__19834\
        );

    \I__4517\ : InMux
    port map (
            O => \N__19837\,
            I => \N__19831\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__19834\,
            I => \c0.tx_transmit_N_274_7\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__19831\,
            I => \c0.tx_transmit_N_274_7\
        );

    \I__4514\ : InMux
    port map (
            O => \N__19826\,
            I => \N__19823\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__19823\,
            I => \N__19818\
        );

    \I__4512\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19814\
        );

    \I__4511\ : InMux
    port map (
            O => \N__19821\,
            I => \N__19810\
        );

    \I__4510\ : Span4Mux_h
    port map (
            O => \N__19818\,
            I => \N__19807\
        );

    \I__4509\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19804\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__19814\,
            I => \N__19801\
        );

    \I__4507\ : InMux
    port map (
            O => \N__19813\,
            I => \N__19798\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__19810\,
            I => \c0.data_out_field_47_N_682_35\
        );

    \I__4505\ : Odrv4
    port map (
            O => \N__19807\,
            I => \c0.data_out_field_47_N_682_35\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__19804\,
            I => \c0.data_out_field_47_N_682_35\
        );

    \I__4503\ : Odrv12
    port map (
            O => \N__19801\,
            I => \c0.data_out_field_47_N_682_35\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__19798\,
            I => \c0.data_out_field_47_N_682_35\
        );

    \I__4501\ : InMux
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__4499\ : Span4Mux_h
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__4498\ : Odrv4
    port map (
            O => \N__19778\,
            I => n10_adj_947
        );

    \I__4497\ : CascadeMux
    port map (
            O => \N__19775\,
            I => \n9_adj_948_cascade_\
        );

    \I__4496\ : InMux
    port map (
            O => \N__19772\,
            I => \N__19769\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__19769\,
            I => \N__19764\
        );

    \I__4494\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19759\
        );

    \I__4493\ : InMux
    port map (
            O => \N__19767\,
            I => \N__19759\
        );

    \I__4492\ : Span4Mux_h
    port map (
            O => \N__19764\,
            I => \N__19755\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__19759\,
            I => \N__19752\
        );

    \I__4490\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19749\
        );

    \I__4489\ : Span4Mux_h
    port map (
            O => \N__19755\,
            I => \N__19746\
        );

    \I__4488\ : Span4Mux_v
    port map (
            O => \N__19752\,
            I => \N__19743\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__19749\,
            I => data_out_field_27
        );

    \I__4486\ : Odrv4
    port map (
            O => \N__19746\,
            I => data_out_field_27
        );

    \I__4485\ : Odrv4
    port map (
            O => \N__19743\,
            I => data_out_field_27
        );

    \I__4484\ : CascadeMux
    port map (
            O => \N__19736\,
            I => \N__19733\
        );

    \I__4483\ : InMux
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__4481\ : Span12Mux_h
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__4480\ : Odrv12
    port map (
            O => \N__19724\,
            I => n4_adj_942
        );

    \I__4479\ : CascadeMux
    port map (
            O => \N__19721\,
            I => \N__19718\
        );

    \I__4478\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__4476\ : Span4Mux_v
    port map (
            O => \N__19712\,
            I => \N__19709\
        );

    \I__4475\ : Odrv4
    port map (
            O => \N__19709\,
            I => \c0.n4531\
        );

    \I__4474\ : InMux
    port map (
            O => \N__19706\,
            I => \N__19703\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__19703\,
            I => \N__19700\
        );

    \I__4472\ : Odrv4
    port map (
            O => \N__19700\,
            I => n8_adj_968
        );

    \I__4471\ : InMux
    port map (
            O => \N__19697\,
            I => \N__19693\
        );

    \I__4470\ : InMux
    port map (
            O => \N__19696\,
            I => \N__19690\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__19693\,
            I => data_out_7_0
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__19690\,
            I => data_out_7_0
        );

    \I__4467\ : InMux
    port map (
            O => \N__19685\,
            I => \N__19679\
        );

    \I__4466\ : InMux
    port map (
            O => \N__19684\,
            I => \N__19679\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__19679\,
            I => data_out_6_0
        );

    \I__4464\ : CascadeMux
    port map (
            O => \N__19676\,
            I => \N__19673\
        );

    \I__4463\ : InMux
    port map (
            O => \N__19673\,
            I => \N__19670\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__19670\,
            I => \N__19667\
        );

    \I__4461\ : Odrv12
    port map (
            O => \N__19667\,
            I => \c0.n4577\
        );

    \I__4460\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19661\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__4458\ : Span4Mux_h
    port map (
            O => \N__19658\,
            I => \N__19652\
        );

    \I__4457\ : InMux
    port map (
            O => \N__19657\,
            I => \N__19649\
        );

    \I__4456\ : InMux
    port map (
            O => \N__19656\,
            I => \N__19644\
        );

    \I__4455\ : InMux
    port map (
            O => \N__19655\,
            I => \N__19644\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__19652\,
            I => data_out_field_6
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__19649\,
            I => data_out_field_6
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__19644\,
            I => data_out_field_6
        );

    \I__4451\ : CascadeMux
    port map (
            O => \N__19637\,
            I => \n1246_cascade_\
        );

    \I__4450\ : CascadeMux
    port map (
            O => \N__19634\,
            I => \N__19629\
        );

    \I__4449\ : InMux
    port map (
            O => \N__19633\,
            I => \N__19625\
        );

    \I__4448\ : InMux
    port map (
            O => \N__19632\,
            I => \N__19622\
        );

    \I__4447\ : InMux
    port map (
            O => \N__19629\,
            I => \N__19619\
        );

    \I__4446\ : InMux
    port map (
            O => \N__19628\,
            I => \N__19616\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__19625\,
            I => data_out_field_22
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__19622\,
            I => data_out_field_22
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__19619\,
            I => data_out_field_22
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__19616\,
            I => data_out_field_22
        );

    \I__4441\ : InMux
    port map (
            O => \N__19607\,
            I => \c0.n3844\
        );

    \I__4440\ : CascadeMux
    port map (
            O => \N__19604\,
            I => \N__19598\
        );

    \I__4439\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19591\
        );

    \I__4438\ : InMux
    port map (
            O => \N__19602\,
            I => \N__19591\
        );

    \I__4437\ : InMux
    port map (
            O => \N__19601\,
            I => \N__19586\
        );

    \I__4436\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19582\
        );

    \I__4435\ : InMux
    port map (
            O => \N__19597\,
            I => \N__19577\
        );

    \I__4434\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19577\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__19591\,
            I => \N__19574\
        );

    \I__4432\ : InMux
    port map (
            O => \N__19590\,
            I => \N__19569\
        );

    \I__4431\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19569\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__19586\,
            I => \N__19562\
        );

    \I__4429\ : InMux
    port map (
            O => \N__19585\,
            I => \N__19558\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__19582\,
            I => \N__19549\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__19577\,
            I => \N__19549\
        );

    \I__4426\ : Span4Mux_v
    port map (
            O => \N__19574\,
            I => \N__19549\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__19569\,
            I => \N__19549\
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__19568\,
            I => \N__19546\
        );

    \I__4423\ : InMux
    port map (
            O => \N__19567\,
            I => \N__19541\
        );

    \I__4422\ : InMux
    port map (
            O => \N__19566\,
            I => \N__19541\
        );

    \I__4421\ : InMux
    port map (
            O => \N__19565\,
            I => \N__19538\
        );

    \I__4420\ : Span4Mux_v
    port map (
            O => \N__19562\,
            I => \N__19535\
        );

    \I__4419\ : InMux
    port map (
            O => \N__19561\,
            I => \N__19532\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__19558\,
            I => \N__19529\
        );

    \I__4417\ : Span4Mux_v
    port map (
            O => \N__19549\,
            I => \N__19526\
        );

    \I__4416\ : InMux
    port map (
            O => \N__19546\,
            I => \N__19523\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__19541\,
            I => \N__19517\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__19538\,
            I => \N__19517\
        );

    \I__4413\ : Span4Mux_h
    port map (
            O => \N__19535\,
            I => \N__19512\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__19532\,
            I => \N__19512\
        );

    \I__4411\ : Span4Mux_h
    port map (
            O => \N__19529\,
            I => \N__19505\
        );

    \I__4410\ : Span4Mux_h
    port map (
            O => \N__19526\,
            I => \N__19505\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__19523\,
            I => \N__19505\
        );

    \I__4408\ : InMux
    port map (
            O => \N__19522\,
            I => \N__19502\
        );

    \I__4407\ : Odrv12
    port map (
            O => \N__19517\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__4406\ : Odrv4
    port map (
            O => \N__19512\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__4405\ : Odrv4
    port map (
            O => \N__19505\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__19502\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__4403\ : InMux
    port map (
            O => \N__19493\,
            I => \c0.n3845\
        );

    \I__4402\ : InMux
    port map (
            O => \N__19490\,
            I => \N__19487\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__19487\,
            I => \c0.byte_transmit_counter_3\
        );

    \I__4400\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19480\
        );

    \I__4399\ : InMux
    port map (
            O => \N__19483\,
            I => \N__19477\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__19480\,
            I => \c0.tx_transmit_N_274_3\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__19477\,
            I => \c0.tx_transmit_N_274_3\
        );

    \I__4396\ : InMux
    port map (
            O => \N__19472\,
            I => \c0.n3846\
        );

    \I__4395\ : InMux
    port map (
            O => \N__19469\,
            I => \N__19466\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__19466\,
            I => \N__19463\
        );

    \I__4393\ : Span12Mux_s7_v
    port map (
            O => \N__19463\,
            I => \N__19460\
        );

    \I__4392\ : Odrv12
    port map (
            O => \N__19460\,
            I => \c0.byte_transmit_counter_4\
        );

    \I__4391\ : InMux
    port map (
            O => \N__19457\,
            I => \N__19454\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__19454\,
            I => \N__19451\
        );

    \I__4389\ : Span4Mux_h
    port map (
            O => \N__19451\,
            I => \N__19448\
        );

    \I__4388\ : Span4Mux_h
    port map (
            O => \N__19448\,
            I => \N__19444\
        );

    \I__4387\ : InMux
    port map (
            O => \N__19447\,
            I => \N__19441\
        );

    \I__4386\ : Odrv4
    port map (
            O => \N__19444\,
            I => \c0.tx_transmit_N_274_4\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__19441\,
            I => \c0.tx_transmit_N_274_4\
        );

    \I__4384\ : InMux
    port map (
            O => \N__19436\,
            I => \c0.n3847\
        );

    \I__4383\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19430\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__19430\,
            I => \N__19427\
        );

    \I__4381\ : Span4Mux_h
    port map (
            O => \N__19427\,
            I => \N__19424\
        );

    \I__4380\ : Span4Mux_h
    port map (
            O => \N__19424\,
            I => \N__19421\
        );

    \I__4379\ : Odrv4
    port map (
            O => \N__19421\,
            I => \c0.byte_transmit_counter_5\
        );

    \I__4378\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19415\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__19415\,
            I => \N__19412\
        );

    \I__4376\ : Span4Mux_h
    port map (
            O => \N__19412\,
            I => \N__19409\
        );

    \I__4375\ : Span4Mux_h
    port map (
            O => \N__19409\,
            I => \N__19405\
        );

    \I__4374\ : InMux
    port map (
            O => \N__19408\,
            I => \N__19402\
        );

    \I__4373\ : Odrv4
    port map (
            O => \N__19405\,
            I => \c0.tx_transmit_N_274_5\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__19402\,
            I => \c0.tx_transmit_N_274_5\
        );

    \I__4371\ : InMux
    port map (
            O => \N__19397\,
            I => \c0.n3848\
        );

    \I__4370\ : InMux
    port map (
            O => \N__19394\,
            I => \N__19391\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__19391\,
            I => \N__19388\
        );

    \I__4368\ : Span4Mux_h
    port map (
            O => \N__19388\,
            I => \N__19385\
        );

    \I__4367\ : Span4Mux_h
    port map (
            O => \N__19385\,
            I => \N__19382\
        );

    \I__4366\ : Odrv4
    port map (
            O => \N__19382\,
            I => \c0.byte_transmit_counter_6\
        );

    \I__4365\ : InMux
    port map (
            O => \N__19379\,
            I => \N__19376\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__19376\,
            I => \N__19373\
        );

    \I__4363\ : Span4Mux_h
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__4362\ : Span4Mux_h
    port map (
            O => \N__19370\,
            I => \N__19366\
        );

    \I__4361\ : InMux
    port map (
            O => \N__19369\,
            I => \N__19363\
        );

    \I__4360\ : Odrv4
    port map (
            O => \N__19366\,
            I => \c0.tx_transmit_N_274_6\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__19363\,
            I => \c0.tx_transmit_N_274_6\
        );

    \I__4358\ : InMux
    port map (
            O => \N__19358\,
            I => \c0.n3849\
        );

    \I__4357\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19352\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__4355\ : Span4Mux_v
    port map (
            O => \N__19349\,
            I => \N__19346\
        );

    \I__4354\ : Span4Mux_h
    port map (
            O => \N__19346\,
            I => \N__19343\
        );

    \I__4353\ : Odrv4
    port map (
            O => \N__19343\,
            I => \c0.byte_transmit_counter_7\
        );

    \I__4352\ : InMux
    port map (
            O => \N__19340\,
            I => \c0.n3850\
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__19337\,
            I => \c0.n4774_cascade_\
        );

    \I__4350\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19331\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__19331\,
            I => \N__19328\
        );

    \I__4348\ : Span4Mux_v
    port map (
            O => \N__19328\,
            I => \N__19325\
        );

    \I__4347\ : Odrv4
    port map (
            O => \N__19325\,
            I => tx_data_6_keep
        );

    \I__4346\ : CascadeMux
    port map (
            O => \N__19322\,
            I => \N__19319\
        );

    \I__4345\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19316\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__19316\,
            I => \N__19313\
        );

    \I__4343\ : Span4Mux_h
    port map (
            O => \N__19313\,
            I => \N__19310\
        );

    \I__4342\ : Odrv4
    port map (
            O => \N__19310\,
            I => n10_adj_971
        );

    \I__4341\ : CascadeMux
    port map (
            O => \N__19307\,
            I => \N__19304\
        );

    \I__4340\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19301\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__19301\,
            I => \N__19298\
        );

    \I__4338\ : Span4Mux_h
    port map (
            O => \N__19298\,
            I => \N__19294\
        );

    \I__4337\ : InMux
    port map (
            O => \N__19297\,
            I => \N__19291\
        );

    \I__4336\ : Odrv4
    port map (
            O => \N__19294\,
            I => \c0.data_12\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__19291\,
            I => \c0.data_12\
        );

    \I__4334\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19282\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__19285\,
            I => \N__19278\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__19282\,
            I => \N__19275\
        );

    \I__4331\ : InMux
    port map (
            O => \N__19281\,
            I => \N__19270\
        );

    \I__4330\ : InMux
    port map (
            O => \N__19278\,
            I => \N__19270\
        );

    \I__4329\ : Odrv12
    port map (
            O => \N__19275\,
            I => data_out_field_7
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__19270\,
            I => data_out_field_7
        );

    \I__4327\ : InMux
    port map (
            O => \N__19265\,
            I => \N__19262\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__19262\,
            I => \N__19258\
        );

    \I__4325\ : CascadeMux
    port map (
            O => \N__19261\,
            I => \N__19253\
        );

    \I__4324\ : Span4Mux_h
    port map (
            O => \N__19258\,
            I => \N__19250\
        );

    \I__4323\ : InMux
    port map (
            O => \N__19257\,
            I => \N__19247\
        );

    \I__4322\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19242\
        );

    \I__4321\ : InMux
    port map (
            O => \N__19253\,
            I => \N__19242\
        );

    \I__4320\ : Odrv4
    port map (
            O => \N__19250\,
            I => \c0.tx.r_Bit_Index_2\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__19247\,
            I => \c0.tx.r_Bit_Index_2\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__19242\,
            I => \c0.tx.r_Bit_Index_2\
        );

    \I__4317\ : InMux
    port map (
            O => \N__19235\,
            I => \N__19232\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__19232\,
            I => \N__19229\
        );

    \I__4315\ : Span12Mux_s3_v
    port map (
            O => \N__19229\,
            I => \N__19223\
        );

    \I__4314\ : InMux
    port map (
            O => \N__19228\,
            I => \N__19216\
        );

    \I__4313\ : InMux
    port map (
            O => \N__19227\,
            I => \N__19216\
        );

    \I__4312\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19216\
        );

    \I__4311\ : Odrv12
    port map (
            O => \N__19223\,
            I => \c0.tx.r_Bit_Index_1\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__19216\,
            I => \c0.tx.r_Bit_Index_1\
        );

    \I__4309\ : InMux
    port map (
            O => \N__19211\,
            I => \N__19203\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__19210\,
            I => \N__19200\
        );

    \I__4307\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19194\
        );

    \I__4306\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19194\
        );

    \I__4305\ : InMux
    port map (
            O => \N__19207\,
            I => \N__19189\
        );

    \I__4304\ : InMux
    port map (
            O => \N__19206\,
            I => \N__19189\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__19203\,
            I => \N__19186\
        );

    \I__4302\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19182\
        );

    \I__4301\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19179\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__19194\,
            I => \N__19172\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__19189\,
            I => \N__19172\
        );

    \I__4298\ : Span4Mux_h
    port map (
            O => \N__19186\,
            I => \N__19172\
        );

    \I__4297\ : InMux
    port map (
            O => \N__19185\,
            I => \N__19169\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__19182\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__19179\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__4294\ : Odrv4
    port map (
            O => \N__19172\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__19169\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__4292\ : InMux
    port map (
            O => \N__19160\,
            I => \N__19156\
        );

    \I__4291\ : InMux
    port map (
            O => \N__19159\,
            I => \N__19153\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__19156\,
            I => data_out_6_5
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__19153\,
            I => data_out_6_5
        );

    \I__4288\ : InMux
    port map (
            O => \N__19148\,
            I => \N__19145\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__19145\,
            I => \c0.n4616\
        );

    \I__4286\ : InMux
    port map (
            O => \N__19142\,
            I => \N__19136\
        );

    \I__4285\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19133\
        );

    \I__4284\ : InMux
    port map (
            O => \N__19140\,
            I => \N__19127\
        );

    \I__4283\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19127\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__19136\,
            I => \N__19122\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__19133\,
            I => \N__19122\
        );

    \I__4280\ : InMux
    port map (
            O => \N__19132\,
            I => \N__19119\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__19127\,
            I => data_out_field_25
        );

    \I__4278\ : Odrv12
    port map (
            O => \N__19122\,
            I => data_out_field_25
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__19119\,
            I => data_out_field_25
        );

    \I__4276\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19107\
        );

    \I__4275\ : InMux
    port map (
            O => \N__19111\,
            I => \N__19102\
        );

    \I__4274\ : InMux
    port map (
            O => \N__19110\,
            I => \N__19099\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__19107\,
            I => \N__19096\
        );

    \I__4272\ : InMux
    port map (
            O => \N__19106\,
            I => \N__19091\
        );

    \I__4271\ : InMux
    port map (
            O => \N__19105\,
            I => \N__19091\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__19102\,
            I => \c0.data_out_field_47_N_682_40\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__19099\,
            I => \c0.data_out_field_47_N_682_40\
        );

    \I__4268\ : Odrv4
    port map (
            O => \N__19096\,
            I => \c0.data_out_field_47_N_682_40\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__19091\,
            I => \c0.data_out_field_47_N_682_40\
        );

    \I__4266\ : InMux
    port map (
            O => \N__19082\,
            I => \N__19079\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__19079\,
            I => \N__19076\
        );

    \I__4264\ : Span4Mux_v
    port map (
            O => \N__19076\,
            I => \N__19073\
        );

    \I__4263\ : Span4Mux_h
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__19070\,
            I => \c0.n4561\
        );

    \I__4261\ : CascadeMux
    port map (
            O => \N__19067\,
            I => \N__19064\
        );

    \I__4260\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__19061\,
            I => \N__19057\
        );

    \I__4258\ : InMux
    port map (
            O => \N__19060\,
            I => \N__19054\
        );

    \I__4257\ : Odrv12
    port map (
            O => \N__19057\,
            I => \c0.data_2\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__19054\,
            I => \c0.data_2\
        );

    \I__4255\ : CascadeMux
    port map (
            O => \N__19049\,
            I => \c0.n4771_cascade_\
        );

    \I__4254\ : InMux
    port map (
            O => \N__19046\,
            I => \N__19043\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__19043\,
            I => n7_adj_935
        );

    \I__4252\ : CascadeMux
    port map (
            O => \N__19040\,
            I => \n8_adj_934_cascade_\
        );

    \I__4251\ : CascadeMux
    port map (
            O => \N__19037\,
            I => \N__19034\
        );

    \I__4250\ : InMux
    port map (
            O => \N__19034\,
            I => \N__19030\
        );

    \I__4249\ : InMux
    port map (
            O => \N__19033\,
            I => \N__19027\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__19030\,
            I => \N__19024\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__19027\,
            I => data_out_7_7
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__19024\,
            I => data_out_7_7
        );

    \I__4245\ : InMux
    port map (
            O => \N__19019\,
            I => \N__19016\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__19016\,
            I => \N__19013\
        );

    \I__4243\ : Span4Mux_h
    port map (
            O => \N__19013\,
            I => \N__19010\
        );

    \I__4242\ : Odrv4
    port map (
            O => \N__19010\,
            I => \c0.n1333\
        );

    \I__4241\ : CascadeMux
    port map (
            O => \N__19007\,
            I => \c0.n4447_cascade_\
        );

    \I__4240\ : InMux
    port map (
            O => \N__19004\,
            I => \N__19001\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__19001\,
            I => n9_adj_972
        );

    \I__4238\ : InMux
    port map (
            O => \N__18998\,
            I => \N__18995\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__18995\,
            I => \N__18992\
        );

    \I__4236\ : Odrv4
    port map (
            O => \N__18992\,
            I => \c0.n4795\
        );

    \I__4235\ : InMux
    port map (
            O => \N__18989\,
            I => \N__18986\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__18986\,
            I => \N__18983\
        );

    \I__4233\ : Odrv4
    port map (
            O => \N__18983\,
            I => n11_adj_945
        );

    \I__4232\ : InMux
    port map (
            O => \N__18980\,
            I => \N__18977\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__18977\,
            I => \N__18974\
        );

    \I__4230\ : Span4Mux_v
    port map (
            O => \N__18974\,
            I => \N__18971\
        );

    \I__4229\ : Odrv4
    port map (
            O => \N__18971\,
            I => n4_adj_970
        );

    \I__4228\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18961\
        );

    \I__4227\ : InMux
    port map (
            O => \N__18967\,
            I => \N__18958\
        );

    \I__4226\ : InMux
    port map (
            O => \N__18966\,
            I => \N__18955\
        );

    \I__4225\ : InMux
    port map (
            O => \N__18965\,
            I => \N__18952\
        );

    \I__4224\ : InMux
    port map (
            O => \N__18964\,
            I => \N__18949\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__18961\,
            I => \N__18946\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__18958\,
            I => data_out_field_16
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__18955\,
            I => data_out_field_16
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__18952\,
            I => data_out_field_16
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__18949\,
            I => data_out_field_16
        );

    \I__4218\ : Odrv4
    port map (
            O => \N__18946\,
            I => data_out_field_16
        );

    \I__4217\ : InMux
    port map (
            O => \N__18935\,
            I => \N__18932\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__18932\,
            I => \c0.n4447\
        );

    \I__4215\ : CascadeMux
    port map (
            O => \N__18929\,
            I => \n7_adj_969_cascade_\
        );

    \I__4214\ : InMux
    port map (
            O => \N__18926\,
            I => \N__18922\
        );

    \I__4213\ : InMux
    port map (
            O => \N__18925\,
            I => \N__18919\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__18922\,
            I => \N__18916\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__18919\,
            I => \N__18913\
        );

    \I__4210\ : Span4Mux_h
    port map (
            O => \N__18916\,
            I => \N__18910\
        );

    \I__4209\ : Odrv12
    port map (
            O => \N__18913\,
            I => \c0.n4380\
        );

    \I__4208\ : Odrv4
    port map (
            O => \N__18910\,
            I => \c0.n4380\
        );

    \I__4207\ : InMux
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__18902\,
            I => \N__18898\
        );

    \I__4205\ : InMux
    port map (
            O => \N__18901\,
            I => \N__18895\
        );

    \I__4204\ : Span4Mux_v
    port map (
            O => \N__18898\,
            I => \N__18889\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__18895\,
            I => \N__18889\
        );

    \I__4202\ : InMux
    port map (
            O => \N__18894\,
            I => \N__18884\
        );

    \I__4201\ : Span4Mux_h
    port map (
            O => \N__18889\,
            I => \N__18881\
        );

    \I__4200\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18878\
        );

    \I__4199\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18875\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__18884\,
            I => \c0.data_out_field_47_N_682_33\
        );

    \I__4197\ : Odrv4
    port map (
            O => \N__18881\,
            I => \c0.data_out_field_47_N_682_33\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__18878\,
            I => \c0.data_out_field_47_N_682_33\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__18875\,
            I => \c0.data_out_field_47_N_682_33\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__18866\,
            I => \N__18863\
        );

    \I__4193\ : InMux
    port map (
            O => \N__18863\,
            I => \N__18860\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__18860\,
            I => \c0.n4393\
        );

    \I__4191\ : InMux
    port map (
            O => \N__18857\,
            I => \N__18854\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__18854\,
            I => \N__18851\
        );

    \I__4189\ : Odrv4
    port map (
            O => \N__18851\,
            I => n12_adj_966
        );

    \I__4188\ : CascadeMux
    port map (
            O => \N__18848\,
            I => \n1677_cascade_\
        );

    \I__4187\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18841\
        );

    \I__4186\ : InMux
    port map (
            O => \N__18844\,
            I => \N__18838\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__18841\,
            I => \N__18835\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__18838\,
            I => data_out_6_7
        );

    \I__4183\ : Odrv4
    port map (
            O => \N__18835\,
            I => data_out_6_7
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__4181\ : InMux
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__18824\,
            I => \c0.n4885\
        );

    \I__4179\ : InMux
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__4177\ : Span4Mux_h
    port map (
            O => \N__18815\,
            I => \N__18811\
        );

    \I__4176\ : InMux
    port map (
            O => \N__18814\,
            I => \N__18808\
        );

    \I__4175\ : Odrv4
    port map (
            O => \N__18811\,
            I => \c0.data_5\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__18808\,
            I => \c0.data_5\
        );

    \I__4173\ : CascadeMux
    port map (
            O => \N__18803\,
            I => \c0.n6_adj_904_cascade_\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__18800\,
            I => \n7_adj_938_cascade_\
        );

    \I__4171\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__18794\,
            I => \N__18790\
        );

    \I__4169\ : InMux
    port map (
            O => \N__18793\,
            I => \N__18787\
        );

    \I__4168\ : Span4Mux_v
    port map (
            O => \N__18790\,
            I => \N__18782\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__18787\,
            I => \N__18782\
        );

    \I__4166\ : Span4Mux_h
    port map (
            O => \N__18782\,
            I => \N__18779\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__18779\,
            I => data_out_6_3
        );

    \I__4164\ : InMux
    port map (
            O => \N__18776\,
            I => \N__18772\
        );

    \I__4163\ : InMux
    port map (
            O => \N__18775\,
            I => \N__18769\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__18772\,
            I => \c0.delay_counter_6\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__18769\,
            I => \c0.delay_counter_6\
        );

    \I__4160\ : CascadeMux
    port map (
            O => \N__18764\,
            I => \N__18761\
        );

    \I__4159\ : InMux
    port map (
            O => \N__18761\,
            I => \N__18757\
        );

    \I__4158\ : InMux
    port map (
            O => \N__18760\,
            I => \N__18754\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__18757\,
            I => \c0.delay_counter_0\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__18754\,
            I => \c0.delay_counter_0\
        );

    \I__4155\ : CascadeMux
    port map (
            O => \N__18749\,
            I => \N__18745\
        );

    \I__4154\ : InMux
    port map (
            O => \N__18748\,
            I => \N__18742\
        );

    \I__4153\ : InMux
    port map (
            O => \N__18745\,
            I => \N__18739\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__18742\,
            I => \c0.delay_counter_2\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__18739\,
            I => \c0.delay_counter_2\
        );

    \I__4150\ : InMux
    port map (
            O => \N__18734\,
            I => \N__18730\
        );

    \I__4149\ : InMux
    port map (
            O => \N__18733\,
            I => \N__18727\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__18730\,
            I => \c0.delay_counter_4\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__18727\,
            I => \c0.delay_counter_4\
        );

    \I__4146\ : InMux
    port map (
            O => \N__18722\,
            I => \N__18718\
        );

    \I__4145\ : InMux
    port map (
            O => \N__18721\,
            I => \N__18715\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__18718\,
            I => \c0.delay_counter_5\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__18715\,
            I => \c0.delay_counter_5\
        );

    \I__4142\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18706\
        );

    \I__4141\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18703\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__18706\,
            I => \c0.delay_counter_1\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__18703\,
            I => \c0.delay_counter_1\
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__18698\,
            I => \N__18694\
        );

    \I__4137\ : InMux
    port map (
            O => \N__18697\,
            I => \N__18691\
        );

    \I__4136\ : InMux
    port map (
            O => \N__18694\,
            I => \N__18688\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__18691\,
            I => \c0.delay_counter_7\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__18688\,
            I => \c0.delay_counter_7\
        );

    \I__4133\ : InMux
    port map (
            O => \N__18683\,
            I => \N__18679\
        );

    \I__4132\ : InMux
    port map (
            O => \N__18682\,
            I => \N__18676\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__18679\,
            I => \c0.delay_counter_3\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__18676\,
            I => \c0.delay_counter_3\
        );

    \I__4129\ : InMux
    port map (
            O => \N__18671\,
            I => \N__18668\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__18668\,
            I => \c0.n13\
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__18665\,
            I => \c0.n14_adj_902_cascade_\
        );

    \I__4126\ : InMux
    port map (
            O => \N__18662\,
            I => \N__18659\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__18659\,
            I => \N__18655\
        );

    \I__4124\ : InMux
    port map (
            O => \N__18658\,
            I => \N__18652\
        );

    \I__4123\ : Odrv12
    port map (
            O => \N__18655\,
            I => \c0.data_4\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__18652\,
            I => \c0.data_4\
        );

    \I__4121\ : CascadeMux
    port map (
            O => \N__18647\,
            I => \n3580_cascade_\
        );

    \I__4120\ : CascadeMux
    port map (
            O => \N__18644\,
            I => \N__18641\
        );

    \I__4119\ : InMux
    port map (
            O => \N__18641\,
            I => \N__18638\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__18638\,
            I => \N__18635\
        );

    \I__4117\ : Span4Mux_h
    port map (
            O => \N__18635\,
            I => \N__18631\
        );

    \I__4116\ : InMux
    port map (
            O => \N__18634\,
            I => \N__18628\
        );

    \I__4115\ : Odrv4
    port map (
            O => \N__18631\,
            I => \c0.data_11\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__18628\,
            I => \c0.data_11\
        );

    \I__4113\ : CascadeMux
    port map (
            O => \N__18623\,
            I => \N__18620\
        );

    \I__4112\ : InMux
    port map (
            O => \N__18620\,
            I => \N__18617\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__18617\,
            I => \N__18614\
        );

    \I__4110\ : Span4Mux_h
    port map (
            O => \N__18614\,
            I => \N__18610\
        );

    \I__4109\ : InMux
    port map (
            O => \N__18613\,
            I => \N__18607\
        );

    \I__4108\ : Odrv4
    port map (
            O => \N__18610\,
            I => \c0.data_3\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__18607\,
            I => \c0.data_3\
        );

    \I__4106\ : InMux
    port map (
            O => \N__18602\,
            I => \N__18599\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__18599\,
            I => n7_adj_933
        );

    \I__4104\ : InMux
    port map (
            O => \N__18596\,
            I => \N__18593\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__18593\,
            I => \N__18589\
        );

    \I__4102\ : InMux
    port map (
            O => \N__18592\,
            I => \N__18586\
        );

    \I__4101\ : Span4Mux_s3_v
    port map (
            O => \N__18589\,
            I => \N__18579\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__18586\,
            I => \N__18579\
        );

    \I__4099\ : InMux
    port map (
            O => \N__18585\,
            I => \N__18576\
        );

    \I__4098\ : InMux
    port map (
            O => \N__18584\,
            I => \N__18573\
        );

    \I__4097\ : Span4Mux_h
    port map (
            O => \N__18579\,
            I => \N__18570\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__18576\,
            I => \c0.data_out_field_47_N_682_41\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__18573\,
            I => \c0.data_out_field_47_N_682_41\
        );

    \I__4094\ : Odrv4
    port map (
            O => \N__18570\,
            I => \c0.data_out_field_47_N_682_41\
        );

    \I__4093\ : InMux
    port map (
            O => \N__18563\,
            I => \N__18559\
        );

    \I__4092\ : InMux
    port map (
            O => \N__18562\,
            I => \N__18553\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__18559\,
            I => \N__18550\
        );

    \I__4090\ : InMux
    port map (
            O => \N__18558\,
            I => \N__18547\
        );

    \I__4089\ : CascadeMux
    port map (
            O => \N__18557\,
            I => \N__18544\
        );

    \I__4088\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18541\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__18553\,
            I => \N__18538\
        );

    \I__4086\ : Span4Mux_v
    port map (
            O => \N__18550\,
            I => \N__18533\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__18547\,
            I => \N__18533\
        );

    \I__4084\ : InMux
    port map (
            O => \N__18544\,
            I => \N__18530\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__18541\,
            I => \N__18523\
        );

    \I__4082\ : Span4Mux_h
    port map (
            O => \N__18538\,
            I => \N__18523\
        );

    \I__4081\ : Span4Mux_h
    port map (
            O => \N__18533\,
            I => \N__18523\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__18530\,
            I => \c0.data_out_field_47_N_682_34\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__18523\,
            I => \c0.data_out_field_47_N_682_34\
        );

    \I__4078\ : CascadeMux
    port map (
            O => \N__18518\,
            I => \c0.n1384_cascade_\
        );

    \I__4077\ : InMux
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__18512\,
            I => \N__18505\
        );

    \I__4075\ : InMux
    port map (
            O => \N__18511\,
            I => \N__18502\
        );

    \I__4074\ : InMux
    port map (
            O => \N__18510\,
            I => \N__18497\
        );

    \I__4073\ : InMux
    port map (
            O => \N__18509\,
            I => \N__18497\
        );

    \I__4072\ : InMux
    port map (
            O => \N__18508\,
            I => \N__18494\
        );

    \I__4071\ : Span4Mux_v
    port map (
            O => \N__18505\,
            I => \N__18491\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__18502\,
            I => \N__18486\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__18497\,
            I => \N__18486\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__18494\,
            I => \c0.data_out_field_47_N_682_32\
        );

    \I__4067\ : Odrv4
    port map (
            O => \N__18491\,
            I => \c0.data_out_field_47_N_682_32\
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__18486\,
            I => \c0.data_out_field_47_N_682_32\
        );

    \I__4065\ : InMux
    port map (
            O => \N__18479\,
            I => \N__18476\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__18476\,
            I => \N__18472\
        );

    \I__4063\ : InMux
    port map (
            O => \N__18475\,
            I => \N__18467\
        );

    \I__4062\ : Span4Mux_h
    port map (
            O => \N__18472\,
            I => \N__18464\
        );

    \I__4061\ : InMux
    port map (
            O => \N__18471\,
            I => \N__18459\
        );

    \I__4060\ : InMux
    port map (
            O => \N__18470\,
            I => \N__18459\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__18467\,
            I => data_out_field_3
        );

    \I__4058\ : Odrv4
    port map (
            O => \N__18464\,
            I => data_out_field_3
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__18459\,
            I => data_out_field_3
        );

    \I__4056\ : InMux
    port map (
            O => \N__18452\,
            I => \N__18447\
        );

    \I__4055\ : CascadeMux
    port map (
            O => \N__18451\,
            I => \N__18443\
        );

    \I__4054\ : InMux
    port map (
            O => \N__18450\,
            I => \N__18440\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__18447\,
            I => \N__18437\
        );

    \I__4052\ : InMux
    port map (
            O => \N__18446\,
            I => \N__18432\
        );

    \I__4051\ : InMux
    port map (
            O => \N__18443\,
            I => \N__18432\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__18440\,
            I => \N__18427\
        );

    \I__4049\ : Span4Mux_v
    port map (
            O => \N__18437\,
            I => \N__18427\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__18432\,
            I => \N__18424\
        );

    \I__4047\ : Odrv4
    port map (
            O => \N__18427\,
            I => data_out_field_4
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__18424\,
            I => data_out_field_4
        );

    \I__4045\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18416\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__18416\,
            I => \N__18413\
        );

    \I__4043\ : Span4Mux_h
    port map (
            O => \N__18413\,
            I => \N__18410\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__18410\,
            I => \c0.n4529\
        );

    \I__4041\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18404\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__4039\ : Span4Mux_v
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__4038\ : Odrv4
    port map (
            O => \N__18398\,
            I => n7_adj_937
        );

    \I__4037\ : InMux
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__18392\,
            I => \N__18389\
        );

    \I__4035\ : Odrv4
    port map (
            O => \N__18389\,
            I => \c0.n4565\
        );

    \I__4034\ : CascadeMux
    port map (
            O => \N__18386\,
            I => \n11_adj_967_cascade_\
        );

    \I__4033\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18380\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__18380\,
            I => \N__18376\
        );

    \I__4031\ : InMux
    port map (
            O => \N__18379\,
            I => \N__18373\
        );

    \I__4030\ : Span4Mux_v
    port map (
            O => \N__18376\,
            I => \N__18370\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__18373\,
            I => data_out_7_4
        );

    \I__4028\ : Odrv4
    port map (
            O => \N__18370\,
            I => data_out_7_4
        );

    \I__4027\ : InMux
    port map (
            O => \N__18365\,
            I => \N__18361\
        );

    \I__4026\ : InMux
    port map (
            O => \N__18364\,
            I => \N__18358\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__18361\,
            I => \N__18353\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__18358\,
            I => \N__18350\
        );

    \I__4023\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18347\
        );

    \I__4022\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18344\
        );

    \I__4021\ : Span4Mux_h
    port map (
            O => \N__18353\,
            I => \N__18337\
        );

    \I__4020\ : Span4Mux_h
    port map (
            O => \N__18350\,
            I => \N__18337\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__18347\,
            I => \N__18337\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__18344\,
            I => data_out_field_11
        );

    \I__4017\ : Odrv4
    port map (
            O => \N__18337\,
            I => data_out_field_11
        );

    \I__4016\ : CascadeMux
    port map (
            O => \N__18332\,
            I => \c0.n6_cascade_\
        );

    \I__4015\ : InMux
    port map (
            O => \N__18329\,
            I => \N__18324\
        );

    \I__4014\ : InMux
    port map (
            O => \N__18328\,
            I => \N__18321\
        );

    \I__4013\ : InMux
    port map (
            O => \N__18327\,
            I => \N__18318\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__18324\,
            I => \N__18315\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__18321\,
            I => \N__18309\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__18318\,
            I => \N__18309\
        );

    \I__4009\ : Span4Mux_h
    port map (
            O => \N__18315\,
            I => \N__18306\
        );

    \I__4008\ : InMux
    port map (
            O => \N__18314\,
            I => \N__18303\
        );

    \I__4007\ : Span4Mux_v
    port map (
            O => \N__18309\,
            I => \N__18300\
        );

    \I__4006\ : Span4Mux_v
    port map (
            O => \N__18306\,
            I => \N__18297\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__18303\,
            I => data_out_field_24
        );

    \I__4004\ : Odrv4
    port map (
            O => \N__18300\,
            I => data_out_field_24
        );

    \I__4003\ : Odrv4
    port map (
            O => \N__18297\,
            I => data_out_field_24
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__18290\,
            I => \c0.n4456_cascade_\
        );

    \I__4001\ : CascadeMux
    port map (
            O => \N__18287\,
            I => \N__18284\
        );

    \I__4000\ : InMux
    port map (
            O => \N__18284\,
            I => \N__18281\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__18281\,
            I => \N__18278\
        );

    \I__3998\ : Span4Mux_v
    port map (
            O => \N__18278\,
            I => \N__18274\
        );

    \I__3997\ : InMux
    port map (
            O => \N__18277\,
            I => \N__18271\
        );

    \I__3996\ : Odrv4
    port map (
            O => \N__18274\,
            I => \c0.data_0\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__18271\,
            I => \c0.data_0\
        );

    \I__3994\ : InMux
    port map (
            O => \N__18266\,
            I => \N__18262\
        );

    \I__3993\ : InMux
    port map (
            O => \N__18265\,
            I => \N__18258\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__18262\,
            I => \N__18255\
        );

    \I__3991\ : InMux
    port map (
            O => \N__18261\,
            I => \N__18252\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__18258\,
            I => data_out_field_17
        );

    \I__3989\ : Odrv4
    port map (
            O => \N__18255\,
            I => data_out_field_17
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__18252\,
            I => data_out_field_17
        );

    \I__3987\ : InMux
    port map (
            O => \N__18245\,
            I => \N__18242\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__18242\,
            I => \N__18239\
        );

    \I__3985\ : Span4Mux_h
    port map (
            O => \N__18239\,
            I => \N__18236\
        );

    \I__3984\ : Odrv4
    port map (
            O => \N__18236\,
            I => \c0.n4562\
        );

    \I__3983\ : InMux
    port map (
            O => \N__18233\,
            I => \N__18230\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__18230\,
            I => \N__18226\
        );

    \I__3981\ : InMux
    port map (
            O => \N__18229\,
            I => \N__18223\
        );

    \I__3980\ : Span4Mux_v
    port map (
            O => \N__18226\,
            I => \N__18220\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__18223\,
            I => data_out_7_2
        );

    \I__3978\ : Odrv4
    port map (
            O => \N__18220\,
            I => data_out_7_2
        );

    \I__3977\ : InMux
    port map (
            O => \N__18215\,
            I => \N__18211\
        );

    \I__3976\ : InMux
    port map (
            O => \N__18214\,
            I => \N__18208\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__18211\,
            I => \N__18203\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__18208\,
            I => \N__18203\
        );

    \I__3973\ : Odrv12
    port map (
            O => \N__18203\,
            I => data_out_7_1
        );

    \I__3972\ : InMux
    port map (
            O => \N__18200\,
            I => \N__18197\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__18197\,
            I => \N__18194\
        );

    \I__3970\ : Odrv12
    port map (
            O => \N__18194\,
            I => \c0.n4574\
        );

    \I__3969\ : InMux
    port map (
            O => \N__18191\,
            I => \N__18188\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__18188\,
            I => \N__18185\
        );

    \I__3967\ : Span12Mux_h
    port map (
            O => \N__18185\,
            I => \N__18181\
        );

    \I__3966\ : InMux
    port map (
            O => \N__18184\,
            I => \N__18178\
        );

    \I__3965\ : Odrv12
    port map (
            O => \N__18181\,
            I => \c0.data_10\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__18178\,
            I => \c0.data_10\
        );

    \I__3963\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18169\
        );

    \I__3962\ : InMux
    port map (
            O => \N__18172\,
            I => \N__18166\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__18169\,
            I => \N__18162\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__18166\,
            I => \N__18159\
        );

    \I__3959\ : InMux
    port map (
            O => \N__18165\,
            I => \N__18156\
        );

    \I__3958\ : Span4Mux_v
    port map (
            O => \N__18162\,
            I => \N__18153\
        );

    \I__3957\ : Span4Mux_h
    port map (
            O => \N__18159\,
            I => \N__18150\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__18156\,
            I => data_out_field_19
        );

    \I__3955\ : Odrv4
    port map (
            O => \N__18153\,
            I => data_out_field_19
        );

    \I__3954\ : Odrv4
    port map (
            O => \N__18150\,
            I => data_out_field_19
        );

    \I__3953\ : InMux
    port map (
            O => \N__18143\,
            I => \N__18140\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__18140\,
            I => n8_adj_936
        );

    \I__3951\ : InMux
    port map (
            O => \N__18137\,
            I => \N__18133\
        );

    \I__3950\ : InMux
    port map (
            O => \N__18136\,
            I => \N__18130\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__18133\,
            I => \N__18127\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__18130\,
            I => data_out_6_2
        );

    \I__3947\ : Odrv4
    port map (
            O => \N__18127\,
            I => data_out_6_2
        );

    \I__3946\ : InMux
    port map (
            O => \N__18122\,
            I => \N__18119\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__18119\,
            I => \c0.n2429\
        );

    \I__3944\ : CascadeMux
    port map (
            O => \N__18116\,
            I => \N__18113\
        );

    \I__3943\ : InMux
    port map (
            O => \N__18113\,
            I => \N__18110\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__18110\,
            I => \N__18107\
        );

    \I__3941\ : Span4Mux_h
    port map (
            O => \N__18107\,
            I => \N__18103\
        );

    \I__3940\ : InMux
    port map (
            O => \N__18106\,
            I => \N__18100\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__18103\,
            I => \c0.data_6\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__18100\,
            I => \c0.data_6\
        );

    \I__3937\ : InMux
    port map (
            O => \N__18095\,
            I => \N__18092\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__18092\,
            I => \N__18089\
        );

    \I__3935\ : Span4Mux_h
    port map (
            O => \N__18089\,
            I => \N__18085\
        );

    \I__3934\ : InMux
    port map (
            O => \N__18088\,
            I => \N__18082\
        );

    \I__3933\ : Odrv4
    port map (
            O => \N__18085\,
            I => \c0.data_7\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__18082\,
            I => \c0.data_7\
        );

    \I__3931\ : CascadeMux
    port map (
            O => \N__18077\,
            I => \N__18074\
        );

    \I__3930\ : InMux
    port map (
            O => \N__18074\,
            I => \N__18071\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__18071\,
            I => \N__18068\
        );

    \I__3928\ : Span4Mux_h
    port map (
            O => \N__18068\,
            I => \N__18064\
        );

    \I__3927\ : InMux
    port map (
            O => \N__18067\,
            I => \N__18061\
        );

    \I__3926\ : Odrv4
    port map (
            O => \N__18064\,
            I => \c0.data_14\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__18061\,
            I => \c0.data_14\
        );

    \I__3924\ : InMux
    port map (
            O => \N__18056\,
            I => \N__18052\
        );

    \I__3923\ : InMux
    port map (
            O => \N__18055\,
            I => \N__18049\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__18052\,
            I => \N__18046\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__18049\,
            I => \N__18041\
        );

    \I__3920\ : Span4Mux_v
    port map (
            O => \N__18046\,
            I => \N__18041\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__18041\,
            I => data_out_7_3
        );

    \I__3918\ : CascadeMux
    port map (
            O => \N__18038\,
            I => \N__18035\
        );

    \I__3917\ : InMux
    port map (
            O => \N__18035\,
            I => \N__18032\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__18032\,
            I => \N__18029\
        );

    \I__3915\ : Span4Mux_h
    port map (
            O => \N__18029\,
            I => \N__18025\
        );

    \I__3914\ : InMux
    port map (
            O => \N__18028\,
            I => \N__18022\
        );

    \I__3913\ : Odrv4
    port map (
            O => \N__18025\,
            I => \c0.data_8\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__18022\,
            I => \c0.data_8\
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__18017\,
            I => \n8_adj_932_cascade_\
        );

    \I__3910\ : InMux
    port map (
            O => \N__18014\,
            I => \c0.n3901\
        );

    \I__3909\ : InMux
    port map (
            O => \N__18011\,
            I => \c0.n3902\
        );

    \I__3908\ : InMux
    port map (
            O => \N__18008\,
            I => \c0.n3903\
        );

    \I__3907\ : InMux
    port map (
            O => \N__18005\,
            I => \c0.n3904\
        );

    \I__3906\ : InMux
    port map (
            O => \N__18002\,
            I => \c0.n3905\
        );

    \I__3905\ : InMux
    port map (
            O => \N__17999\,
            I => \N__17996\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__17996\,
            I => \N__17992\
        );

    \I__3903\ : InMux
    port map (
            O => \N__17995\,
            I => \N__17989\
        );

    \I__3902\ : Span4Mux_h
    port map (
            O => \N__17992\,
            I => \N__17986\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__17989\,
            I => data_out_6_1
        );

    \I__3900\ : Odrv4
    port map (
            O => \N__17986\,
            I => data_out_6_1
        );

    \I__3899\ : InMux
    port map (
            O => \N__17981\,
            I => \N__17978\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__17978\,
            I => \N__17974\
        );

    \I__3897\ : InMux
    port map (
            O => \N__17977\,
            I => \N__17971\
        );

    \I__3896\ : Span4Mux_h
    port map (
            O => \N__17974\,
            I => \N__17968\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__17971\,
            I => \c0.data_15\
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__17968\,
            I => \c0.data_15\
        );

    \I__3893\ : InMux
    port map (
            O => \N__17963\,
            I => \N__17960\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__17960\,
            I => \N__17957\
        );

    \I__3891\ : Odrv12
    port map (
            O => \N__17957\,
            I => \c0.n4888\
        );

    \I__3890\ : InMux
    port map (
            O => \N__17954\,
            I => \N__17951\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__17951\,
            I => \c0.rx.n4093\
        );

    \I__3888\ : InMux
    port map (
            O => \N__17948\,
            I => \N__17945\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__17945\,
            I => \c0.rx.n4378\
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__17942\,
            I => \c0.rx.n13_cascade_\
        );

    \I__3885\ : InMux
    port map (
            O => \N__17939\,
            I => \N__17936\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__17936\,
            I => \c0.rx.n6\
        );

    \I__3883\ : CascadeMux
    port map (
            O => \N__17933\,
            I => \N__17926\
        );

    \I__3882\ : InMux
    port map (
            O => \N__17932\,
            I => \N__17921\
        );

    \I__3881\ : InMux
    port map (
            O => \N__17931\,
            I => \N__17914\
        );

    \I__3880\ : InMux
    port map (
            O => \N__17930\,
            I => \N__17914\
        );

    \I__3879\ : InMux
    port map (
            O => \N__17929\,
            I => \N__17914\
        );

    \I__3878\ : InMux
    port map (
            O => \N__17926\,
            I => \N__17907\
        );

    \I__3877\ : InMux
    port map (
            O => \N__17925\,
            I => \N__17907\
        );

    \I__3876\ : InMux
    port map (
            O => \N__17924\,
            I => \N__17907\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__17921\,
            I => n1554
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__17914\,
            I => n1554
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__17907\,
            I => n1554
        );

    \I__3872\ : InMux
    port map (
            O => \N__17900\,
            I => \N__17897\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__17897\,
            I => \N__17894\
        );

    \I__3870\ : Odrv4
    port map (
            O => \N__17894\,
            I => n220
        );

    \I__3869\ : InMux
    port map (
            O => \N__17891\,
            I => \N__17883\
        );

    \I__3868\ : InMux
    port map (
            O => \N__17890\,
            I => \N__17880\
        );

    \I__3867\ : InMux
    port map (
            O => \N__17889\,
            I => \N__17875\
        );

    \I__3866\ : InMux
    port map (
            O => \N__17888\,
            I => \N__17875\
        );

    \I__3865\ : InMux
    port map (
            O => \N__17887\,
            I => \N__17870\
        );

    \I__3864\ : InMux
    port map (
            O => \N__17886\,
            I => \N__17870\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__17883\,
            I => n573
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__17880\,
            I => n573
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__17875\,
            I => n573
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__17870\,
            I => n573
        );

    \I__3859\ : CascadeMux
    port map (
            O => \N__17861\,
            I => \n1554_cascade_\
        );

    \I__3858\ : InMux
    port map (
            O => \N__17858\,
            I => \N__17852\
        );

    \I__3857\ : InMux
    port map (
            O => \N__17857\,
            I => \N__17847\
        );

    \I__3856\ : InMux
    port map (
            O => \N__17856\,
            I => \N__17847\
        );

    \I__3855\ : InMux
    port map (
            O => \N__17855\,
            I => \N__17843\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__17852\,
            I => \N__17838\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__17847\,
            I => \N__17838\
        );

    \I__3852\ : InMux
    port map (
            O => \N__17846\,
            I => \N__17834\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__17843\,
            I => \N__17831\
        );

    \I__3850\ : Span4Mux_v
    port map (
            O => \N__17838\,
            I => \N__17828\
        );

    \I__3849\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17825\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__17834\,
            I => \r_Clock_Count_6\
        );

    \I__3847\ : Odrv4
    port map (
            O => \N__17831\,
            I => \r_Clock_Count_6\
        );

    \I__3846\ : Odrv4
    port map (
            O => \N__17828\,
            I => \r_Clock_Count_6\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__17825\,
            I => \r_Clock_Count_6\
        );

    \I__3844\ : InMux
    port map (
            O => \N__17816\,
            I => \N__17813\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__17813\,
            I => \N__17810\
        );

    \I__3842\ : Span4Mux_s1_v
    port map (
            O => \N__17810\,
            I => \N__17804\
        );

    \I__3841\ : InMux
    port map (
            O => \N__17809\,
            I => \N__17801\
        );

    \I__3840\ : InMux
    port map (
            O => \N__17808\,
            I => \N__17796\
        );

    \I__3839\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17796\
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__17804\,
            I => \c0.rx.n2179\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__17801\,
            I => \c0.rx.n2179\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__17796\,
            I => \c0.rx.n2179\
        );

    \I__3835\ : CascadeMux
    port map (
            O => \N__17789\,
            I => \N__17785\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__17788\,
            I => \N__17782\
        );

    \I__3833\ : InMux
    port map (
            O => \N__17785\,
            I => \N__17773\
        );

    \I__3832\ : InMux
    port map (
            O => \N__17782\,
            I => \N__17773\
        );

    \I__3831\ : InMux
    port map (
            O => \N__17781\,
            I => \N__17768\
        );

    \I__3830\ : InMux
    port map (
            O => \N__17780\,
            I => \N__17768\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__17779\,
            I => \N__17763\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__17778\,
            I => \N__17757\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__17773\,
            I => \N__17753\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__17768\,
            I => \N__17750\
        );

    \I__3825\ : InMux
    port map (
            O => \N__17767\,
            I => \N__17745\
        );

    \I__3824\ : InMux
    port map (
            O => \N__17766\,
            I => \N__17745\
        );

    \I__3823\ : InMux
    port map (
            O => \N__17763\,
            I => \N__17736\
        );

    \I__3822\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17736\
        );

    \I__3821\ : InMux
    port map (
            O => \N__17761\,
            I => \N__17736\
        );

    \I__3820\ : InMux
    port map (
            O => \N__17760\,
            I => \N__17736\
        );

    \I__3819\ : InMux
    port map (
            O => \N__17757\,
            I => \N__17733\
        );

    \I__3818\ : InMux
    port map (
            O => \N__17756\,
            I => \N__17730\
        );

    \I__3817\ : Span4Mux_h
    port map (
            O => \N__17753\,
            I => \N__17727\
        );

    \I__3816\ : Span4Mux_v
    port map (
            O => \N__17750\,
            I => \N__17720\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__17745\,
            I => \N__17720\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__17736\,
            I => \N__17720\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__17733\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__17730\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__3811\ : Odrv4
    port map (
            O => \N__17727\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__3810\ : Odrv4
    port map (
            O => \N__17720\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__3809\ : InMux
    port map (
            O => \N__17711\,
            I => \N__17702\
        );

    \I__3808\ : InMux
    port map (
            O => \N__17710\,
            I => \N__17697\
        );

    \I__3807\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17697\
        );

    \I__3806\ : InMux
    port map (
            O => \N__17708\,
            I => \N__17688\
        );

    \I__3805\ : InMux
    port map (
            O => \N__17707\,
            I => \N__17688\
        );

    \I__3804\ : InMux
    port map (
            O => \N__17706\,
            I => \N__17688\
        );

    \I__3803\ : InMux
    port map (
            O => \N__17705\,
            I => \N__17688\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__17702\,
            I => \N__17680\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__17697\,
            I => \N__17675\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__17688\,
            I => \N__17675\
        );

    \I__3799\ : InMux
    port map (
            O => \N__17687\,
            I => \N__17672\
        );

    \I__3798\ : InMux
    port map (
            O => \N__17686\,
            I => \N__17669\
        );

    \I__3797\ : InMux
    port map (
            O => \N__17685\,
            I => \N__17666\
        );

    \I__3796\ : InMux
    port map (
            O => \N__17684\,
            I => \N__17663\
        );

    \I__3795\ : InMux
    port map (
            O => \N__17683\,
            I => \N__17660\
        );

    \I__3794\ : Span4Mux_h
    port map (
            O => \N__17680\,
            I => \N__17655\
        );

    \I__3793\ : Span4Mux_h
    port map (
            O => \N__17675\,
            I => \N__17655\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__17672\,
            I => \N__17646\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__17669\,
            I => \N__17646\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__17666\,
            I => \N__17646\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__17663\,
            I => \N__17646\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__17660\,
            I => \r_Rx_Data\
        );

    \I__3787\ : Odrv4
    port map (
            O => \N__17655\,
            I => \r_Rx_Data\
        );

    \I__3786\ : Odrv12
    port map (
            O => \N__17646\,
            I => \r_Rx_Data\
        );

    \I__3785\ : InMux
    port map (
            O => \N__17639\,
            I => \N__17634\
        );

    \I__3784\ : InMux
    port map (
            O => \N__17638\,
            I => \N__17622\
        );

    \I__3783\ : InMux
    port map (
            O => \N__17637\,
            I => \N__17622\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__17634\,
            I => \N__17615\
        );

    \I__3781\ : InMux
    port map (
            O => \N__17633\,
            I => \N__17612\
        );

    \I__3780\ : InMux
    port map (
            O => \N__17632\,
            I => \N__17607\
        );

    \I__3779\ : InMux
    port map (
            O => \N__17631\,
            I => \N__17607\
        );

    \I__3778\ : InMux
    port map (
            O => \N__17630\,
            I => \N__17598\
        );

    \I__3777\ : InMux
    port map (
            O => \N__17629\,
            I => \N__17598\
        );

    \I__3776\ : InMux
    port map (
            O => \N__17628\,
            I => \N__17598\
        );

    \I__3775\ : InMux
    port map (
            O => \N__17627\,
            I => \N__17598\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__17622\,
            I => \N__17595\
        );

    \I__3773\ : InMux
    port map (
            O => \N__17621\,
            I => \N__17588\
        );

    \I__3772\ : InMux
    port map (
            O => \N__17620\,
            I => \N__17588\
        );

    \I__3771\ : InMux
    port map (
            O => \N__17619\,
            I => \N__17588\
        );

    \I__3770\ : InMux
    port map (
            O => \N__17618\,
            I => \N__17585\
        );

    \I__3769\ : Span4Mux_h
    port map (
            O => \N__17615\,
            I => \N__17576\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__17612\,
            I => \N__17576\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__17607\,
            I => \N__17576\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__17598\,
            I => \N__17576\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__17595\,
            I => \c0.rx.r_SM_Main_2\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__17588\,
            I => \c0.rx.r_SM_Main_2\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__17585\,
            I => \c0.rx.r_SM_Main_2\
        );

    \I__3762\ : Odrv4
    port map (
            O => \N__17576\,
            I => \c0.rx.r_SM_Main_2\
        );

    \I__3761\ : CascadeMux
    port map (
            O => \N__17567\,
            I => \c0.rx.n4666_cascade_\
        );

    \I__3760\ : InMux
    port map (
            O => \N__17564\,
            I => \N__17561\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__17561\,
            I => \c0.rx.n4667\
        );

    \I__3758\ : InMux
    port map (
            O => \N__17558\,
            I => \N__17545\
        );

    \I__3757\ : InMux
    port map (
            O => \N__17557\,
            I => \N__17545\
        );

    \I__3756\ : InMux
    port map (
            O => \N__17556\,
            I => \N__17537\
        );

    \I__3755\ : InMux
    port map (
            O => \N__17555\,
            I => \N__17537\
        );

    \I__3754\ : InMux
    port map (
            O => \N__17554\,
            I => \N__17528\
        );

    \I__3753\ : InMux
    port map (
            O => \N__17553\,
            I => \N__17528\
        );

    \I__3752\ : InMux
    port map (
            O => \N__17552\,
            I => \N__17528\
        );

    \I__3751\ : InMux
    port map (
            O => \N__17551\,
            I => \N__17528\
        );

    \I__3750\ : CascadeMux
    port map (
            O => \N__17550\,
            I => \N__17525\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__17545\,
            I => \N__17521\
        );

    \I__3748\ : CascadeMux
    port map (
            O => \N__17544\,
            I => \N__17518\
        );

    \I__3747\ : InMux
    port map (
            O => \N__17543\,
            I => \N__17513\
        );

    \I__3746\ : InMux
    port map (
            O => \N__17542\,
            I => \N__17510\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__17537\,
            I => \N__17507\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__17528\,
            I => \N__17504\
        );

    \I__3743\ : InMux
    port map (
            O => \N__17525\,
            I => \N__17499\
        );

    \I__3742\ : InMux
    port map (
            O => \N__17524\,
            I => \N__17499\
        );

    \I__3741\ : Span4Mux_h
    port map (
            O => \N__17521\,
            I => \N__17496\
        );

    \I__3740\ : InMux
    port map (
            O => \N__17518\,
            I => \N__17489\
        );

    \I__3739\ : InMux
    port map (
            O => \N__17517\,
            I => \N__17489\
        );

    \I__3738\ : InMux
    port map (
            O => \N__17516\,
            I => \N__17489\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__17513\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__17510\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__3735\ : Odrv12
    port map (
            O => \N__17507\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__3734\ : Odrv4
    port map (
            O => \N__17504\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__17499\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__3732\ : Odrv4
    port map (
            O => \N__17496\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__17489\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__3730\ : InMux
    port map (
            O => \N__17474\,
            I => \c0.n3899\
        );

    \I__3729\ : InMux
    port map (
            O => \N__17471\,
            I => \c0.n3900\
        );

    \I__3728\ : CascadeMux
    port map (
            O => \N__17468\,
            I => \N__17465\
        );

    \I__3727\ : InMux
    port map (
            O => \N__17465\,
            I => \N__17462\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__17462\,
            I => \N__17459\
        );

    \I__3725\ : Span4Mux_v
    port map (
            O => \N__17459\,
            I => \N__17455\
        );

    \I__3724\ : InMux
    port map (
            O => \N__17458\,
            I => \N__17452\
        );

    \I__3723\ : Sp12to4
    port map (
            O => \N__17455\,
            I => \N__17446\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__17452\,
            I => \N__17446\
        );

    \I__3721\ : InMux
    port map (
            O => \N__17451\,
            I => \N__17443\
        );

    \I__3720\ : Odrv12
    port map (
            O => \N__17446\,
            I => data_in_5_1
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__17443\,
            I => data_in_5_1
        );

    \I__3718\ : CascadeMux
    port map (
            O => \N__17438\,
            I => \N__17435\
        );

    \I__3717\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17432\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__17432\,
            I => \N__17429\
        );

    \I__3715\ : Span4Mux_h
    port map (
            O => \N__17429\,
            I => \N__17426\
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__17426\,
            I => n224
        );

    \I__3713\ : InMux
    port map (
            O => \N__17423\,
            I => \N__17420\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__17420\,
            I => \N__17413\
        );

    \I__3711\ : InMux
    port map (
            O => \N__17419\,
            I => \N__17410\
        );

    \I__3710\ : InMux
    port map (
            O => \N__17418\,
            I => \N__17407\
        );

    \I__3709\ : InMux
    port map (
            O => \N__17417\,
            I => \N__17404\
        );

    \I__3708\ : InMux
    port map (
            O => \N__17416\,
            I => \N__17401\
        );

    \I__3707\ : Span4Mux_h
    port map (
            O => \N__17413\,
            I => \N__17396\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__17410\,
            I => \N__17396\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__17407\,
            I => \r_Clock_Count_2\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__17404\,
            I => \r_Clock_Count_2\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__17401\,
            I => \r_Clock_Count_2\
        );

    \I__3702\ : Odrv4
    port map (
            O => \N__17396\,
            I => \r_Clock_Count_2\
        );

    \I__3701\ : InMux
    port map (
            O => \N__17387\,
            I => \N__17384\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__17384\,
            I => \N__17381\
        );

    \I__3699\ : Odrv12
    port map (
            O => \N__17381\,
            I => \c0.n4528\
        );

    \I__3698\ : InMux
    port map (
            O => \N__17378\,
            I => \N__17375\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__17375\,
            I => \N__17369\
        );

    \I__3696\ : InMux
    port map (
            O => \N__17374\,
            I => \N__17364\
        );

    \I__3695\ : InMux
    port map (
            O => \N__17373\,
            I => \N__17360\
        );

    \I__3694\ : InMux
    port map (
            O => \N__17372\,
            I => \N__17357\
        );

    \I__3693\ : Span4Mux_s2_v
    port map (
            O => \N__17369\,
            I => \N__17354\
        );

    \I__3692\ : InMux
    port map (
            O => \N__17368\,
            I => \N__17349\
        );

    \I__3691\ : InMux
    port map (
            O => \N__17367\,
            I => \N__17349\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__17364\,
            I => \N__17346\
        );

    \I__3689\ : InMux
    port map (
            O => \N__17363\,
            I => \N__17343\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__17360\,
            I => \c0.rx.r_SM_Main_2_N_816_2\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__17357\,
            I => \c0.rx.r_SM_Main_2_N_816_2\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__17354\,
            I => \c0.rx.r_SM_Main_2_N_816_2\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__17349\,
            I => \c0.rx.r_SM_Main_2_N_816_2\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__17346\,
            I => \c0.rx.r_SM_Main_2_N_816_2\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__17343\,
            I => \c0.rx.r_SM_Main_2_N_816_2\
        );

    \I__3682\ : SRMux
    port map (
            O => \N__17330\,
            I => \N__17327\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__17327\,
            I => \N__17324\
        );

    \I__3680\ : Odrv4
    port map (
            O => \N__17324\,
            I => \c0.rx.n1024\
        );

    \I__3679\ : InMux
    port map (
            O => \N__17321\,
            I => \N__17318\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__17318\,
            I => \c0.tx.o_Tx_Serial_N_790\
        );

    \I__3677\ : InMux
    port map (
            O => \N__17315\,
            I => \N__17312\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__17312\,
            I => \c0.tx.n12\
        );

    \I__3675\ : CascadeMux
    port map (
            O => \N__17309\,
            I => \c0.rx.n6_cascade_\
        );

    \I__3674\ : InMux
    port map (
            O => \N__17306\,
            I => \N__17297\
        );

    \I__3673\ : InMux
    port map (
            O => \N__17305\,
            I => \N__17297\
        );

    \I__3672\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17297\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__17297\,
            I => \c0.rx.n357\
        );

    \I__3670\ : InMux
    port map (
            O => \N__17294\,
            I => \N__17291\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__17291\,
            I => \N__17288\
        );

    \I__3668\ : Span4Mux_h
    port map (
            O => \N__17288\,
            I => \N__17284\
        );

    \I__3667\ : InMux
    port map (
            O => \N__17287\,
            I => \N__17281\
        );

    \I__3666\ : Odrv4
    port map (
            O => \N__17284\,
            I => rx_data_1
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__17281\,
            I => rx_data_1
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__17276\,
            I => \N__17273\
        );

    \I__3663\ : InMux
    port map (
            O => \N__17273\,
            I => \N__17269\
        );

    \I__3662\ : InMux
    port map (
            O => \N__17272\,
            I => \N__17266\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__17269\,
            I => \N__17262\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__17266\,
            I => \N__17258\
        );

    \I__3659\ : InMux
    port map (
            O => \N__17265\,
            I => \N__17255\
        );

    \I__3658\ : Span4Mux_v
    port map (
            O => \N__17262\,
            I => \N__17252\
        );

    \I__3657\ : InMux
    port map (
            O => \N__17261\,
            I => \N__17249\
        );

    \I__3656\ : Span4Mux_h
    port map (
            O => \N__17258\,
            I => \N__17242\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__17255\,
            I => \N__17242\
        );

    \I__3654\ : Span4Mux_s2_v
    port map (
            O => \N__17252\,
            I => \N__17242\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__17249\,
            I => data_in_7_1
        );

    \I__3652\ : Odrv4
    port map (
            O => \N__17242\,
            I => data_in_7_1
        );

    \I__3651\ : InMux
    port map (
            O => \N__17237\,
            I => \N__17233\
        );

    \I__3650\ : InMux
    port map (
            O => \N__17236\,
            I => \N__17230\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__17233\,
            I => \N__17227\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__17230\,
            I => \r_Tx_Data_1\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__17227\,
            I => \r_Tx_Data_1\
        );

    \I__3646\ : InMux
    port map (
            O => \N__17222\,
            I => \N__17218\
        );

    \I__3645\ : InMux
    port map (
            O => \N__17221\,
            I => \N__17215\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__17218\,
            I => \N__17212\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__17215\,
            I => \r_Tx_Data_0\
        );

    \I__3642\ : Odrv4
    port map (
            O => \N__17212\,
            I => \r_Tx_Data_0\
        );

    \I__3641\ : InMux
    port map (
            O => \N__17207\,
            I => \N__17203\
        );

    \I__3640\ : InMux
    port map (
            O => \N__17206\,
            I => \N__17200\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__17203\,
            I => \N__17197\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__17200\,
            I => \r_Tx_Data_3\
        );

    \I__3637\ : Odrv12
    port map (
            O => \N__17197\,
            I => \r_Tx_Data_3\
        );

    \I__3636\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17188\
        );

    \I__3635\ : InMux
    port map (
            O => \N__17191\,
            I => \N__17185\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__17188\,
            I => \N__17182\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__17185\,
            I => \r_Tx_Data_2\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__17182\,
            I => \r_Tx_Data_2\
        );

    \I__3631\ : InMux
    port map (
            O => \N__17177\,
            I => \N__17174\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__17174\,
            I => \c0.tx.n4558\
        );

    \I__3629\ : CascadeMux
    port map (
            O => \N__17171\,
            I => \c0.tx.n4559_cascade_\
        );

    \I__3628\ : InMux
    port map (
            O => \N__17168\,
            I => \N__17165\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__17165\,
            I => \c0.tx.n4837\
        );

    \I__3626\ : IoInMux
    port map (
            O => \N__17162\,
            I => \N__17159\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__17159\,
            I => \N__17155\
        );

    \I__3624\ : InMux
    port map (
            O => \N__17158\,
            I => \N__17152\
        );

    \I__3623\ : Span4Mux_s1_v
    port map (
            O => \N__17155\,
            I => \N__17149\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__17152\,
            I => \N__17146\
        );

    \I__3621\ : Sp12to4
    port map (
            O => \N__17149\,
            I => \N__17142\
        );

    \I__3620\ : Span4Mux_s1_v
    port map (
            O => \N__17146\,
            I => \N__17139\
        );

    \I__3619\ : InMux
    port map (
            O => \N__17145\,
            I => \N__17136\
        );

    \I__3618\ : Odrv12
    port map (
            O => \N__17142\,
            I => tx_o
        );

    \I__3617\ : Odrv4
    port map (
            O => \N__17139\,
            I => tx_o
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__17136\,
            I => tx_o
        );

    \I__3615\ : InMux
    port map (
            O => \N__17129\,
            I => \N__17121\
        );

    \I__3614\ : InMux
    port map (
            O => \N__17128\,
            I => \N__17121\
        );

    \I__3613\ : CascadeMux
    port map (
            O => \N__17127\,
            I => \N__17117\
        );

    \I__3612\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17113\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__17121\,
            I => \N__17110\
        );

    \I__3610\ : InMux
    port map (
            O => \N__17120\,
            I => \N__17103\
        );

    \I__3609\ : InMux
    port map (
            O => \N__17117\,
            I => \N__17103\
        );

    \I__3608\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17103\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__17113\,
            I => \N__17080\
        );

    \I__3606\ : Span4Mux_h
    port map (
            O => \N__17110\,
            I => \N__17080\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__17103\,
            I => \N__17080\
        );

    \I__3604\ : InMux
    port map (
            O => \N__17102\,
            I => \N__17075\
        );

    \I__3603\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17075\
        );

    \I__3602\ : InMux
    port map (
            O => \N__17100\,
            I => \N__17070\
        );

    \I__3601\ : InMux
    port map (
            O => \N__17099\,
            I => \N__17070\
        );

    \I__3600\ : CascadeMux
    port map (
            O => \N__17098\,
            I => \N__17066\
        );

    \I__3599\ : InMux
    port map (
            O => \N__17097\,
            I => \N__17053\
        );

    \I__3598\ : InMux
    port map (
            O => \N__17096\,
            I => \N__17050\
        );

    \I__3597\ : InMux
    port map (
            O => \N__17095\,
            I => \N__17046\
        );

    \I__3596\ : InMux
    port map (
            O => \N__17094\,
            I => \N__17041\
        );

    \I__3595\ : InMux
    port map (
            O => \N__17093\,
            I => \N__17041\
        );

    \I__3594\ : InMux
    port map (
            O => \N__17092\,
            I => \N__17038\
        );

    \I__3593\ : InMux
    port map (
            O => \N__17091\,
            I => \N__17033\
        );

    \I__3592\ : InMux
    port map (
            O => \N__17090\,
            I => \N__17033\
        );

    \I__3591\ : InMux
    port map (
            O => \N__17089\,
            I => \N__17028\
        );

    \I__3590\ : InMux
    port map (
            O => \N__17088\,
            I => \N__17028\
        );

    \I__3589\ : InMux
    port map (
            O => \N__17087\,
            I => \N__17025\
        );

    \I__3588\ : Span4Mux_v
    port map (
            O => \N__17080\,
            I => \N__17012\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__17075\,
            I => \N__17012\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__17070\,
            I => \N__17012\
        );

    \I__3585\ : InMux
    port map (
            O => \N__17069\,
            I => \N__17003\
        );

    \I__3584\ : InMux
    port map (
            O => \N__17066\,
            I => \N__17003\
        );

    \I__3583\ : InMux
    port map (
            O => \N__17065\,
            I => \N__17003\
        );

    \I__3582\ : InMux
    port map (
            O => \N__17064\,
            I => \N__17003\
        );

    \I__3581\ : InMux
    port map (
            O => \N__17063\,
            I => \N__16989\
        );

    \I__3580\ : InMux
    port map (
            O => \N__17062\,
            I => \N__16989\
        );

    \I__3579\ : InMux
    port map (
            O => \N__17061\,
            I => \N__16989\
        );

    \I__3578\ : InMux
    port map (
            O => \N__17060\,
            I => \N__16974\
        );

    \I__3577\ : InMux
    port map (
            O => \N__17059\,
            I => \N__16974\
        );

    \I__3576\ : InMux
    port map (
            O => \N__17058\,
            I => \N__16974\
        );

    \I__3575\ : InMux
    port map (
            O => \N__17057\,
            I => \N__16974\
        );

    \I__3574\ : InMux
    port map (
            O => \N__17056\,
            I => \N__16974\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__17053\,
            I => \N__16965\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__17050\,
            I => \N__16965\
        );

    \I__3571\ : InMux
    port map (
            O => \N__17049\,
            I => \N__16962\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__17046\,
            I => \N__16957\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__17041\,
            I => \N__16957\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__17038\,
            I => \N__16954\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__17033\,
            I => \N__16951\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__17028\,
            I => \N__16946\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__17025\,
            I => \N__16946\
        );

    \I__3564\ : InMux
    port map (
            O => \N__17024\,
            I => \N__16943\
        );

    \I__3563\ : InMux
    port map (
            O => \N__17023\,
            I => \N__16940\
        );

    \I__3562\ : InMux
    port map (
            O => \N__17022\,
            I => \N__16937\
        );

    \I__3561\ : InMux
    port map (
            O => \N__17021\,
            I => \N__16932\
        );

    \I__3560\ : InMux
    port map (
            O => \N__17020\,
            I => \N__16932\
        );

    \I__3559\ : InMux
    port map (
            O => \N__17019\,
            I => \N__16929\
        );

    \I__3558\ : Span4Mux_s1_v
    port map (
            O => \N__17012\,
            I => \N__16924\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__17003\,
            I => \N__16924\
        );

    \I__3556\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16908\
        );

    \I__3555\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16908\
        );

    \I__3554\ : InMux
    port map (
            O => \N__17000\,
            I => \N__16908\
        );

    \I__3553\ : InMux
    port map (
            O => \N__16999\,
            I => \N__16908\
        );

    \I__3552\ : InMux
    port map (
            O => \N__16998\,
            I => \N__16902\
        );

    \I__3551\ : InMux
    port map (
            O => \N__16997\,
            I => \N__16899\
        );

    \I__3550\ : InMux
    port map (
            O => \N__16996\,
            I => \N__16896\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__16989\,
            I => \N__16893\
        );

    \I__3548\ : InMux
    port map (
            O => \N__16988\,
            I => \N__16884\
        );

    \I__3547\ : InMux
    port map (
            O => \N__16987\,
            I => \N__16884\
        );

    \I__3546\ : InMux
    port map (
            O => \N__16986\,
            I => \N__16884\
        );

    \I__3545\ : InMux
    port map (
            O => \N__16985\,
            I => \N__16884\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__16974\,
            I => \N__16881\
        );

    \I__3543\ : InMux
    port map (
            O => \N__16973\,
            I => \N__16874\
        );

    \I__3542\ : InMux
    port map (
            O => \N__16972\,
            I => \N__16874\
        );

    \I__3541\ : InMux
    port map (
            O => \N__16971\,
            I => \N__16874\
        );

    \I__3540\ : InMux
    port map (
            O => \N__16970\,
            I => \N__16871\
        );

    \I__3539\ : Span4Mux_v
    port map (
            O => \N__16965\,
            I => \N__16866\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__16962\,
            I => \N__16866\
        );

    \I__3537\ : Span4Mux_s2_v
    port map (
            O => \N__16957\,
            I => \N__16863\
        );

    \I__3536\ : Span4Mux_h
    port map (
            O => \N__16954\,
            I => \N__16856\
        );

    \I__3535\ : Span4Mux_h
    port map (
            O => \N__16951\,
            I => \N__16856\
        );

    \I__3534\ : Span4Mux_v
    port map (
            O => \N__16946\,
            I => \N__16856\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__16943\,
            I => \N__16843\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__16940\,
            I => \N__16843\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__16937\,
            I => \N__16843\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__16932\,
            I => \N__16843\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__16929\,
            I => \N__16843\
        );

    \I__3528\ : Sp12to4
    port map (
            O => \N__16924\,
            I => \N__16843\
        );

    \I__3527\ : InMux
    port map (
            O => \N__16923\,
            I => \N__16832\
        );

    \I__3526\ : InMux
    port map (
            O => \N__16922\,
            I => \N__16832\
        );

    \I__3525\ : InMux
    port map (
            O => \N__16921\,
            I => \N__16832\
        );

    \I__3524\ : InMux
    port map (
            O => \N__16920\,
            I => \N__16832\
        );

    \I__3523\ : InMux
    port map (
            O => \N__16919\,
            I => \N__16832\
        );

    \I__3522\ : InMux
    port map (
            O => \N__16918\,
            I => \N__16827\
        );

    \I__3521\ : InMux
    port map (
            O => \N__16917\,
            I => \N__16827\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__16908\,
            I => \N__16824\
        );

    \I__3519\ : InMux
    port map (
            O => \N__16907\,
            I => \N__16821\
        );

    \I__3518\ : InMux
    port map (
            O => \N__16906\,
            I => \N__16816\
        );

    \I__3517\ : InMux
    port map (
            O => \N__16905\,
            I => \N__16816\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__16902\,
            I => \N__16811\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__16899\,
            I => \N__16811\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__16896\,
            I => \N__16806\
        );

    \I__3513\ : Span4Mux_v
    port map (
            O => \N__16893\,
            I => \N__16806\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__16884\,
            I => \N__16801\
        );

    \I__3511\ : Span4Mux_h
    port map (
            O => \N__16881\,
            I => \N__16801\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__16874\,
            I => \N__16790\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__16871\,
            I => \N__16790\
        );

    \I__3508\ : Span4Mux_s2_v
    port map (
            O => \N__16866\,
            I => \N__16790\
        );

    \I__3507\ : Span4Mux_h
    port map (
            O => \N__16863\,
            I => \N__16790\
        );

    \I__3506\ : Span4Mux_v
    port map (
            O => \N__16856\,
            I => \N__16790\
        );

    \I__3505\ : Span12Mux_s5_h
    port map (
            O => \N__16843\,
            I => \N__16787\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__16832\,
            I => \N__16780\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__16827\,
            I => \N__16780\
        );

    \I__3502\ : Span12Mux_v
    port map (
            O => \N__16824\,
            I => \N__16780\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__16821\,
            I => rx_data_ready_keep
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__16816\,
            I => rx_data_ready_keep
        );

    \I__3499\ : Odrv4
    port map (
            O => \N__16811\,
            I => rx_data_ready_keep
        );

    \I__3498\ : Odrv4
    port map (
            O => \N__16806\,
            I => rx_data_ready_keep
        );

    \I__3497\ : Odrv4
    port map (
            O => \N__16801\,
            I => rx_data_ready_keep
        );

    \I__3496\ : Odrv4
    port map (
            O => \N__16790\,
            I => rx_data_ready_keep
        );

    \I__3495\ : Odrv12
    port map (
            O => \N__16787\,
            I => rx_data_ready_keep
        );

    \I__3494\ : Odrv12
    port map (
            O => \N__16780\,
            I => rx_data_ready_keep
        );

    \I__3493\ : InMux
    port map (
            O => \N__16763\,
            I => \N__16759\
        );

    \I__3492\ : InMux
    port map (
            O => \N__16762\,
            I => \N__16756\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__16759\,
            I => \N__16753\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__16756\,
            I => \N__16746\
        );

    \I__3489\ : Span4Mux_s2_v
    port map (
            O => \N__16753\,
            I => \N__16746\
        );

    \I__3488\ : InMux
    port map (
            O => \N__16752\,
            I => \N__16743\
        );

    \I__3487\ : InMux
    port map (
            O => \N__16751\,
            I => \N__16740\
        );

    \I__3486\ : Odrv4
    port map (
            O => \N__16746\,
            I => data_in_6_1
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__16743\,
            I => data_in_6_1
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__16740\,
            I => data_in_6_1
        );

    \I__3483\ : InMux
    port map (
            O => \N__16733\,
            I => \N__16730\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__16730\,
            I => \c0.n4789\
        );

    \I__3481\ : CascadeMux
    port map (
            O => \N__16727\,
            I => \tx_data_4_keep_cascade_\
        );

    \I__3480\ : InMux
    port map (
            O => \N__16724\,
            I => \N__16720\
        );

    \I__3479\ : InMux
    port map (
            O => \N__16723\,
            I => \N__16717\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__16720\,
            I => \r_Tx_Data_4\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__16717\,
            I => \r_Tx_Data_4\
        );

    \I__3476\ : InMux
    port map (
            O => \N__16712\,
            I => \N__16709\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__16709\,
            I => \c0.n4576\
        );

    \I__3474\ : InMux
    port map (
            O => \N__16706\,
            I => \N__16703\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__16703\,
            I => \N__16700\
        );

    \I__3472\ : Odrv4
    port map (
            O => \N__16700\,
            I => \c0.tx.n4589\
        );

    \I__3471\ : InMux
    port map (
            O => \N__16697\,
            I => \N__16694\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__16694\,
            I => \c0.tx.n4588\
        );

    \I__3469\ : CascadeMux
    port map (
            O => \N__16691\,
            I => \tx_data_5_keep_cascade_\
        );

    \I__3468\ : InMux
    port map (
            O => \N__16688\,
            I => \N__16684\
        );

    \I__3467\ : InMux
    port map (
            O => \N__16687\,
            I => \N__16681\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__16684\,
            I => \r_Tx_Data_5\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__16681\,
            I => \r_Tx_Data_5\
        );

    \I__3464\ : CascadeMux
    port map (
            O => \N__16676\,
            I => \N__16672\
        );

    \I__3463\ : InMux
    port map (
            O => \N__16675\,
            I => \N__16667\
        );

    \I__3462\ : InMux
    port map (
            O => \N__16672\,
            I => \N__16667\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__16667\,
            I => \N__16664\
        );

    \I__3460\ : Odrv12
    port map (
            O => \N__16664\,
            I => \c0.tx.n1588\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__16661\,
            I => \c0.tx.n4715_cascade_\
        );

    \I__3458\ : InMux
    port map (
            O => \N__16658\,
            I => \N__16654\
        );

    \I__3457\ : InMux
    port map (
            O => \N__16657\,
            I => \N__16651\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__16654\,
            I => \r_Tx_Data_7\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__16651\,
            I => \r_Tx_Data_7\
        );

    \I__3454\ : InMux
    port map (
            O => \N__16646\,
            I => \N__16643\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__16643\,
            I => \c0.n4585\
        );

    \I__3452\ : InMux
    port map (
            O => \N__16640\,
            I => \N__16634\
        );

    \I__3451\ : InMux
    port map (
            O => \N__16639\,
            I => \N__16634\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__16634\,
            I => \r_Tx_Data_6\
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__16631\,
            I => \c0.n4861_cascade_\
        );

    \I__3448\ : CascadeMux
    port map (
            O => \N__16628\,
            I => \tx_data_0_keep_cascade_\
        );

    \I__3447\ : CascadeMux
    port map (
            O => \N__16625\,
            I => \N__16622\
        );

    \I__3446\ : InMux
    port map (
            O => \N__16622\,
            I => \N__16619\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__16619\,
            I => \c0.n4586\
        );

    \I__3444\ : InMux
    port map (
            O => \N__16616\,
            I => \N__16613\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__16613\,
            I => \N__16610\
        );

    \I__3442\ : Odrv4
    port map (
            O => \N__16610\,
            I => \c0.n4573\
        );

    \I__3441\ : InMux
    port map (
            O => \N__16607\,
            I => \N__16604\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__16604\,
            I => \c0.n4621\
        );

    \I__3439\ : InMux
    port map (
            O => \N__16601\,
            I => \N__16598\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__16598\,
            I => \c0.n4525\
        );

    \I__3437\ : InMux
    port map (
            O => \N__16595\,
            I => \N__16592\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__16592\,
            I => \N__16588\
        );

    \I__3435\ : InMux
    port map (
            O => \N__16591\,
            I => \N__16585\
        );

    \I__3434\ : Span4Mux_s2_v
    port map (
            O => \N__16588\,
            I => \N__16582\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__16585\,
            I => \N__16579\
        );

    \I__3432\ : Span4Mux_h
    port map (
            O => \N__16582\,
            I => \N__16572\
        );

    \I__3431\ : Span4Mux_h
    port map (
            O => \N__16579\,
            I => \N__16572\
        );

    \I__3430\ : InMux
    port map (
            O => \N__16578\,
            I => \N__16567\
        );

    \I__3429\ : InMux
    port map (
            O => \N__16577\,
            I => \N__16567\
        );

    \I__3428\ : Odrv4
    port map (
            O => \N__16572\,
            I => data_in_6_3
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__16567\,
            I => data_in_6_3
        );

    \I__3426\ : InMux
    port map (
            O => \N__16562\,
            I => \N__16558\
        );

    \I__3425\ : InMux
    port map (
            O => \N__16561\,
            I => \N__16555\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__16558\,
            I => \N__16552\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__16555\,
            I => \N__16549\
        );

    \I__3422\ : Span12Mux_s6_h
    port map (
            O => \N__16552\,
            I => \N__16545\
        );

    \I__3421\ : Span4Mux_h
    port map (
            O => \N__16549\,
            I => \N__16542\
        );

    \I__3420\ : InMux
    port map (
            O => \N__16548\,
            I => \N__16539\
        );

    \I__3419\ : Odrv12
    port map (
            O => \N__16545\,
            I => data_in_5_3
        );

    \I__3418\ : Odrv4
    port map (
            O => \N__16542\,
            I => data_in_5_3
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__16539\,
            I => data_in_5_3
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__16532\,
            I => \c0.n4768_cascade_\
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__16529\,
            I => \tx_data_7_keep_cascade_\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__16526\,
            I => \c0.n4843_cascade_\
        );

    \I__3413\ : CascadeMux
    port map (
            O => \N__16523\,
            I => \tx_data_1_keep_cascade_\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__16520\,
            I => \c0.rx.n4641_cascade_\
        );

    \I__3411\ : InMux
    port map (
            O => \N__16517\,
            I => \N__16514\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__16514\,
            I => \c0.rx.n8\
        );

    \I__3409\ : InMux
    port map (
            O => \N__16511\,
            I => \N__16508\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__16508\,
            I => \c0.rx.n4\
        );

    \I__3407\ : CascadeMux
    port map (
            O => \N__16505\,
            I => \N__16502\
        );

    \I__3406\ : InMux
    port map (
            O => \N__16502\,
            I => \N__16499\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__16499\,
            I => \N__16496\
        );

    \I__3404\ : Odrv12
    port map (
            O => \N__16496\,
            I => \c0.rx.n7\
        );

    \I__3403\ : CascadeMux
    port map (
            O => \N__16493\,
            I => \c0.rx.n4093_cascade_\
        );

    \I__3402\ : InMux
    port map (
            O => \N__16490\,
            I => \N__16487\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__16487\,
            I => \c0.rx.n2246\
        );

    \I__3400\ : CascadeMux
    port map (
            O => \N__16484\,
            I => \N__16481\
        );

    \I__3399\ : InMux
    port map (
            O => \N__16481\,
            I => \N__16478\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__16478\,
            I => n221
        );

    \I__3397\ : InMux
    port map (
            O => \N__16475\,
            I => \N__16470\
        );

    \I__3396\ : InMux
    port map (
            O => \N__16474\,
            I => \N__16467\
        );

    \I__3395\ : InMux
    port map (
            O => \N__16473\,
            I => \N__16464\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__16470\,
            I => \r_Clock_Count_5\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__16467\,
            I => \r_Clock_Count_5\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__16464\,
            I => \r_Clock_Count_5\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__16457\,
            I => \c0.n4783_cascade_\
        );

    \I__3390\ : InMux
    port map (
            O => \N__16454\,
            I => \N__16451\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__16451\,
            I => \N__16448\
        );

    \I__3388\ : Span4Mux_v
    port map (
            O => \N__16448\,
            I => \N__16445\
        );

    \I__3387\ : Odrv4
    port map (
            O => \N__16445\,
            I => \c0.n4526\
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__16442\,
            I => \tx_data_3_keep_cascade_\
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__16439\,
            I => \N__16436\
        );

    \I__3384\ : InMux
    port map (
            O => \N__16436\,
            I => \N__16433\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__16433\,
            I => \c0.n4622\
        );

    \I__3382\ : InMux
    port map (
            O => \N__16430\,
            I => \N__16425\
        );

    \I__3381\ : InMux
    port map (
            O => \N__16429\,
            I => \N__16421\
        );

    \I__3380\ : InMux
    port map (
            O => \N__16428\,
            I => \N__16418\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__16425\,
            I => \N__16415\
        );

    \I__3378\ : InMux
    port map (
            O => \N__16424\,
            I => \N__16412\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__16421\,
            I => \r_Clock_Count_3\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__16418\,
            I => \r_Clock_Count_3\
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__16415\,
            I => \r_Clock_Count_3\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__16412\,
            I => \r_Clock_Count_3\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__16403\,
            I => \c0.rx.n214_cascade_\
        );

    \I__3372\ : CascadeMux
    port map (
            O => \N__16400\,
            I => \c0.rx.n4_cascade_\
        );

    \I__3371\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16388\
        );

    \I__3370\ : InMux
    port map (
            O => \N__16396\,
            I => \N__16383\
        );

    \I__3369\ : InMux
    port map (
            O => \N__16395\,
            I => \N__16383\
        );

    \I__3368\ : InMux
    port map (
            O => \N__16394\,
            I => \N__16378\
        );

    \I__3367\ : InMux
    port map (
            O => \N__16393\,
            I => \N__16378\
        );

    \I__3366\ : InMux
    port map (
            O => \N__16392\,
            I => \N__16373\
        );

    \I__3365\ : InMux
    port map (
            O => \N__16391\,
            I => \N__16373\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__16388\,
            I => \r_Bit_Index_2\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__16383\,
            I => \r_Bit_Index_2\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__16378\,
            I => \r_Bit_Index_2\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__16373\,
            I => \r_Bit_Index_2\
        );

    \I__3360\ : InMux
    port map (
            O => \N__16364\,
            I => \N__16355\
        );

    \I__3359\ : InMux
    port map (
            O => \N__16363\,
            I => \N__16352\
        );

    \I__3358\ : InMux
    port map (
            O => \N__16362\,
            I => \N__16349\
        );

    \I__3357\ : InMux
    port map (
            O => \N__16361\,
            I => \N__16344\
        );

    \I__3356\ : InMux
    port map (
            O => \N__16360\,
            I => \N__16344\
        );

    \I__3355\ : InMux
    port map (
            O => \N__16359\,
            I => \N__16339\
        );

    \I__3354\ : InMux
    port map (
            O => \N__16358\,
            I => \N__16339\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__16355\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__16352\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__16349\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__16344\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__16339\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__3348\ : InMux
    port map (
            O => \N__16328\,
            I => \N__16322\
        );

    \I__3347\ : InMux
    port map (
            O => \N__16327\,
            I => \N__16322\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__16322\,
            I => \N__16319\
        );

    \I__3345\ : Odrv4
    port map (
            O => \N__16319\,
            I => n4_adj_951
        );

    \I__3344\ : InMux
    port map (
            O => \N__16316\,
            I => \N__16313\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__16313\,
            I => \c0.rx.n4679\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__16310\,
            I => \N__16307\
        );

    \I__3341\ : InMux
    port map (
            O => \N__16307\,
            I => \N__16301\
        );

    \I__3340\ : InMux
    port map (
            O => \N__16306\,
            I => \N__16298\
        );

    \I__3339\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16293\
        );

    \I__3338\ : InMux
    port map (
            O => \N__16304\,
            I => \N__16293\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__16301\,
            I => \N__16290\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__16298\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__16293\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__3334\ : Odrv12
    port map (
            O => \N__16290\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__3333\ : InMux
    port map (
            O => \N__16283\,
            I => \N__16280\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__16280\,
            I => n219
        );

    \I__3331\ : InMux
    port map (
            O => \N__16277\,
            I => \N__16274\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__16274\,
            I => \N__16267\
        );

    \I__3329\ : InMux
    port map (
            O => \N__16273\,
            I => \N__16264\
        );

    \I__3328\ : InMux
    port map (
            O => \N__16272\,
            I => \N__16261\
        );

    \I__3327\ : InMux
    port map (
            O => \N__16271\,
            I => \N__16256\
        );

    \I__3326\ : InMux
    port map (
            O => \N__16270\,
            I => \N__16256\
        );

    \I__3325\ : Odrv4
    port map (
            O => \N__16267\,
            I => \r_Clock_Count_7\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__16264\,
            I => \r_Clock_Count_7\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__16261\,
            I => \r_Clock_Count_7\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__16256\,
            I => \r_Clock_Count_7\
        );

    \I__3321\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16244\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__16244\,
            I => \N__16241\
        );

    \I__3319\ : Odrv12
    port map (
            O => \N__16241\,
            I => \c0.rx.n4677\
        );

    \I__3318\ : InMux
    port map (
            O => \N__16238\,
            I => \N__16235\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__16235\,
            I => \N__16232\
        );

    \I__3316\ : Odrv4
    port map (
            O => \N__16232\,
            I => n226
        );

    \I__3315\ : CascadeMux
    port map (
            O => \N__16229\,
            I => \n573_cascade_\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__16226\,
            I => \N__16221\
        );

    \I__3313\ : InMux
    port map (
            O => \N__16225\,
            I => \N__16218\
        );

    \I__3312\ : InMux
    port map (
            O => \N__16224\,
            I => \N__16214\
        );

    \I__3311\ : InMux
    port map (
            O => \N__16221\,
            I => \N__16211\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__16218\,
            I => \N__16208\
        );

    \I__3309\ : InMux
    port map (
            O => \N__16217\,
            I => \N__16205\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__16214\,
            I => \r_Clock_Count_0\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__16211\,
            I => \r_Clock_Count_0\
        );

    \I__3306\ : Odrv4
    port map (
            O => \N__16208\,
            I => \r_Clock_Count_0\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__16205\,
            I => \r_Clock_Count_0\
        );

    \I__3304\ : CascadeMux
    port map (
            O => \N__16196\,
            I => \N__16193\
        );

    \I__3303\ : InMux
    port map (
            O => \N__16193\,
            I => \N__16190\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__16190\,
            I => \N__16187\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__16187\,
            I => n222
        );

    \I__3300\ : InMux
    port map (
            O => \N__16184\,
            I => \N__16181\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__16181\,
            I => \N__16176\
        );

    \I__3298\ : InMux
    port map (
            O => \N__16180\,
            I => \N__16173\
        );

    \I__3297\ : InMux
    port map (
            O => \N__16179\,
            I => \N__16170\
        );

    \I__3296\ : Odrv4
    port map (
            O => \N__16176\,
            I => \r_Clock_Count_4\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__16173\,
            I => \r_Clock_Count_4\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__16170\,
            I => \r_Clock_Count_4\
        );

    \I__3293\ : CascadeMux
    port map (
            O => \N__16163\,
            I => \N__16159\
        );

    \I__3292\ : InMux
    port map (
            O => \N__16162\,
            I => \N__16151\
        );

    \I__3291\ : InMux
    port map (
            O => \N__16159\,
            I => \N__16151\
        );

    \I__3290\ : InMux
    port map (
            O => \N__16158\,
            I => \N__16151\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__16151\,
            I => n1527
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__16148\,
            I => \n1527_cascade_\
        );

    \I__3287\ : InMux
    port map (
            O => \N__16145\,
            I => \N__16136\
        );

    \I__3286\ : InMux
    port map (
            O => \N__16144\,
            I => \N__16136\
        );

    \I__3285\ : InMux
    port map (
            O => \N__16143\,
            I => \N__16136\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__16136\,
            I => n2142
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__16133\,
            I => \N__16128\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__16132\,
            I => \N__16125\
        );

    \I__3281\ : InMux
    port map (
            O => \N__16131\,
            I => \N__16122\
        );

    \I__3280\ : InMux
    port map (
            O => \N__16128\,
            I => \N__16119\
        );

    \I__3279\ : InMux
    port map (
            O => \N__16125\,
            I => \N__16115\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__16122\,
            I => \N__16112\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__16119\,
            I => \N__16109\
        );

    \I__3276\ : InMux
    port map (
            O => \N__16118\,
            I => \N__16106\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__16115\,
            I => \N__16103\
        );

    \I__3274\ : Span4Mux_h
    port map (
            O => \N__16112\,
            I => \N__16100\
        );

    \I__3273\ : Span4Mux_h
    port map (
            O => \N__16109\,
            I => \N__16097\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__16106\,
            I => data_in_7_0
        );

    \I__3271\ : Odrv4
    port map (
            O => \N__16103\,
            I => data_in_7_0
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__16100\,
            I => data_in_7_0
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__16097\,
            I => data_in_7_0
        );

    \I__3268\ : InMux
    port map (
            O => \N__16088\,
            I => \N__16082\
        );

    \I__3267\ : InMux
    port map (
            O => \N__16087\,
            I => \N__16079\
        );

    \I__3266\ : InMux
    port map (
            O => \N__16086\,
            I => \N__16076\
        );

    \I__3265\ : InMux
    port map (
            O => \N__16085\,
            I => \N__16073\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__16082\,
            I => \N__16070\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__16079\,
            I => \N__16067\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__16076\,
            I => data_in_6_0
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__16073\,
            I => data_in_6_0
        );

    \I__3260\ : Odrv12
    port map (
            O => \N__16070\,
            I => data_in_6_0
        );

    \I__3259\ : Odrv4
    port map (
            O => \N__16067\,
            I => data_in_6_0
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__16058\,
            I => \N__16055\
        );

    \I__3257\ : InMux
    port map (
            O => \N__16055\,
            I => \N__16052\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__16052\,
            I => \c0.rx.n232\
        );

    \I__3255\ : CascadeMux
    port map (
            O => \N__16049\,
            I => \c0.rx.r_SM_Main_2_N_816_2_cascade_\
        );

    \I__3254\ : InMux
    port map (
            O => \N__16046\,
            I => \N__16043\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__16043\,
            I => \N__16040\
        );

    \I__3252\ : Span4Mux_s2_v
    port map (
            O => \N__16040\,
            I => \N__16037\
        );

    \I__3251\ : Odrv4
    port map (
            O => \N__16037\,
            I => \c0.rx.n4678\
        );

    \I__3250\ : CascadeMux
    port map (
            O => \N__16034\,
            I => \N__16028\
        );

    \I__3249\ : InMux
    port map (
            O => \N__16033\,
            I => \N__16021\
        );

    \I__3248\ : InMux
    port map (
            O => \N__16032\,
            I => \N__16021\
        );

    \I__3247\ : InMux
    port map (
            O => \N__16031\,
            I => \N__16016\
        );

    \I__3246\ : InMux
    port map (
            O => \N__16028\,
            I => \N__16016\
        );

    \I__3245\ : InMux
    port map (
            O => \N__16027\,
            I => \N__16011\
        );

    \I__3244\ : InMux
    port map (
            O => \N__16026\,
            I => \N__16011\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__16021\,
            I => \r_Bit_Index_0\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__16016\,
            I => \r_Bit_Index_0\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__16011\,
            I => \r_Bit_Index_0\
        );

    \I__3240\ : CascadeMux
    port map (
            O => \N__16004\,
            I => \N__16001\
        );

    \I__3239\ : InMux
    port map (
            O => \N__16001\,
            I => \N__15997\
        );

    \I__3238\ : InMux
    port map (
            O => \N__16000\,
            I => \N__15994\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__15997\,
            I => n4_adj_943
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__15994\,
            I => n4_adj_943
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__15989\,
            I => \N__15986\
        );

    \I__3234\ : InMux
    port map (
            O => \N__15986\,
            I => \N__15983\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__15983\,
            I => \N__15980\
        );

    \I__3232\ : Odrv4
    port map (
            O => \N__15980\,
            I => n223
        );

    \I__3231\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15974\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__15974\,
            I => \N__15970\
        );

    \I__3229\ : InMux
    port map (
            O => \N__15973\,
            I => \N__15967\
        );

    \I__3228\ : Odrv4
    port map (
            O => \N__15970\,
            I => \c0.rx.n214\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__15967\,
            I => \c0.rx.n214\
        );

    \I__3226\ : InMux
    port map (
            O => \N__15962\,
            I => \N__15959\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__15959\,
            I => \N__15956\
        );

    \I__3224\ : Span4Mux_h
    port map (
            O => \N__15956\,
            I => \N__15953\
        );

    \I__3223\ : Odrv4
    port map (
            O => \N__15953\,
            I => \c0.n4408\
        );

    \I__3222\ : InMux
    port map (
            O => \N__15950\,
            I => \N__15947\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__15947\,
            I => \N__15944\
        );

    \I__3220\ : Span4Mux_h
    port map (
            O => \N__15944\,
            I => \N__15940\
        );

    \I__3219\ : InMux
    port map (
            O => \N__15943\,
            I => \N__15937\
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__15940\,
            I => \c0.n1271\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__15937\,
            I => \c0.n1271\
        );

    \I__3216\ : InMux
    port map (
            O => \N__15932\,
            I => \N__15929\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__15929\,
            I => \N__15926\
        );

    \I__3214\ : Span4Mux_h
    port map (
            O => \N__15926\,
            I => \N__15923\
        );

    \I__3213\ : Odrv4
    port map (
            O => \N__15923\,
            I => \c0.n4409\
        );

    \I__3212\ : CascadeMux
    port map (
            O => \N__15920\,
            I => \c0.rx.n232_cascade_\
        );

    \I__3211\ : InMux
    port map (
            O => \N__15917\,
            I => \N__15914\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__15914\,
            I => \N__15911\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__15911\,
            I => \c0.n4516\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__15908\,
            I => \c0.rx.n1464_cascade_\
        );

    \I__3207\ : CascadeMux
    port map (
            O => \N__15905\,
            I => \N__15902\
        );

    \I__3206\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15899\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__15899\,
            I => \N__15895\
        );

    \I__3204\ : InMux
    port map (
            O => \N__15898\,
            I => \N__15892\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__15895\,
            I => \c0.data_1\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__15892\,
            I => \c0.data_1\
        );

    \I__3201\ : InMux
    port map (
            O => \N__15887\,
            I => \N__15884\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__15884\,
            I => \N__15879\
        );

    \I__3199\ : CascadeMux
    port map (
            O => \N__15883\,
            I => \N__15875\
        );

    \I__3198\ : InMux
    port map (
            O => \N__15882\,
            I => \N__15872\
        );

    \I__3197\ : Span4Mux_h
    port map (
            O => \N__15879\,
            I => \N__15869\
        );

    \I__3196\ : InMux
    port map (
            O => \N__15878\,
            I => \N__15866\
        );

    \I__3195\ : InMux
    port map (
            O => \N__15875\,
            I => \N__15863\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__15872\,
            I => data_in_7_2
        );

    \I__3193\ : Odrv4
    port map (
            O => \N__15869\,
            I => data_in_7_2
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__15866\,
            I => data_in_7_2
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__15863\,
            I => data_in_7_2
        );

    \I__3190\ : InMux
    port map (
            O => \N__15854\,
            I => \N__15849\
        );

    \I__3189\ : InMux
    port map (
            O => \N__15853\,
            I => \N__15846\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__15852\,
            I => \N__15842\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__15849\,
            I => \N__15839\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__15846\,
            I => \N__15836\
        );

    \I__3185\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15833\
        );

    \I__3184\ : InMux
    port map (
            O => \N__15842\,
            I => \N__15830\
        );

    \I__3183\ : Span4Mux_h
    port map (
            O => \N__15839\,
            I => \N__15825\
        );

    \I__3182\ : Span4Mux_h
    port map (
            O => \N__15836\,
            I => \N__15825\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__15833\,
            I => data_in_6_2
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__15830\,
            I => data_in_6_2
        );

    \I__3179\ : Odrv4
    port map (
            O => \N__15825\,
            I => data_in_6_2
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__15818\,
            I => \c0.n4517_cascade_\
        );

    \I__3177\ : CascadeMux
    port map (
            O => \N__15815\,
            I => \c0.n4867_cascade_\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__15812\,
            I => \tx_data_2_keep_cascade_\
        );

    \I__3175\ : InMux
    port map (
            O => \N__15809\,
            I => \N__15806\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__15806\,
            I => \c0.n4564\
        );

    \I__3173\ : InMux
    port map (
            O => \N__15803\,
            I => \c0.n3916\
        );

    \I__3172\ : InMux
    port map (
            O => \N__15800\,
            I => \c0.n3917\
        );

    \I__3171\ : InMux
    port map (
            O => \N__15797\,
            I => \c0.n3918\
        );

    \I__3170\ : InMux
    port map (
            O => \N__15794\,
            I => \c0.n3919\
        );

    \I__3169\ : InMux
    port map (
            O => \N__15791\,
            I => \c0.n3920\
        );

    \I__3168\ : CascadeMux
    port map (
            O => \N__15788\,
            I => \N__15779\
        );

    \I__3167\ : CascadeMux
    port map (
            O => \N__15787\,
            I => \N__15774\
        );

    \I__3166\ : CascadeMux
    port map (
            O => \N__15786\,
            I => \N__15771\
        );

    \I__3165\ : CascadeMux
    port map (
            O => \N__15785\,
            I => \N__15768\
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__15784\,
            I => \N__15762\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__15783\,
            I => \N__15757\
        );

    \I__3162\ : CascadeMux
    port map (
            O => \N__15782\,
            I => \N__15754\
        );

    \I__3161\ : InMux
    port map (
            O => \N__15779\,
            I => \N__15751\
        );

    \I__3160\ : InMux
    port map (
            O => \N__15778\,
            I => \N__15748\
        );

    \I__3159\ : CascadeMux
    port map (
            O => \N__15777\,
            I => \N__15743\
        );

    \I__3158\ : InMux
    port map (
            O => \N__15774\,
            I => \N__15740\
        );

    \I__3157\ : InMux
    port map (
            O => \N__15771\,
            I => \N__15735\
        );

    \I__3156\ : InMux
    port map (
            O => \N__15768\,
            I => \N__15735\
        );

    \I__3155\ : InMux
    port map (
            O => \N__15767\,
            I => \N__15732\
        );

    \I__3154\ : InMux
    port map (
            O => \N__15766\,
            I => \N__15728\
        );

    \I__3153\ : InMux
    port map (
            O => \N__15765\,
            I => \N__15723\
        );

    \I__3152\ : InMux
    port map (
            O => \N__15762\,
            I => \N__15723\
        );

    \I__3151\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15720\
        );

    \I__3150\ : InMux
    port map (
            O => \N__15760\,
            I => \N__15717\
        );

    \I__3149\ : InMux
    port map (
            O => \N__15757\,
            I => \N__15714\
        );

    \I__3148\ : InMux
    port map (
            O => \N__15754\,
            I => \N__15711\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__15751\,
            I => \N__15706\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__15748\,
            I => \N__15706\
        );

    \I__3145\ : InMux
    port map (
            O => \N__15747\,
            I => \N__15698\
        );

    \I__3144\ : InMux
    port map (
            O => \N__15746\,
            I => \N__15698\
        );

    \I__3143\ : InMux
    port map (
            O => \N__15743\,
            I => \N__15698\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__15740\,
            I => \N__15693\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__15735\,
            I => \N__15693\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__15732\,
            I => \N__15690\
        );

    \I__3139\ : InMux
    port map (
            O => \N__15731\,
            I => \N__15687\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__15728\,
            I => \N__15672\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__15723\,
            I => \N__15672\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__15720\,
            I => \N__15672\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__15717\,
            I => \N__15672\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__15714\,
            I => \N__15672\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__15711\,
            I => \N__15672\
        );

    \I__3132\ : Span4Mux_s1_h
    port map (
            O => \N__15706\,
            I => \N__15672\
        );

    \I__3131\ : InMux
    port map (
            O => \N__15705\,
            I => \N__15669\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__15698\,
            I => \N__15664\
        );

    \I__3129\ : Span4Mux_h
    port map (
            O => \N__15693\,
            I => \N__15664\
        );

    \I__3128\ : Span4Mux_h
    port map (
            O => \N__15690\,
            I => \N__15661\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__15687\,
            I => \N__15656\
        );

    \I__3126\ : Span4Mux_v
    port map (
            O => \N__15672\,
            I => \N__15656\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__15669\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__3124\ : Odrv4
    port map (
            O => \N__15664\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__15661\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__15656\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__3121\ : InMux
    port map (
            O => \N__15647\,
            I => \N__15641\
        );

    \I__3120\ : InMux
    port map (
            O => \N__15646\,
            I => \N__15641\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__15641\,
            I => \N__15632\
        );

    \I__3118\ : InMux
    port map (
            O => \N__15640\,
            I => \N__15629\
        );

    \I__3117\ : InMux
    port map (
            O => \N__15639\,
            I => \N__15626\
        );

    \I__3116\ : InMux
    port map (
            O => \N__15638\,
            I => \N__15623\
        );

    \I__3115\ : InMux
    port map (
            O => \N__15637\,
            I => \N__15620\
        );

    \I__3114\ : InMux
    port map (
            O => \N__15636\,
            I => \N__15617\
        );

    \I__3113\ : InMux
    port map (
            O => \N__15635\,
            I => \N__15614\
        );

    \I__3112\ : Span4Mux_s2_h
    port map (
            O => \N__15632\,
            I => \N__15609\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__15629\,
            I => \N__15609\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__15626\,
            I => \N__15605\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__15623\,
            I => \N__15601\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__15620\,
            I => \N__15598\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__15617\,
            I => \N__15595\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__15614\,
            I => \N__15590\
        );

    \I__3105\ : Span4Mux_v
    port map (
            O => \N__15609\,
            I => \N__15590\
        );

    \I__3104\ : InMux
    port map (
            O => \N__15608\,
            I => \N__15587\
        );

    \I__3103\ : Span4Mux_h
    port map (
            O => \N__15605\,
            I => \N__15584\
        );

    \I__3102\ : InMux
    port map (
            O => \N__15604\,
            I => \N__15581\
        );

    \I__3101\ : Span4Mux_h
    port map (
            O => \N__15601\,
            I => \N__15578\
        );

    \I__3100\ : Span4Mux_v
    port map (
            O => \N__15598\,
            I => \N__15571\
        );

    \I__3099\ : Span4Mux_v
    port map (
            O => \N__15595\,
            I => \N__15571\
        );

    \I__3098\ : Span4Mux_s2_h
    port map (
            O => \N__15590\,
            I => \N__15571\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__15587\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__15584\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__15581\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__3094\ : Odrv4
    port map (
            O => \N__15578\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__3093\ : Odrv4
    port map (
            O => \N__15571\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__3092\ : InMux
    port map (
            O => \N__15560\,
            I => \N__15555\
        );

    \I__3091\ : InMux
    port map (
            O => \N__15559\,
            I => \N__15552\
        );

    \I__3090\ : InMux
    port map (
            O => \N__15558\,
            I => \N__15549\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__15555\,
            I => \N__15537\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__15552\,
            I => \N__15537\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__15549\,
            I => \N__15537\
        );

    \I__3086\ : InMux
    port map (
            O => \N__15548\,
            I => \N__15532\
        );

    \I__3085\ : InMux
    port map (
            O => \N__15547\,
            I => \N__15532\
        );

    \I__3084\ : CascadeMux
    port map (
            O => \N__15546\,
            I => \N__15529\
        );

    \I__3083\ : InMux
    port map (
            O => \N__15545\,
            I => \N__15522\
        );

    \I__3082\ : InMux
    port map (
            O => \N__15544\,
            I => \N__15507\
        );

    \I__3081\ : Span4Mux_v
    port map (
            O => \N__15537\,
            I => \N__15502\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__15532\,
            I => \N__15502\
        );

    \I__3079\ : InMux
    port map (
            O => \N__15529\,
            I => \N__15499\
        );

    \I__3078\ : InMux
    port map (
            O => \N__15528\,
            I => \N__15496\
        );

    \I__3077\ : InMux
    port map (
            O => \N__15527\,
            I => \N__15492\
        );

    \I__3076\ : InMux
    port map (
            O => \N__15526\,
            I => \N__15487\
        );

    \I__3075\ : InMux
    port map (
            O => \N__15525\,
            I => \N__15487\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__15522\,
            I => \N__15484\
        );

    \I__3073\ : InMux
    port map (
            O => \N__15521\,
            I => \N__15481\
        );

    \I__3072\ : InMux
    port map (
            O => \N__15520\,
            I => \N__15478\
        );

    \I__3071\ : InMux
    port map (
            O => \N__15519\,
            I => \N__15475\
        );

    \I__3070\ : InMux
    port map (
            O => \N__15518\,
            I => \N__15472\
        );

    \I__3069\ : InMux
    port map (
            O => \N__15517\,
            I => \N__15461\
        );

    \I__3068\ : InMux
    port map (
            O => \N__15516\,
            I => \N__15461\
        );

    \I__3067\ : InMux
    port map (
            O => \N__15515\,
            I => \N__15454\
        );

    \I__3066\ : InMux
    port map (
            O => \N__15514\,
            I => \N__15454\
        );

    \I__3065\ : InMux
    port map (
            O => \N__15513\,
            I => \N__15454\
        );

    \I__3064\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15449\
        );

    \I__3063\ : InMux
    port map (
            O => \N__15511\,
            I => \N__15449\
        );

    \I__3062\ : InMux
    port map (
            O => \N__15510\,
            I => \N__15446\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__15507\,
            I => \N__15443\
        );

    \I__3060\ : Span4Mux_s3_v
    port map (
            O => \N__15502\,
            I => \N__15436\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__15499\,
            I => \N__15436\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__15496\,
            I => \N__15436\
        );

    \I__3057\ : CascadeMux
    port map (
            O => \N__15495\,
            I => \N__15433\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__15492\,
            I => \N__15427\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__15487\,
            I => \N__15418\
        );

    \I__3054\ : Span4Mux_v
    port map (
            O => \N__15484\,
            I => \N__15418\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__15481\,
            I => \N__15418\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__15478\,
            I => \N__15418\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__15475\,
            I => \N__15413\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__15472\,
            I => \N__15413\
        );

    \I__3049\ : InMux
    port map (
            O => \N__15471\,
            I => \N__15410\
        );

    \I__3048\ : InMux
    port map (
            O => \N__15470\,
            I => \N__15407\
        );

    \I__3047\ : InMux
    port map (
            O => \N__15469\,
            I => \N__15402\
        );

    \I__3046\ : InMux
    port map (
            O => \N__15468\,
            I => \N__15402\
        );

    \I__3045\ : InMux
    port map (
            O => \N__15467\,
            I => \N__15397\
        );

    \I__3044\ : InMux
    port map (
            O => \N__15466\,
            I => \N__15397\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__15461\,
            I => \N__15390\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__15454\,
            I => \N__15390\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__15449\,
            I => \N__15390\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__15446\,
            I => \N__15383\
        );

    \I__3039\ : Span4Mux_s3_v
    port map (
            O => \N__15443\,
            I => \N__15383\
        );

    \I__3038\ : Span4Mux_h
    port map (
            O => \N__15436\,
            I => \N__15383\
        );

    \I__3037\ : InMux
    port map (
            O => \N__15433\,
            I => \N__15380\
        );

    \I__3036\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15377\
        );

    \I__3035\ : InMux
    port map (
            O => \N__15431\,
            I => \N__15374\
        );

    \I__3034\ : InMux
    port map (
            O => \N__15430\,
            I => \N__15371\
        );

    \I__3033\ : Span4Mux_v
    port map (
            O => \N__15427\,
            I => \N__15364\
        );

    \I__3032\ : Span4Mux_v
    port map (
            O => \N__15418\,
            I => \N__15364\
        );

    \I__3031\ : Span4Mux_v
    port map (
            O => \N__15413\,
            I => \N__15364\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__15410\,
            I => \N__15355\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__15407\,
            I => \N__15355\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__15402\,
            I => \N__15355\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__15397\,
            I => \N__15355\
        );

    \I__3026\ : Span4Mux_h
    port map (
            O => \N__15390\,
            I => \N__15352\
        );

    \I__3025\ : Span4Mux_v
    port map (
            O => \N__15383\,
            I => \N__15349\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__15380\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__15377\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__15374\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__15371\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__3020\ : Odrv4
    port map (
            O => \N__15364\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__3019\ : Odrv12
    port map (
            O => \N__15355\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__3018\ : Odrv4
    port map (
            O => \N__15352\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__15349\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__3016\ : InMux
    port map (
            O => \N__15332\,
            I => \N__15329\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__15329\,
            I => \N__15324\
        );

    \I__3014\ : InMux
    port map (
            O => \N__15328\,
            I => \N__15321\
        );

    \I__3013\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15318\
        );

    \I__3012\ : Span4Mux_h
    port map (
            O => \N__15324\,
            I => \N__15315\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__15321\,
            I => \N__15310\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__15318\,
            I => \N__15310\
        );

    \I__3009\ : Odrv4
    port map (
            O => \N__15315\,
            I => \c0.FRAME_MATCHER_wait_for_transmission_N_423\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__15310\,
            I => \c0.FRAME_MATCHER_wait_for_transmission_N_423\
        );

    \I__3007\ : CascadeMux
    port map (
            O => \N__15305\,
            I => \N__15302\
        );

    \I__3006\ : InMux
    port map (
            O => \N__15302\,
            I => \N__15298\
        );

    \I__3005\ : InMux
    port map (
            O => \N__15301\,
            I => \N__15295\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__15298\,
            I => \c0.data_9\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__15295\,
            I => \c0.data_9\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__15290\,
            I => \c0.n4619_cascade_\
        );

    \I__3001\ : InMux
    port map (
            O => \N__15287\,
            I => \c0.n3907\
        );

    \I__3000\ : InMux
    port map (
            O => \N__15284\,
            I => \c0.n3908\
        );

    \I__2999\ : InMux
    port map (
            O => \N__15281\,
            I => \c0.n3909\
        );

    \I__2998\ : InMux
    port map (
            O => \N__15278\,
            I => \c0.n3910\
        );

    \I__2997\ : InMux
    port map (
            O => \N__15275\,
            I => \c0.n3911\
        );

    \I__2996\ : InMux
    port map (
            O => \N__15272\,
            I => \c0.n3912\
        );

    \I__2995\ : InMux
    port map (
            O => \N__15269\,
            I => \bfn_6_26_0_\
        );

    \I__2994\ : InMux
    port map (
            O => \N__15266\,
            I => \c0.n3914\
        );

    \I__2993\ : InMux
    port map (
            O => \N__15263\,
            I => \c0.n3915\
        );

    \I__2992\ : InMux
    port map (
            O => \N__15260\,
            I => \c0.rx.n3886\
        );

    \I__2991\ : InMux
    port map (
            O => \N__15257\,
            I => \c0.rx.n3887\
        );

    \I__2990\ : InMux
    port map (
            O => \N__15254\,
            I => \c0.rx.n3888\
        );

    \I__2989\ : InMux
    port map (
            O => \N__15251\,
            I => \c0.rx.n3889\
        );

    \I__2988\ : InMux
    port map (
            O => \N__15248\,
            I => \c0.rx.n3890\
        );

    \I__2987\ : InMux
    port map (
            O => \N__15245\,
            I => \N__15242\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__15242\,
            I => \N__15239\
        );

    \I__2985\ : Span4Mux_h
    port map (
            O => \N__15239\,
            I => \N__15236\
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__15236\,
            I => n1695
        );

    \I__2983\ : InMux
    port map (
            O => \N__15233\,
            I => \N__15230\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__15230\,
            I => \N__15219\
        );

    \I__2981\ : InMux
    port map (
            O => \N__15229\,
            I => \N__15208\
        );

    \I__2980\ : InMux
    port map (
            O => \N__15228\,
            I => \N__15208\
        );

    \I__2979\ : InMux
    port map (
            O => \N__15227\,
            I => \N__15208\
        );

    \I__2978\ : InMux
    port map (
            O => \N__15226\,
            I => \N__15208\
        );

    \I__2977\ : InMux
    port map (
            O => \N__15225\,
            I => \N__15208\
        );

    \I__2976\ : InMux
    port map (
            O => \N__15224\,
            I => \N__15201\
        );

    \I__2975\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15201\
        );

    \I__2974\ : InMux
    port map (
            O => \N__15222\,
            I => \N__15201\
        );

    \I__2973\ : Odrv12
    port map (
            O => \N__15219\,
            I => n6_adj_940
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__15208\,
            I => n6_adj_940
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__15201\,
            I => n6_adj_940
        );

    \I__2970\ : InMux
    port map (
            O => \N__15194\,
            I => \N__15189\
        );

    \I__2969\ : InMux
    port map (
            O => \N__15193\,
            I => \N__15186\
        );

    \I__2968\ : InMux
    port map (
            O => \N__15192\,
            I => \N__15183\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__15189\,
            I => \N__15178\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__15186\,
            I => \N__15178\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__15183\,
            I => \N__15175\
        );

    \I__2964\ : Span4Mux_h
    port map (
            O => \N__15178\,
            I => \N__15172\
        );

    \I__2963\ : Span4Mux_h
    port map (
            O => \N__15175\,
            I => \N__15169\
        );

    \I__2962\ : Odrv4
    port map (
            O => \N__15172\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__2961\ : Odrv4
    port map (
            O => \N__15169\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__2960\ : InMux
    port map (
            O => \N__15164\,
            I => \bfn_6_25_0_\
        );

    \I__2959\ : InMux
    port map (
            O => \N__15161\,
            I => \c0.n3906\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__15158\,
            I => \n1222_cascade_\
        );

    \I__2957\ : InMux
    port map (
            O => \N__15155\,
            I => \N__15151\
        );

    \I__2956\ : InMux
    port map (
            O => \N__15154\,
            I => \N__15148\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__15151\,
            I => rx_data_0
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__15148\,
            I => rx_data_0
        );

    \I__2953\ : InMux
    port map (
            O => \N__15143\,
            I => \N__15139\
        );

    \I__2952\ : InMux
    port map (
            O => \N__15142\,
            I => \N__15136\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__15139\,
            I => \N__15131\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__15136\,
            I => \N__15131\
        );

    \I__2949\ : Odrv12
    port map (
            O => \N__15131\,
            I => n4_adj_950
        );

    \I__2948\ : InMux
    port map (
            O => \N__15128\,
            I => \N__15122\
        );

    \I__2947\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15122\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__15122\,
            I => n4
        );

    \I__2945\ : InMux
    port map (
            O => \N__15119\,
            I => \N__15116\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__15116\,
            I => \c0.rx.n2269\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__15113\,
            I => \c0.rx.n2269_cascade_\
        );

    \I__2942\ : InMux
    port map (
            O => \N__15110\,
            I => \N__15107\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__15107\,
            I => \N__15102\
        );

    \I__2940\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15097\
        );

    \I__2939\ : InMux
    port map (
            O => \N__15105\,
            I => \N__15097\
        );

    \I__2938\ : Odrv4
    port map (
            O => \N__15102\,
            I => n1227
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__15097\,
            I => n1227
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__15092\,
            I => \n1227_cascade_\
        );

    \I__2935\ : InMux
    port map (
            O => \N__15089\,
            I => \bfn_5_32_0_\
        );

    \I__2934\ : InMux
    port map (
            O => \N__15086\,
            I => \c0.rx.n3884\
        );

    \I__2933\ : InMux
    port map (
            O => \N__15083\,
            I => \c0.rx.n3885\
        );

    \I__2932\ : InMux
    port map (
            O => \N__15080\,
            I => \N__15075\
        );

    \I__2931\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15072\
        );

    \I__2930\ : InMux
    port map (
            O => \N__15078\,
            I => \N__15068\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__15075\,
            I => \N__15065\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__15072\,
            I => \N__15062\
        );

    \I__2927\ : InMux
    port map (
            O => \N__15071\,
            I => \N__15059\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__15068\,
            I => \N__15056\
        );

    \I__2925\ : Odrv12
    port map (
            O => \N__15065\,
            I => data_in_1_2
        );

    \I__2924\ : Odrv4
    port map (
            O => \N__15062\,
            I => data_in_1_2
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__15059\,
            I => data_in_1_2
        );

    \I__2922\ : Odrv4
    port map (
            O => \N__15056\,
            I => data_in_1_2
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__15047\,
            I => \N__15039\
        );

    \I__2920\ : InMux
    port map (
            O => \N__15046\,
            I => \N__15006\
        );

    \I__2919\ : InMux
    port map (
            O => \N__15045\,
            I => \N__15001\
        );

    \I__2918\ : InMux
    port map (
            O => \N__15044\,
            I => \N__15001\
        );

    \I__2917\ : CascadeMux
    port map (
            O => \N__15043\,
            I => \N__14998\
        );

    \I__2916\ : InMux
    port map (
            O => \N__15042\,
            I => \N__14994\
        );

    \I__2915\ : InMux
    port map (
            O => \N__15039\,
            I => \N__14989\
        );

    \I__2914\ : InMux
    port map (
            O => \N__15038\,
            I => \N__14989\
        );

    \I__2913\ : InMux
    port map (
            O => \N__15037\,
            I => \N__14984\
        );

    \I__2912\ : InMux
    port map (
            O => \N__15036\,
            I => \N__14984\
        );

    \I__2911\ : InMux
    port map (
            O => \N__15035\,
            I => \N__14979\
        );

    \I__2910\ : InMux
    port map (
            O => \N__15034\,
            I => \N__14979\
        );

    \I__2909\ : InMux
    port map (
            O => \N__15033\,
            I => \N__14974\
        );

    \I__2908\ : InMux
    port map (
            O => \N__15032\,
            I => \N__14965\
        );

    \I__2907\ : InMux
    port map (
            O => \N__15031\,
            I => \N__14965\
        );

    \I__2906\ : InMux
    port map (
            O => \N__15030\,
            I => \N__14965\
        );

    \I__2905\ : InMux
    port map (
            O => \N__15029\,
            I => \N__14965\
        );

    \I__2904\ : InMux
    port map (
            O => \N__15028\,
            I => \N__14953\
        );

    \I__2903\ : InMux
    port map (
            O => \N__15027\,
            I => \N__14950\
        );

    \I__2902\ : InMux
    port map (
            O => \N__15026\,
            I => \N__14947\
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__15025\,
            I => \N__14941\
        );

    \I__2900\ : InMux
    port map (
            O => \N__15024\,
            I => \N__14919\
        );

    \I__2899\ : InMux
    port map (
            O => \N__15023\,
            I => \N__14919\
        );

    \I__2898\ : InMux
    port map (
            O => \N__15022\,
            I => \N__14919\
        );

    \I__2897\ : InMux
    port map (
            O => \N__15021\,
            I => \N__14919\
        );

    \I__2896\ : InMux
    port map (
            O => \N__15020\,
            I => \N__14914\
        );

    \I__2895\ : InMux
    port map (
            O => \N__15019\,
            I => \N__14914\
        );

    \I__2894\ : InMux
    port map (
            O => \N__15018\,
            I => \N__14901\
        );

    \I__2893\ : InMux
    port map (
            O => \N__15017\,
            I => \N__14901\
        );

    \I__2892\ : InMux
    port map (
            O => \N__15016\,
            I => \N__14901\
        );

    \I__2891\ : InMux
    port map (
            O => \N__15015\,
            I => \N__14901\
        );

    \I__2890\ : InMux
    port map (
            O => \N__15014\,
            I => \N__14901\
        );

    \I__2889\ : InMux
    port map (
            O => \N__15013\,
            I => \N__14901\
        );

    \I__2888\ : InMux
    port map (
            O => \N__15012\,
            I => \N__14892\
        );

    \I__2887\ : InMux
    port map (
            O => \N__15011\,
            I => \N__14892\
        );

    \I__2886\ : InMux
    port map (
            O => \N__15010\,
            I => \N__14892\
        );

    \I__2885\ : InMux
    port map (
            O => \N__15009\,
            I => \N__14892\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__15006\,
            I => \N__14889\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__15001\,
            I => \N__14886\
        );

    \I__2882\ : InMux
    port map (
            O => \N__14998\,
            I => \N__14881\
        );

    \I__2881\ : InMux
    port map (
            O => \N__14997\,
            I => \N__14881\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__14994\,
            I => \N__14872\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__14989\,
            I => \N__14872\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__14984\,
            I => \N__14872\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__14979\,
            I => \N__14872\
        );

    \I__2876\ : InMux
    port map (
            O => \N__14978\,
            I => \N__14867\
        );

    \I__2875\ : InMux
    port map (
            O => \N__14977\,
            I => \N__14867\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__14974\,
            I => \N__14864\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__14965\,
            I => \N__14861\
        );

    \I__2872\ : InMux
    port map (
            O => \N__14964\,
            I => \N__14856\
        );

    \I__2871\ : InMux
    port map (
            O => \N__14963\,
            I => \N__14856\
        );

    \I__2870\ : InMux
    port map (
            O => \N__14962\,
            I => \N__14853\
        );

    \I__2869\ : InMux
    port map (
            O => \N__14961\,
            I => \N__14850\
        );

    \I__2868\ : InMux
    port map (
            O => \N__14960\,
            I => \N__14839\
        );

    \I__2867\ : InMux
    port map (
            O => \N__14959\,
            I => \N__14839\
        );

    \I__2866\ : InMux
    port map (
            O => \N__14958\,
            I => \N__14839\
        );

    \I__2865\ : InMux
    port map (
            O => \N__14957\,
            I => \N__14839\
        );

    \I__2864\ : InMux
    port map (
            O => \N__14956\,
            I => \N__14839\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__14953\,
            I => \N__14836\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__14950\,
            I => \N__14831\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__14947\,
            I => \N__14831\
        );

    \I__2860\ : InMux
    port map (
            O => \N__14946\,
            I => \N__14826\
        );

    \I__2859\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14826\
        );

    \I__2858\ : InMux
    port map (
            O => \N__14944\,
            I => \N__14823\
        );

    \I__2857\ : InMux
    port map (
            O => \N__14941\,
            I => \N__14818\
        );

    \I__2856\ : InMux
    port map (
            O => \N__14940\,
            I => \N__14818\
        );

    \I__2855\ : InMux
    port map (
            O => \N__14939\,
            I => \N__14811\
        );

    \I__2854\ : InMux
    port map (
            O => \N__14938\,
            I => \N__14811\
        );

    \I__2853\ : InMux
    port map (
            O => \N__14937\,
            I => \N__14811\
        );

    \I__2852\ : InMux
    port map (
            O => \N__14936\,
            I => \N__14804\
        );

    \I__2851\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14804\
        );

    \I__2850\ : InMux
    port map (
            O => \N__14934\,
            I => \N__14804\
        );

    \I__2849\ : InMux
    port map (
            O => \N__14933\,
            I => \N__14791\
        );

    \I__2848\ : InMux
    port map (
            O => \N__14932\,
            I => \N__14791\
        );

    \I__2847\ : InMux
    port map (
            O => \N__14931\,
            I => \N__14791\
        );

    \I__2846\ : InMux
    port map (
            O => \N__14930\,
            I => \N__14791\
        );

    \I__2845\ : InMux
    port map (
            O => \N__14929\,
            I => \N__14791\
        );

    \I__2844\ : InMux
    port map (
            O => \N__14928\,
            I => \N__14791\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__14919\,
            I => \N__14786\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__14914\,
            I => \N__14786\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__14901\,
            I => \N__14777\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__14892\,
            I => \N__14777\
        );

    \I__2839\ : Span4Mux_s2_v
    port map (
            O => \N__14889\,
            I => \N__14777\
        );

    \I__2838\ : Span4Mux_v
    port map (
            O => \N__14886\,
            I => \N__14777\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__14881\,
            I => \N__14772\
        );

    \I__2836\ : Span4Mux_h
    port map (
            O => \N__14872\,
            I => \N__14772\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__14867\,
            I => \N__14765\
        );

    \I__2834\ : Span4Mux_v
    port map (
            O => \N__14864\,
            I => \N__14765\
        );

    \I__2833\ : Span4Mux_h
    port map (
            O => \N__14861\,
            I => \N__14765\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__14856\,
            I => \N__14762\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__14853\,
            I => \N__14751\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__14850\,
            I => \N__14751\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__14839\,
            I => \N__14751\
        );

    \I__2828\ : Span4Mux_v
    port map (
            O => \N__14836\,
            I => \N__14751\
        );

    \I__2827\ : Span4Mux_h
    port map (
            O => \N__14831\,
            I => \N__14751\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__14826\,
            I => \c0.n1197\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__14823\,
            I => \c0.n1197\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__14818\,
            I => \c0.n1197\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__14811\,
            I => \c0.n1197\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__14804\,
            I => \c0.n1197\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__14791\,
            I => \c0.n1197\
        );

    \I__2820\ : Odrv12
    port map (
            O => \N__14786\,
            I => \c0.n1197\
        );

    \I__2819\ : Odrv4
    port map (
            O => \N__14777\,
            I => \c0.n1197\
        );

    \I__2818\ : Odrv4
    port map (
            O => \N__14772\,
            I => \c0.n1197\
        );

    \I__2817\ : Odrv4
    port map (
            O => \N__14765\,
            I => \c0.n1197\
        );

    \I__2816\ : Odrv12
    port map (
            O => \N__14762\,
            I => \c0.n1197\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__14751\,
            I => \c0.n1197\
        );

    \I__2814\ : CascadeMux
    port map (
            O => \N__14726\,
            I => \N__14717\
        );

    \I__2813\ : CascadeMux
    port map (
            O => \N__14725\,
            I => \N__14708\
        );

    \I__2812\ : CascadeMux
    port map (
            O => \N__14724\,
            I => \N__14699\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__14723\,
            I => \N__14696\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__14722\,
            I => \N__14690\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__14721\,
            I => \N__14681\
        );

    \I__2808\ : InMux
    port map (
            O => \N__14720\,
            I => \N__14674\
        );

    \I__2807\ : InMux
    port map (
            O => \N__14717\,
            I => \N__14674\
        );

    \I__2806\ : InMux
    port map (
            O => \N__14716\,
            I => \N__14674\
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__14715\,
            I => \N__14671\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__14714\,
            I => \N__14666\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__14713\,
            I => \N__14662\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__14712\,
            I => \N__14659\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__14711\,
            I => \N__14656\
        );

    \I__2800\ : InMux
    port map (
            O => \N__14708\,
            I => \N__14647\
        );

    \I__2799\ : InMux
    port map (
            O => \N__14707\,
            I => \N__14647\
        );

    \I__2798\ : CascadeMux
    port map (
            O => \N__14706\,
            I => \N__14636\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__14705\,
            I => \N__14633\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__14704\,
            I => \N__14630\
        );

    \I__2795\ : CascadeMux
    port map (
            O => \N__14703\,
            I => \N__14625\
        );

    \I__2794\ : CascadeMux
    port map (
            O => \N__14702\,
            I => \N__14622\
        );

    \I__2793\ : InMux
    port map (
            O => \N__14699\,
            I => \N__14612\
        );

    \I__2792\ : InMux
    port map (
            O => \N__14696\,
            I => \N__14612\
        );

    \I__2791\ : InMux
    port map (
            O => \N__14695\,
            I => \N__14612\
        );

    \I__2790\ : InMux
    port map (
            O => \N__14694\,
            I => \N__14612\
        );

    \I__2789\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14607\
        );

    \I__2788\ : InMux
    port map (
            O => \N__14690\,
            I => \N__14607\
        );

    \I__2787\ : InMux
    port map (
            O => \N__14689\,
            I => \N__14598\
        );

    \I__2786\ : InMux
    port map (
            O => \N__14688\,
            I => \N__14598\
        );

    \I__2785\ : InMux
    port map (
            O => \N__14687\,
            I => \N__14598\
        );

    \I__2784\ : InMux
    port map (
            O => \N__14686\,
            I => \N__14598\
        );

    \I__2783\ : CascadeMux
    port map (
            O => \N__14685\,
            I => \N__14595\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__14684\,
            I => \N__14592\
        );

    \I__2781\ : InMux
    port map (
            O => \N__14681\,
            I => \N__14586\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__14674\,
            I => \N__14583\
        );

    \I__2779\ : InMux
    port map (
            O => \N__14671\,
            I => \N__14580\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__14670\,
            I => \N__14575\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__14669\,
            I => \N__14571\
        );

    \I__2776\ : InMux
    port map (
            O => \N__14666\,
            I => \N__14567\
        );

    \I__2775\ : InMux
    port map (
            O => \N__14665\,
            I => \N__14562\
        );

    \I__2774\ : InMux
    port map (
            O => \N__14662\,
            I => \N__14562\
        );

    \I__2773\ : InMux
    port map (
            O => \N__14659\,
            I => \N__14555\
        );

    \I__2772\ : InMux
    port map (
            O => \N__14656\,
            I => \N__14555\
        );

    \I__2771\ : InMux
    port map (
            O => \N__14655\,
            I => \N__14555\
        );

    \I__2770\ : InMux
    port map (
            O => \N__14654\,
            I => \N__14548\
        );

    \I__2769\ : InMux
    port map (
            O => \N__14653\,
            I => \N__14548\
        );

    \I__2768\ : InMux
    port map (
            O => \N__14652\,
            I => \N__14548\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__14647\,
            I => \N__14545\
        );

    \I__2766\ : InMux
    port map (
            O => \N__14646\,
            I => \N__14542\
        );

    \I__2765\ : InMux
    port map (
            O => \N__14645\,
            I => \N__14531\
        );

    \I__2764\ : InMux
    port map (
            O => \N__14644\,
            I => \N__14531\
        );

    \I__2763\ : InMux
    port map (
            O => \N__14643\,
            I => \N__14531\
        );

    \I__2762\ : InMux
    port map (
            O => \N__14642\,
            I => \N__14531\
        );

    \I__2761\ : InMux
    port map (
            O => \N__14641\,
            I => \N__14531\
        );

    \I__2760\ : InMux
    port map (
            O => \N__14640\,
            I => \N__14518\
        );

    \I__2759\ : InMux
    port map (
            O => \N__14639\,
            I => \N__14518\
        );

    \I__2758\ : InMux
    port map (
            O => \N__14636\,
            I => \N__14518\
        );

    \I__2757\ : InMux
    port map (
            O => \N__14633\,
            I => \N__14518\
        );

    \I__2756\ : InMux
    port map (
            O => \N__14630\,
            I => \N__14518\
        );

    \I__2755\ : InMux
    port map (
            O => \N__14629\,
            I => \N__14518\
        );

    \I__2754\ : InMux
    port map (
            O => \N__14628\,
            I => \N__14509\
        );

    \I__2753\ : InMux
    port map (
            O => \N__14625\,
            I => \N__14509\
        );

    \I__2752\ : InMux
    port map (
            O => \N__14622\,
            I => \N__14509\
        );

    \I__2751\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14509\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__14612\,
            I => \N__14502\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__14607\,
            I => \N__14502\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__14598\,
            I => \N__14502\
        );

    \I__2747\ : InMux
    port map (
            O => \N__14595\,
            I => \N__14496\
        );

    \I__2746\ : InMux
    port map (
            O => \N__14592\,
            I => \N__14496\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__14591\,
            I => \N__14490\
        );

    \I__2744\ : CascadeMux
    port map (
            O => \N__14590\,
            I => \N__14487\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__14589\,
            I => \N__14481\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__14586\,
            I => \N__14474\
        );

    \I__2741\ : Span4Mux_s3_v
    port map (
            O => \N__14583\,
            I => \N__14474\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__14580\,
            I => \N__14474\
        );

    \I__2739\ : CascadeMux
    port map (
            O => \N__14579\,
            I => \N__14469\
        );

    \I__2738\ : CascadeMux
    port map (
            O => \N__14578\,
            I => \N__14466\
        );

    \I__2737\ : InMux
    port map (
            O => \N__14575\,
            I => \N__14459\
        );

    \I__2736\ : InMux
    port map (
            O => \N__14574\,
            I => \N__14459\
        );

    \I__2735\ : InMux
    port map (
            O => \N__14571\,
            I => \N__14454\
        );

    \I__2734\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14454\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__14567\,
            I => \N__14451\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__14562\,
            I => \N__14432\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__14555\,
            I => \N__14432\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__14548\,
            I => \N__14432\
        );

    \I__2729\ : Span4Mux_s2_h
    port map (
            O => \N__14545\,
            I => \N__14432\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__14542\,
            I => \N__14432\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__14531\,
            I => \N__14432\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__14518\,
            I => \N__14432\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__14509\,
            I => \N__14432\
        );

    \I__2724\ : Span4Mux_s3_v
    port map (
            O => \N__14502\,
            I => \N__14432\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__14501\,
            I => \N__14429\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__14496\,
            I => \N__14425\
        );

    \I__2721\ : InMux
    port map (
            O => \N__14495\,
            I => \N__14420\
        );

    \I__2720\ : InMux
    port map (
            O => \N__14494\,
            I => \N__14420\
        );

    \I__2719\ : InMux
    port map (
            O => \N__14493\,
            I => \N__14407\
        );

    \I__2718\ : InMux
    port map (
            O => \N__14490\,
            I => \N__14407\
        );

    \I__2717\ : InMux
    port map (
            O => \N__14487\,
            I => \N__14407\
        );

    \I__2716\ : InMux
    port map (
            O => \N__14486\,
            I => \N__14407\
        );

    \I__2715\ : InMux
    port map (
            O => \N__14485\,
            I => \N__14407\
        );

    \I__2714\ : InMux
    port map (
            O => \N__14484\,
            I => \N__14407\
        );

    \I__2713\ : InMux
    port map (
            O => \N__14481\,
            I => \N__14401\
        );

    \I__2712\ : Span4Mux_v
    port map (
            O => \N__14474\,
            I => \N__14398\
        );

    \I__2711\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14389\
        );

    \I__2710\ : InMux
    port map (
            O => \N__14472\,
            I => \N__14389\
        );

    \I__2709\ : InMux
    port map (
            O => \N__14469\,
            I => \N__14389\
        );

    \I__2708\ : InMux
    port map (
            O => \N__14466\,
            I => \N__14389\
        );

    \I__2707\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14384\
        );

    \I__2706\ : InMux
    port map (
            O => \N__14464\,
            I => \N__14384\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__14459\,
            I => \N__14381\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__14454\,
            I => \N__14376\
        );

    \I__2703\ : Span4Mux_s3_h
    port map (
            O => \N__14451\,
            I => \N__14376\
        );

    \I__2702\ : Span4Mux_v
    port map (
            O => \N__14432\,
            I => \N__14373\
        );

    \I__2701\ : InMux
    port map (
            O => \N__14429\,
            I => \N__14370\
        );

    \I__2700\ : InMux
    port map (
            O => \N__14428\,
            I => \N__14367\
        );

    \I__2699\ : Span4Mux_v
    port map (
            O => \N__14425\,
            I => \N__14362\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__14420\,
            I => \N__14362\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__14407\,
            I => \N__14359\
        );

    \I__2696\ : InMux
    port map (
            O => \N__14406\,
            I => \N__14354\
        );

    \I__2695\ : InMux
    port map (
            O => \N__14405\,
            I => \N__14354\
        );

    \I__2694\ : InMux
    port map (
            O => \N__14404\,
            I => \N__14351\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__14401\,
            I => \N__14346\
        );

    \I__2692\ : Span4Mux_s0_h
    port map (
            O => \N__14398\,
            I => \N__14346\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__14389\,
            I => \N__14337\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__14384\,
            I => \N__14337\
        );

    \I__2689\ : Span4Mux_s3_h
    port map (
            O => \N__14381\,
            I => \N__14337\
        );

    \I__2688\ : Span4Mux_v
    port map (
            O => \N__14376\,
            I => \N__14337\
        );

    \I__2687\ : Span4Mux_s2_h
    port map (
            O => \N__14373\,
            I => \N__14334\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__14370\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__14367\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__14362\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__2683\ : Odrv12
    port map (
            O => \N__14359\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__14354\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__14351\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__14346\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__14337\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__14334\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__2677\ : InMux
    port map (
            O => \N__14315\,
            I => \N__14312\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__14312\,
            I => \N__14307\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__14311\,
            I => \N__14304\
        );

    \I__2674\ : InMux
    port map (
            O => \N__14310\,
            I => \N__14301\
        );

    \I__2673\ : Span4Mux_v
    port map (
            O => \N__14307\,
            I => \N__14298\
        );

    \I__2672\ : InMux
    port map (
            O => \N__14304\,
            I => \N__14295\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__14301\,
            I => \c0.data_in_field_10\
        );

    \I__2670\ : Odrv4
    port map (
            O => \N__14298\,
            I => \c0.data_in_field_10\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__14295\,
            I => \c0.data_in_field_10\
        );

    \I__2668\ : InMux
    port map (
            O => \N__14288\,
            I => \N__14284\
        );

    \I__2667\ : InMux
    port map (
            O => \N__14287\,
            I => \N__14281\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__14284\,
            I => n2651
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__14281\,
            I => n2651
        );

    \I__2664\ : CascadeMux
    port map (
            O => \N__14276\,
            I => \N__14273\
        );

    \I__2663\ : InMux
    port map (
            O => \N__14273\,
            I => \N__14268\
        );

    \I__2662\ : InMux
    port map (
            O => \N__14272\,
            I => \N__14265\
        );

    \I__2661\ : InMux
    port map (
            O => \N__14271\,
            I => \N__14262\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__14268\,
            I => data_in_5_0
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__14265\,
            I => data_in_5_0
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__14262\,
            I => data_in_5_0
        );

    \I__2657\ : InMux
    port map (
            O => \N__14255\,
            I => \N__14251\
        );

    \I__2656\ : InMux
    port map (
            O => \N__14254\,
            I => \N__14248\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__14251\,
            I => \N__14242\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__14248\,
            I => \N__14242\
        );

    \I__2653\ : InMux
    port map (
            O => \N__14247\,
            I => \N__14239\
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__14242\,
            I => data_in_4_0
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__14239\,
            I => data_in_4_0
        );

    \I__2650\ : InMux
    port map (
            O => \N__14234\,
            I => \N__14231\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__14231\,
            I => \N__14228\
        );

    \I__2648\ : Span4Mux_h
    port map (
            O => \N__14228\,
            I => \N__14223\
        );

    \I__2647\ : InMux
    port map (
            O => \N__14227\,
            I => \N__14220\
        );

    \I__2646\ : InMux
    port map (
            O => \N__14226\,
            I => \N__14217\
        );

    \I__2645\ : Odrv4
    port map (
            O => \N__14223\,
            I => data_in_4_3
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__14220\,
            I => data_in_4_3
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__14217\,
            I => data_in_4_3
        );

    \I__2642\ : InMux
    port map (
            O => \N__14210\,
            I => \N__14206\
        );

    \I__2641\ : InMux
    port map (
            O => \N__14209\,
            I => \N__14203\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__14206\,
            I => \N__14198\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__14203\,
            I => \N__14195\
        );

    \I__2638\ : InMux
    port map (
            O => \N__14202\,
            I => \N__14192\
        );

    \I__2637\ : InMux
    port map (
            O => \N__14201\,
            I => \N__14189\
        );

    \I__2636\ : Span4Mux_v
    port map (
            O => \N__14198\,
            I => \N__14182\
        );

    \I__2635\ : Span4Mux_s2_v
    port map (
            O => \N__14195\,
            I => \N__14182\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__14192\,
            I => \N__14182\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__14189\,
            I => data_in_3_3
        );

    \I__2632\ : Odrv4
    port map (
            O => \N__14182\,
            I => data_in_3_3
        );

    \I__2631\ : CascadeMux
    port map (
            O => \N__14177\,
            I => \N__14174\
        );

    \I__2630\ : InMux
    port map (
            O => \N__14174\,
            I => \N__14170\
        );

    \I__2629\ : InMux
    port map (
            O => \N__14173\,
            I => \N__14167\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__14170\,
            I => \N__14162\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__14167\,
            I => \N__14162\
        );

    \I__2626\ : Span4Mux_v
    port map (
            O => \N__14162\,
            I => \N__14158\
        );

    \I__2625\ : InMux
    port map (
            O => \N__14161\,
            I => \N__14155\
        );

    \I__2624\ : Odrv4
    port map (
            O => \N__14158\,
            I => data_in_5_2
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__14155\,
            I => data_in_5_2
        );

    \I__2622\ : InMux
    port map (
            O => \N__14150\,
            I => \N__14146\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__14149\,
            I => \N__14143\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__14146\,
            I => \N__14139\
        );

    \I__2619\ : InMux
    port map (
            O => \N__14143\,
            I => \N__14134\
        );

    \I__2618\ : InMux
    port map (
            O => \N__14142\,
            I => \N__14134\
        );

    \I__2617\ : Odrv12
    port map (
            O => \N__14139\,
            I => n1222
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__14134\,
            I => n1222
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__14129\,
            I => \N__14125\
        );

    \I__2614\ : InMux
    port map (
            O => \N__14128\,
            I => \N__14122\
        );

    \I__2613\ : InMux
    port map (
            O => \N__14125\,
            I => \N__14119\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__14122\,
            I => \N__14115\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__14119\,
            I => \N__14111\
        );

    \I__2610\ : InMux
    port map (
            O => \N__14118\,
            I => \N__14108\
        );

    \I__2609\ : Span4Mux_h
    port map (
            O => \N__14115\,
            I => \N__14105\
        );

    \I__2608\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14102\
        );

    \I__2607\ : Span4Mux_h
    port map (
            O => \N__14111\,
            I => \N__14099\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__14108\,
            I => data_in_7_3
        );

    \I__2605\ : Odrv4
    port map (
            O => \N__14105\,
            I => data_in_7_3
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__14102\,
            I => data_in_7_3
        );

    \I__2603\ : Odrv4
    port map (
            O => \N__14099\,
            I => data_in_7_3
        );

    \I__2602\ : InMux
    port map (
            O => \N__14090\,
            I => \N__14087\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__14087\,
            I => \N__14081\
        );

    \I__2600\ : InMux
    port map (
            O => \N__14086\,
            I => \N__14078\
        );

    \I__2599\ : InMux
    port map (
            O => \N__14085\,
            I => \N__14073\
        );

    \I__2598\ : InMux
    port map (
            O => \N__14084\,
            I => \N__14073\
        );

    \I__2597\ : Span4Mux_v
    port map (
            O => \N__14081\,
            I => \N__14070\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__14078\,
            I => \N__14067\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__14073\,
            I => data_in_7_6
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__14070\,
            I => data_in_7_6
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__14067\,
            I => data_in_7_6
        );

    \I__2592\ : IoInMux
    port map (
            O => \N__14060\,
            I => \N__14057\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__14057\,
            I => \N__14053\
        );

    \I__2590\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14050\
        );

    \I__2589\ : Span4Mux_s3_h
    port map (
            O => \N__14053\,
            I => \N__14046\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__14050\,
            I => \N__14043\
        );

    \I__2587\ : InMux
    port map (
            O => \N__14049\,
            I => \N__14040\
        );

    \I__2586\ : Odrv4
    port map (
            O => \N__14046\,
            I => tx2_o_adj_949
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__14043\,
            I => tx2_o_adj_949
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__14040\,
            I => tx2_o_adj_949
        );

    \I__2583\ : IoInMux
    port map (
            O => \N__14033\,
            I => \N__14030\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__14030\,
            I => \N__14027\
        );

    \I__2581\ : Span4Mux_s0_h
    port map (
            O => \N__14027\,
            I => \N__14024\
        );

    \I__2580\ : Span4Mux_h
    port map (
            O => \N__14024\,
            I => \N__14021\
        );

    \I__2579\ : Odrv4
    port map (
            O => \N__14021\,
            I => tx2_enable
        );

    \I__2578\ : InMux
    port map (
            O => \N__14018\,
            I => \N__14015\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__14015\,
            I => \N__14009\
        );

    \I__2576\ : CascadeMux
    port map (
            O => \N__14014\,
            I => \N__14006\
        );

    \I__2575\ : InMux
    port map (
            O => \N__14013\,
            I => \N__14002\
        );

    \I__2574\ : InMux
    port map (
            O => \N__14012\,
            I => \N__13999\
        );

    \I__2573\ : Span12Mux_h
    port map (
            O => \N__14009\,
            I => \N__13996\
        );

    \I__2572\ : InMux
    port map (
            O => \N__14006\,
            I => \N__13993\
        );

    \I__2571\ : InMux
    port map (
            O => \N__14005\,
            I => \N__13990\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__14002\,
            I => \N__13987\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__13999\,
            I => \c0.data_in_field_12\
        );

    \I__2568\ : Odrv12
    port map (
            O => \N__13996\,
            I => \c0.data_in_field_12\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__13993\,
            I => \c0.data_in_field_12\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__13990\,
            I => \c0.data_in_field_12\
        );

    \I__2565\ : Odrv12
    port map (
            O => \N__13987\,
            I => \c0.data_in_field_12\
        );

    \I__2564\ : InMux
    port map (
            O => \N__13976\,
            I => \N__13973\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__13973\,
            I => \N__13968\
        );

    \I__2562\ : InMux
    port map (
            O => \N__13972\,
            I => \N__13965\
        );

    \I__2561\ : InMux
    port map (
            O => \N__13971\,
            I => \N__13960\
        );

    \I__2560\ : Sp12to4
    port map (
            O => \N__13968\,
            I => \N__13955\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__13965\,
            I => \N__13955\
        );

    \I__2558\ : InMux
    port map (
            O => \N__13964\,
            I => \N__13952\
        );

    \I__2557\ : InMux
    port map (
            O => \N__13963\,
            I => \N__13949\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__13960\,
            I => \c0.data_in_field_40\
        );

    \I__2555\ : Odrv12
    port map (
            O => \N__13955\,
            I => \c0.data_in_field_40\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__13952\,
            I => \c0.data_in_field_40\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__13949\,
            I => \c0.data_in_field_40\
        );

    \I__2552\ : InMux
    port map (
            O => \N__13940\,
            I => \N__13936\
        );

    \I__2551\ : InMux
    port map (
            O => \N__13939\,
            I => \N__13932\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__13936\,
            I => \N__13929\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__13935\,
            I => \N__13925\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__13932\,
            I => \N__13922\
        );

    \I__2547\ : Span4Mux_h
    port map (
            O => \N__13929\,
            I => \N__13919\
        );

    \I__2546\ : InMux
    port map (
            O => \N__13928\,
            I => \N__13914\
        );

    \I__2545\ : InMux
    port map (
            O => \N__13925\,
            I => \N__13914\
        );

    \I__2544\ : Odrv12
    port map (
            O => \N__13922\,
            I => data_in_6_6
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__13919\,
            I => data_in_6_6
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__13914\,
            I => data_in_6_6
        );

    \I__2541\ : CascadeMux
    port map (
            O => \N__13907\,
            I => \N__13903\
        );

    \I__2540\ : InMux
    port map (
            O => \N__13906\,
            I => \N__13900\
        );

    \I__2539\ : InMux
    port map (
            O => \N__13903\,
            I => \N__13897\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__13900\,
            I => \N__13890\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__13897\,
            I => \N__13890\
        );

    \I__2536\ : InMux
    port map (
            O => \N__13896\,
            I => \N__13887\
        );

    \I__2535\ : InMux
    port map (
            O => \N__13895\,
            I => \N__13883\
        );

    \I__2534\ : Span4Mux_h
    port map (
            O => \N__13890\,
            I => \N__13880\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__13887\,
            I => \N__13877\
        );

    \I__2532\ : InMux
    port map (
            O => \N__13886\,
            I => \N__13874\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__13883\,
            I => \c0.data_in_field_41\
        );

    \I__2530\ : Odrv4
    port map (
            O => \N__13880\,
            I => \c0.data_in_field_41\
        );

    \I__2529\ : Odrv12
    port map (
            O => \N__13877\,
            I => \c0.data_in_field_41\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__13874\,
            I => \c0.data_in_field_41\
        );

    \I__2527\ : InMux
    port map (
            O => \N__13865\,
            I => \N__13862\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__13862\,
            I => \N__13859\
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__13859\,
            I => \c0.n12_adj_878\
        );

    \I__2524\ : InMux
    port map (
            O => \N__13856\,
            I => \N__13853\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__13853\,
            I => \N__13849\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__13852\,
            I => \N__13846\
        );

    \I__2521\ : Span4Mux_h
    port map (
            O => \N__13849\,
            I => \N__13843\
        );

    \I__2520\ : InMux
    port map (
            O => \N__13846\,
            I => \N__13840\
        );

    \I__2519\ : Odrv4
    port map (
            O => \N__13843\,
            I => rx_data_4
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__13840\,
            I => rx_data_4
        );

    \I__2517\ : InMux
    port map (
            O => \N__13835\,
            I => \N__13832\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__13832\,
            I => \N__13828\
        );

    \I__2515\ : CascadeMux
    port map (
            O => \N__13831\,
            I => \N__13825\
        );

    \I__2514\ : Span4Mux_h
    port map (
            O => \N__13828\,
            I => \N__13822\
        );

    \I__2513\ : InMux
    port map (
            O => \N__13825\,
            I => \N__13817\
        );

    \I__2512\ : Span4Mux_v
    port map (
            O => \N__13822\,
            I => \N__13814\
        );

    \I__2511\ : InMux
    port map (
            O => \N__13821\,
            I => \N__13811\
        );

    \I__2510\ : InMux
    port map (
            O => \N__13820\,
            I => \N__13808\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__13817\,
            I => \N__13805\
        );

    \I__2508\ : Odrv4
    port map (
            O => \N__13814\,
            I => data_in_7_4
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__13811\,
            I => data_in_7_4
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__13808\,
            I => data_in_7_4
        );

    \I__2505\ : Odrv4
    port map (
            O => \N__13805\,
            I => data_in_7_4
        );

    \I__2504\ : InMux
    port map (
            O => \N__13796\,
            I => \N__13793\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__13793\,
            I => \N__13789\
        );

    \I__2502\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13786\
        );

    \I__2501\ : Span4Mux_h
    port map (
            O => \N__13789\,
            I => \N__13781\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__13786\,
            I => \N__13778\
        );

    \I__2499\ : InMux
    port map (
            O => \N__13785\,
            I => \N__13775\
        );

    \I__2498\ : InMux
    port map (
            O => \N__13784\,
            I => \N__13772\
        );

    \I__2497\ : Odrv4
    port map (
            O => \N__13781\,
            I => data_in_3_0
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__13778\,
            I => data_in_3_0
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__13775\,
            I => data_in_3_0
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__13772\,
            I => data_in_3_0
        );

    \I__2493\ : InMux
    port map (
            O => \N__13763\,
            I => \N__13760\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__13760\,
            I => \N__13756\
        );

    \I__2491\ : InMux
    port map (
            O => \N__13759\,
            I => \N__13753\
        );

    \I__2490\ : Span4Mux_v
    port map (
            O => \N__13756\,
            I => \N__13746\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__13753\,
            I => \N__13746\
        );

    \I__2488\ : InMux
    port map (
            O => \N__13752\,
            I => \N__13743\
        );

    \I__2487\ : InMux
    port map (
            O => \N__13751\,
            I => \N__13739\
        );

    \I__2486\ : Span4Mux_h
    port map (
            O => \N__13746\,
            I => \N__13734\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__13743\,
            I => \N__13734\
        );

    \I__2484\ : InMux
    port map (
            O => \N__13742\,
            I => \N__13731\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__13739\,
            I => \c0.data_in_field_24\
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__13734\,
            I => \c0.data_in_field_24\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__13731\,
            I => \c0.data_in_field_24\
        );

    \I__2480\ : InMux
    port map (
            O => \N__13724\,
            I => \N__13719\
        );

    \I__2479\ : InMux
    port map (
            O => \N__13723\,
            I => \N__13716\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__13722\,
            I => \N__13713\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__13719\,
            I => \N__13709\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__13716\,
            I => \N__13706\
        );

    \I__2475\ : InMux
    port map (
            O => \N__13713\,
            I => \N__13703\
        );

    \I__2474\ : InMux
    port map (
            O => \N__13712\,
            I => \N__13700\
        );

    \I__2473\ : Span4Mux_v
    port map (
            O => \N__13709\,
            I => \N__13697\
        );

    \I__2472\ : Span4Mux_v
    port map (
            O => \N__13706\,
            I => \N__13692\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__13703\,
            I => \N__13692\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__13700\,
            I => data_in_7_7
        );

    \I__2469\ : Odrv4
    port map (
            O => \N__13697\,
            I => data_in_7_7
        );

    \I__2468\ : Odrv4
    port map (
            O => \N__13692\,
            I => data_in_7_7
        );

    \I__2467\ : InMux
    port map (
            O => \N__13685\,
            I => \N__13682\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__13682\,
            I => \N__13678\
        );

    \I__2465\ : InMux
    port map (
            O => \N__13681\,
            I => \N__13675\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__13678\,
            I => \N__13670\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__13675\,
            I => \N__13667\
        );

    \I__2462\ : InMux
    port map (
            O => \N__13674\,
            I => \N__13664\
        );

    \I__2461\ : InMux
    port map (
            O => \N__13673\,
            I => \N__13661\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__13670\,
            I => data_in_6_7
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__13667\,
            I => data_in_6_7
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__13664\,
            I => data_in_6_7
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__13661\,
            I => data_in_6_7
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__13652\,
            I => \N__13649\
        );

    \I__2455\ : InMux
    port map (
            O => \N__13649\,
            I => \N__13646\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__13646\,
            I => \N__13640\
        );

    \I__2453\ : InMux
    port map (
            O => \N__13645\,
            I => \N__13637\
        );

    \I__2452\ : InMux
    port map (
            O => \N__13644\,
            I => \N__13631\
        );

    \I__2451\ : InMux
    port map (
            O => \N__13643\,
            I => \N__13631\
        );

    \I__2450\ : Span4Mux_h
    port map (
            O => \N__13640\,
            I => \N__13628\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__13637\,
            I => \N__13625\
        );

    \I__2448\ : InMux
    port map (
            O => \N__13636\,
            I => \N__13622\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__13631\,
            I => \c0.data_in_field_35\
        );

    \I__2446\ : Odrv4
    port map (
            O => \N__13628\,
            I => \c0.data_in_field_35\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__13625\,
            I => \c0.data_in_field_35\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__13622\,
            I => \c0.data_in_field_35\
        );

    \I__2443\ : InMux
    port map (
            O => \N__13613\,
            I => \N__13609\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__13612\,
            I => \N__13605\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__13609\,
            I => \N__13602\
        );

    \I__2440\ : InMux
    port map (
            O => \N__13608\,
            I => \N__13599\
        );

    \I__2439\ : InMux
    port map (
            O => \N__13605\,
            I => \N__13594\
        );

    \I__2438\ : Span4Mux_v
    port map (
            O => \N__13602\,
            I => \N__13591\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__13599\,
            I => \N__13588\
        );

    \I__2436\ : InMux
    port map (
            O => \N__13598\,
            I => \N__13585\
        );

    \I__2435\ : InMux
    port map (
            O => \N__13597\,
            I => \N__13582\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__13594\,
            I => \c0.data_in_field_36\
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__13591\,
            I => \c0.data_in_field_36\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__13588\,
            I => \c0.data_in_field_36\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__13585\,
            I => \c0.data_in_field_36\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__13582\,
            I => \c0.data_in_field_36\
        );

    \I__2429\ : InMux
    port map (
            O => \N__13571\,
            I => \N__13568\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__13568\,
            I => \c0.n11\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__13565\,
            I => \N__13562\
        );

    \I__2426\ : InMux
    port map (
            O => \N__13562\,
            I => \N__13559\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__13559\,
            I => \N__13555\
        );

    \I__2424\ : InMux
    port map (
            O => \N__13558\,
            I => \N__13550\
        );

    \I__2423\ : Span4Mux_h
    port map (
            O => \N__13555\,
            I => \N__13547\
        );

    \I__2422\ : InMux
    port map (
            O => \N__13554\,
            I => \N__13542\
        );

    \I__2421\ : InMux
    port map (
            O => \N__13553\,
            I => \N__13542\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__13550\,
            I => \c0.data_in_field_43\
        );

    \I__2419\ : Odrv4
    port map (
            O => \N__13547\,
            I => \c0.data_in_field_43\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__13542\,
            I => \c0.data_in_field_43\
        );

    \I__2417\ : InMux
    port map (
            O => \N__13535\,
            I => \N__13532\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__13532\,
            I => \N__13527\
        );

    \I__2415\ : InMux
    port map (
            O => \N__13531\,
            I => \N__13522\
        );

    \I__2414\ : InMux
    port map (
            O => \N__13530\,
            I => \N__13519\
        );

    \I__2413\ : Span4Mux_h
    port map (
            O => \N__13527\,
            I => \N__13516\
        );

    \I__2412\ : InMux
    port map (
            O => \N__13526\,
            I => \N__13513\
        );

    \I__2411\ : InMux
    port map (
            O => \N__13525\,
            I => \N__13510\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__13522\,
            I => \c0.data_in_field_26\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__13519\,
            I => \c0.data_in_field_26\
        );

    \I__2408\ : Odrv4
    port map (
            O => \N__13516\,
            I => \c0.data_in_field_26\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__13513\,
            I => \c0.data_in_field_26\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__13510\,
            I => \c0.data_in_field_26\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__13499\,
            I => \c0.n4415_cascade_\
        );

    \I__2404\ : InMux
    port map (
            O => \N__13496\,
            I => \N__13492\
        );

    \I__2403\ : InMux
    port map (
            O => \N__13495\,
            I => \N__13489\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__13492\,
            I => \N__13486\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__13489\,
            I => \N__13482\
        );

    \I__2400\ : Span4Mux_v
    port map (
            O => \N__13486\,
            I => \N__13477\
        );

    \I__2399\ : InMux
    port map (
            O => \N__13485\,
            I => \N__13474\
        );

    \I__2398\ : Span4Mux_s3_h
    port map (
            O => \N__13482\,
            I => \N__13471\
        );

    \I__2397\ : InMux
    port map (
            O => \N__13481\,
            I => \N__13466\
        );

    \I__2396\ : InMux
    port map (
            O => \N__13480\,
            I => \N__13466\
        );

    \I__2395\ : Odrv4
    port map (
            O => \N__13477\,
            I => \c0.data_in_field_9\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__13474\,
            I => \c0.data_in_field_9\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__13471\,
            I => \c0.data_in_field_9\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__13466\,
            I => \c0.data_in_field_9\
        );

    \I__2391\ : InMux
    port map (
            O => \N__13457\,
            I => \N__13454\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__13454\,
            I => \N__13451\
        );

    \I__2389\ : Odrv4
    port map (
            O => \N__13451\,
            I => \c0.n23\
        );

    \I__2388\ : InMux
    port map (
            O => \N__13448\,
            I => \N__13444\
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__13447\,
            I => \N__13440\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__13444\,
            I => \N__13437\
        );

    \I__2385\ : InMux
    port map (
            O => \N__13443\,
            I => \N__13434\
        );

    \I__2384\ : InMux
    port map (
            O => \N__13440\,
            I => \N__13429\
        );

    \I__2383\ : Span4Mux_v
    port map (
            O => \N__13437\,
            I => \N__13426\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__13434\,
            I => \N__13423\
        );

    \I__2381\ : InMux
    port map (
            O => \N__13433\,
            I => \N__13420\
        );

    \I__2380\ : InMux
    port map (
            O => \N__13432\,
            I => \N__13417\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__13429\,
            I => \c0.data_in_field_30\
        );

    \I__2378\ : Odrv4
    port map (
            O => \N__13426\,
            I => \c0.data_in_field_30\
        );

    \I__2377\ : Odrv4
    port map (
            O => \N__13423\,
            I => \c0.data_in_field_30\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__13420\,
            I => \c0.data_in_field_30\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__13417\,
            I => \c0.data_in_field_30\
        );

    \I__2374\ : InMux
    port map (
            O => \N__13406\,
            I => \N__13403\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__13403\,
            I => \N__13400\
        );

    \I__2372\ : Span4Mux_h
    port map (
            O => \N__13400\,
            I => \N__13397\
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__13397\,
            I => \c0.n4927\
        );

    \I__2370\ : InMux
    port map (
            O => \N__13394\,
            I => \N__13390\
        );

    \I__2369\ : InMux
    port map (
            O => \N__13393\,
            I => \N__13387\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__13390\,
            I => \c0.n1267\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__13387\,
            I => \c0.n1267\
        );

    \I__2366\ : InMux
    port map (
            O => \N__13382\,
            I => \N__13379\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__13379\,
            I => \c0.n4421\
        );

    \I__2364\ : InMux
    port map (
            O => \N__13376\,
            I => \N__13373\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__13373\,
            I => \N__13370\
        );

    \I__2362\ : Span4Mux_s3_h
    port map (
            O => \N__13370\,
            I => \N__13363\
        );

    \I__2361\ : InMux
    port map (
            O => \N__13369\,
            I => \N__13360\
        );

    \I__2360\ : InMux
    port map (
            O => \N__13368\,
            I => \N__13357\
        );

    \I__2359\ : InMux
    port map (
            O => \N__13367\,
            I => \N__13352\
        );

    \I__2358\ : InMux
    port map (
            O => \N__13366\,
            I => \N__13352\
        );

    \I__2357\ : Odrv4
    port map (
            O => \N__13363\,
            I => \c0.data_in_field_23\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__13360\,
            I => \c0.data_in_field_23\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__13357\,
            I => \c0.data_in_field_23\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__13352\,
            I => \c0.data_in_field_23\
        );

    \I__2353\ : InMux
    port map (
            O => \N__13343\,
            I => \N__13338\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__13342\,
            I => \N__13335\
        );

    \I__2351\ : InMux
    port map (
            O => \N__13341\,
            I => \N__13332\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__13338\,
            I => \N__13329\
        );

    \I__2349\ : InMux
    port map (
            O => \N__13335\,
            I => \N__13324\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__13332\,
            I => \N__13321\
        );

    \I__2347\ : Span4Mux_h
    port map (
            O => \N__13329\,
            I => \N__13318\
        );

    \I__2346\ : InMux
    port map (
            O => \N__13328\,
            I => \N__13313\
        );

    \I__2345\ : InMux
    port map (
            O => \N__13327\,
            I => \N__13313\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__13324\,
            I => \c0.data_in_field_37\
        );

    \I__2343\ : Odrv12
    port map (
            O => \N__13321\,
            I => \c0.data_in_field_37\
        );

    \I__2342\ : Odrv4
    port map (
            O => \N__13318\,
            I => \c0.data_in_field_37\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__13313\,
            I => \c0.data_in_field_37\
        );

    \I__2340\ : InMux
    port map (
            O => \N__13304\,
            I => \N__13301\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__13301\,
            I => \c0.n8_adj_883\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__13298\,
            I => \N__13294\
        );

    \I__2337\ : InMux
    port map (
            O => \N__13297\,
            I => \N__13290\
        );

    \I__2336\ : InMux
    port map (
            O => \N__13294\,
            I => \N__13285\
        );

    \I__2335\ : InMux
    port map (
            O => \N__13293\,
            I => \N__13285\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__13290\,
            I => \N__13280\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__13285\,
            I => \N__13277\
        );

    \I__2332\ : InMux
    port map (
            O => \N__13284\,
            I => \N__13272\
        );

    \I__2331\ : InMux
    port map (
            O => \N__13283\,
            I => \N__13272\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__13280\,
            I => \c0.data_in_field_25\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__13277\,
            I => \c0.data_in_field_25\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__13272\,
            I => \c0.data_in_field_25\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__13265\,
            I => \N__13260\
        );

    \I__2326\ : InMux
    port map (
            O => \N__13264\,
            I => \N__13257\
        );

    \I__2325\ : InMux
    port map (
            O => \N__13263\,
            I => \N__13254\
        );

    \I__2324\ : InMux
    port map (
            O => \N__13260\,
            I => \N__13251\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__13257\,
            I => \N__13242\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__13254\,
            I => \N__13242\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__13251\,
            I => \N__13242\
        );

    \I__2320\ : InMux
    port map (
            O => \N__13250\,
            I => \N__13237\
        );

    \I__2319\ : InMux
    port map (
            O => \N__13249\,
            I => \N__13237\
        );

    \I__2318\ : Odrv4
    port map (
            O => \N__13242\,
            I => \c0.n1290\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__13237\,
            I => \c0.n1290\
        );

    \I__2316\ : InMux
    port map (
            O => \N__13232\,
            I => \N__13229\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__13226\,
            I => \c0.n4441\
        );

    \I__2313\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13218\
        );

    \I__2312\ : InMux
    port map (
            O => \N__13222\,
            I => \N__13215\
        );

    \I__2311\ : InMux
    port map (
            O => \N__13221\,
            I => \N__13211\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__13218\,
            I => \N__13208\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__13215\,
            I => \N__13205\
        );

    \I__2308\ : InMux
    port map (
            O => \N__13214\,
            I => \N__13202\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__13211\,
            I => \c0.data_in_field_28\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__13208\,
            I => \c0.data_in_field_28\
        );

    \I__2305\ : Odrv4
    port map (
            O => \N__13205\,
            I => \c0.data_in_field_28\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__13202\,
            I => \c0.data_in_field_28\
        );

    \I__2303\ : InMux
    port map (
            O => \N__13193\,
            I => \N__13190\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__13190\,
            I => \N__13186\
        );

    \I__2301\ : InMux
    port map (
            O => \N__13189\,
            I => \N__13179\
        );

    \I__2300\ : Span4Mux_v
    port map (
            O => \N__13186\,
            I => \N__13176\
        );

    \I__2299\ : InMux
    port map (
            O => \N__13185\,
            I => \N__13173\
        );

    \I__2298\ : InMux
    port map (
            O => \N__13184\,
            I => \N__13170\
        );

    \I__2297\ : InMux
    port map (
            O => \N__13183\,
            I => \N__13167\
        );

    \I__2296\ : InMux
    port map (
            O => \N__13182\,
            I => \N__13164\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__13179\,
            I => \c0.data_in_field_42\
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__13176\,
            I => \c0.data_in_field_42\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__13173\,
            I => \c0.data_in_field_42\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__13170\,
            I => \c0.data_in_field_42\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__13167\,
            I => \c0.data_in_field_42\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__13164\,
            I => \c0.data_in_field_42\
        );

    \I__2289\ : InMux
    port map (
            O => \N__13151\,
            I => \N__13148\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__13148\,
            I => \N__13142\
        );

    \I__2287\ : InMux
    port map (
            O => \N__13147\,
            I => \N__13139\
        );

    \I__2286\ : InMux
    port map (
            O => \N__13146\,
            I => \N__13134\
        );

    \I__2285\ : InMux
    port map (
            O => \N__13145\,
            I => \N__13134\
        );

    \I__2284\ : Span4Mux_h
    port map (
            O => \N__13142\,
            I => \N__13131\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__13139\,
            I => \N__13128\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__13134\,
            I => \c0.data_in_field_13\
        );

    \I__2281\ : Odrv4
    port map (
            O => \N__13131\,
            I => \c0.data_in_field_13\
        );

    \I__2280\ : Odrv12
    port map (
            O => \N__13128\,
            I => \c0.data_in_field_13\
        );

    \I__2279\ : InMux
    port map (
            O => \N__13121\,
            I => \N__13117\
        );

    \I__2278\ : InMux
    port map (
            O => \N__13120\,
            I => \N__13114\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__13117\,
            I => \c0.n4414\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__13114\,
            I => \c0.n4414\
        );

    \I__2275\ : CascadeMux
    port map (
            O => \N__13109\,
            I => \c0.n30_adj_892_cascade_\
        );

    \I__2274\ : InMux
    port map (
            O => \N__13106\,
            I => \N__13103\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__13103\,
            I => \c0.n25_adj_893\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__13100\,
            I => \N__13095\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__13099\,
            I => \N__13092\
        );

    \I__2270\ : InMux
    port map (
            O => \N__13098\,
            I => \N__13086\
        );

    \I__2269\ : InMux
    port map (
            O => \N__13095\,
            I => \N__13086\
        );

    \I__2268\ : InMux
    port map (
            O => \N__13092\,
            I => \N__13081\
        );

    \I__2267\ : InMux
    port map (
            O => \N__13091\,
            I => \N__13081\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__13086\,
            I => \c0.n2637\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__13081\,
            I => \c0.n2637\
        );

    \I__2264\ : InMux
    port map (
            O => \N__13076\,
            I => \N__13072\
        );

    \I__2263\ : InMux
    port map (
            O => \N__13075\,
            I => \N__13069\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__13072\,
            I => \N__13065\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__13069\,
            I => \N__13062\
        );

    \I__2260\ : InMux
    port map (
            O => \N__13068\,
            I => \N__13059\
        );

    \I__2259\ : Span4Mux_h
    port map (
            O => \N__13065\,
            I => \N__13056\
        );

    \I__2258\ : Span4Mux_h
    port map (
            O => \N__13062\,
            I => \N__13053\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__13059\,
            I => \c0.n1261\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__13056\,
            I => \c0.n1261\
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__13053\,
            I => \c0.n1261\
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__13046\,
            I => \N__13041\
        );

    \I__2253\ : InMux
    port map (
            O => \N__13045\,
            I => \N__13038\
        );

    \I__2252\ : InMux
    port map (
            O => \N__13044\,
            I => \N__13035\
        );

    \I__2251\ : InMux
    port map (
            O => \N__13041\,
            I => \N__13032\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__13038\,
            I => \N__13028\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__13035\,
            I => \N__13023\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__13032\,
            I => \N__13023\
        );

    \I__2247\ : InMux
    port map (
            O => \N__13031\,
            I => \N__13019\
        );

    \I__2246\ : Span4Mux_h
    port map (
            O => \N__13028\,
            I => \N__13014\
        );

    \I__2245\ : Span4Mux_h
    port map (
            O => \N__13023\,
            I => \N__13014\
        );

    \I__2244\ : InMux
    port map (
            O => \N__13022\,
            I => \N__13011\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__13019\,
            I => \c0.data_in_field_45\
        );

    \I__2242\ : Odrv4
    port map (
            O => \N__13014\,
            I => \c0.data_in_field_45\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__13011\,
            I => \c0.data_in_field_45\
        );

    \I__2240\ : InMux
    port map (
            O => \N__13004\,
            I => \N__13001\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__13001\,
            I => \N__12998\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__12998\,
            I => \c0.n14\
        );

    \I__2237\ : InMux
    port map (
            O => \N__12995\,
            I => \N__12992\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__12992\,
            I => \N__12989\
        );

    \I__2235\ : Span4Mux_h
    port map (
            O => \N__12989\,
            I => \N__12986\
        );

    \I__2234\ : Odrv4
    port map (
            O => \N__12986\,
            I => \c0.n12_adj_873\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__12983\,
            I => \c0.n16_cascade_\
        );

    \I__2232\ : InMux
    port map (
            O => \N__12980\,
            I => \N__12977\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__12977\,
            I => \N__12974\
        );

    \I__2230\ : Span4Mux_h
    port map (
            O => \N__12974\,
            I => \N__12971\
        );

    \I__2229\ : Span4Mux_v
    port map (
            O => \N__12971\,
            I => \N__12968\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__12968\,
            I => \c0.n15\
        );

    \I__2227\ : InMux
    port map (
            O => \N__12965\,
            I => \N__12962\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__12962\,
            I => \c0.n24\
        );

    \I__2225\ : InMux
    port map (
            O => \N__12959\,
            I => \N__12956\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__12956\,
            I => \c0.n4388\
        );

    \I__2223\ : CascadeMux
    port map (
            O => \N__12953\,
            I => \N__12950\
        );

    \I__2222\ : InMux
    port map (
            O => \N__12950\,
            I => \N__12947\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__12947\,
            I => \N__12944\
        );

    \I__2220\ : Span4Mux_h
    port map (
            O => \N__12944\,
            I => \N__12941\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__12941\,
            I => \c0.n4445\
        );

    \I__2218\ : InMux
    port map (
            O => \N__12938\,
            I => \N__12935\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__12935\,
            I => \c0.n26_adj_890\
        );

    \I__2216\ : InMux
    port map (
            O => \N__12932\,
            I => \N__12929\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__12929\,
            I => \N__12925\
        );

    \I__2214\ : InMux
    port map (
            O => \N__12928\,
            I => \N__12922\
        );

    \I__2213\ : Span4Mux_h
    port map (
            O => \N__12925\,
            I => \N__12919\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__12922\,
            I => \c0.data_in_frame_6_2\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__12919\,
            I => \c0.data_in_frame_6_2\
        );

    \I__2210\ : InMux
    port map (
            O => \N__12914\,
            I => \N__12911\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__12911\,
            I => \N__12908\
        );

    \I__2208\ : Span4Mux_h
    port map (
            O => \N__12908\,
            I => \N__12905\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__12905\,
            I => \N__12902\
        );

    \I__2206\ : Odrv4
    port map (
            O => \N__12902\,
            I => \c0.n1280\
        );

    \I__2205\ : InMux
    port map (
            O => \N__12899\,
            I => \N__12896\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__12896\,
            I => \N__12892\
        );

    \I__2203\ : InMux
    port map (
            O => \N__12895\,
            I => \N__12889\
        );

    \I__2202\ : Span4Mux_v
    port map (
            O => \N__12892\,
            I => \N__12886\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__12889\,
            I => \N__12883\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__12886\,
            I => \c0.n4390\
        );

    \I__2199\ : Odrv4
    port map (
            O => \N__12883\,
            I => \c0.n4390\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__12878\,
            I => \N__12873\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__12877\,
            I => \N__12870\
        );

    \I__2196\ : InMux
    port map (
            O => \N__12876\,
            I => \N__12867\
        );

    \I__2195\ : InMux
    port map (
            O => \N__12873\,
            I => \N__12863\
        );

    \I__2194\ : InMux
    port map (
            O => \N__12870\,
            I => \N__12860\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__12867\,
            I => \N__12857\
        );

    \I__2192\ : InMux
    port map (
            O => \N__12866\,
            I => \N__12854\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__12863\,
            I => \N__12851\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__12860\,
            I => \c0.data_in_field_47\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__12857\,
            I => \c0.data_in_field_47\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__12854\,
            I => \c0.data_in_field_47\
        );

    \I__2187\ : Odrv4
    port map (
            O => \N__12851\,
            I => \c0.data_in_field_47\
        );

    \I__2186\ : InMux
    port map (
            O => \N__12842\,
            I => \N__12839\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__12839\,
            I => \c0.n4391\
        );

    \I__2184\ : InMux
    port map (
            O => \N__12836\,
            I => \N__12831\
        );

    \I__2183\ : InMux
    port map (
            O => \N__12835\,
            I => \N__12828\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__12834\,
            I => \N__12825\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__12831\,
            I => \N__12822\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__12828\,
            I => \N__12819\
        );

    \I__2179\ : InMux
    port map (
            O => \N__12825\,
            I => \N__12814\
        );

    \I__2178\ : Span4Mux_v
    port map (
            O => \N__12822\,
            I => \N__12809\
        );

    \I__2177\ : Span4Mux_h
    port map (
            O => \N__12819\,
            I => \N__12809\
        );

    \I__2176\ : InMux
    port map (
            O => \N__12818\,
            I => \N__12806\
        );

    \I__2175\ : InMux
    port map (
            O => \N__12817\,
            I => \N__12803\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__12814\,
            I => \c0.data_in_field_1\
        );

    \I__2173\ : Odrv4
    port map (
            O => \N__12809\,
            I => \c0.data_in_field_1\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__12806\,
            I => \c0.data_in_field_1\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__12803\,
            I => \c0.data_in_field_1\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__12794\,
            I => \N__12791\
        );

    \I__2169\ : InMux
    port map (
            O => \N__12791\,
            I => \N__12787\
        );

    \I__2168\ : InMux
    port map (
            O => \N__12790\,
            I => \N__12783\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__12787\,
            I => \N__12780\
        );

    \I__2166\ : InMux
    port map (
            O => \N__12786\,
            I => \N__12776\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__12783\,
            I => \N__12773\
        );

    \I__2164\ : Span12Mux_v
    port map (
            O => \N__12780\,
            I => \N__12770\
        );

    \I__2163\ : InMux
    port map (
            O => \N__12779\,
            I => \N__12767\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__12776\,
            I => \c0.data_in_field_14\
        );

    \I__2161\ : Odrv12
    port map (
            O => \N__12773\,
            I => \c0.data_in_field_14\
        );

    \I__2160\ : Odrv12
    port map (
            O => \N__12770\,
            I => \c0.data_in_field_14\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__12767\,
            I => \c0.data_in_field_14\
        );

    \I__2158\ : InMux
    port map (
            O => \N__12758\,
            I => \N__12755\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__12755\,
            I => \c0.n4474\
        );

    \I__2156\ : InMux
    port map (
            O => \N__12752\,
            I => \N__12749\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__12749\,
            I => \c0.n12_adj_887\
        );

    \I__2154\ : InMux
    port map (
            O => \N__12746\,
            I => \c0.n3922\
        );

    \I__2153\ : SRMux
    port map (
            O => \N__12743\,
            I => \N__12740\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__12740\,
            I => \N__12737\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__12737\,
            I => \c0.n1675\
        );

    \I__2150\ : CEMux
    port map (
            O => \N__12734\,
            I => \N__12731\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__12731\,
            I => \N__12728\
        );

    \I__2148\ : Odrv12
    port map (
            O => \N__12728\,
            I => \c0.n688\
        );

    \I__2147\ : InMux
    port map (
            O => \N__12725\,
            I => \N__12720\
        );

    \I__2146\ : InMux
    port map (
            O => \N__12724\,
            I => \N__12715\
        );

    \I__2145\ : InMux
    port map (
            O => \N__12723\,
            I => \N__12715\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__12720\,
            I => tx2_active
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__12715\,
            I => tx2_active
        );

    \I__2142\ : InMux
    port map (
            O => \N__12710\,
            I => \N__12707\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__12707\,
            I => \c0.n2643\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__12704\,
            I => \c0.n2643_cascade_\
        );

    \I__2139\ : CascadeMux
    port map (
            O => \N__12701\,
            I => \N__12698\
        );

    \I__2138\ : InMux
    port map (
            O => \N__12698\,
            I => \N__12695\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__12695\,
            I => \N__12689\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__12694\,
            I => \N__12685\
        );

    \I__2135\ : InMux
    port map (
            O => \N__12693\,
            I => \N__12680\
        );

    \I__2134\ : InMux
    port map (
            O => \N__12692\,
            I => \N__12680\
        );

    \I__2133\ : Span4Mux_h
    port map (
            O => \N__12689\,
            I => \N__12677\
        );

    \I__2132\ : InMux
    port map (
            O => \N__12688\,
            I => \N__12672\
        );

    \I__2131\ : InMux
    port map (
            O => \N__12685\,
            I => \N__12672\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__12680\,
            I => \c0.tx2_transmit\
        );

    \I__2129\ : Odrv4
    port map (
            O => \N__12677\,
            I => \c0.tx2_transmit\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__12672\,
            I => \c0.tx2_transmit\
        );

    \I__2127\ : InMux
    port map (
            O => \N__12665\,
            I => \N__12662\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__12662\,
            I => \c0.n21\
        );

    \I__2125\ : CascadeMux
    port map (
            O => \N__12659\,
            I => \N__12656\
        );

    \I__2124\ : InMux
    port map (
            O => \N__12656\,
            I => \N__12653\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__12653\,
            I => \c0.n22_adj_881\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__12650\,
            I => \N__12645\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__12649\,
            I => \N__12641\
        );

    \I__2120\ : InMux
    port map (
            O => \N__12648\,
            I => \N__12631\
        );

    \I__2119\ : InMux
    port map (
            O => \N__12645\,
            I => \N__12631\
        );

    \I__2118\ : InMux
    port map (
            O => \N__12644\,
            I => \N__12631\
        );

    \I__2117\ : InMux
    port map (
            O => \N__12641\,
            I => \N__12628\
        );

    \I__2116\ : InMux
    port map (
            O => \N__12640\,
            I => \N__12625\
        );

    \I__2115\ : InMux
    port map (
            O => \N__12639\,
            I => \N__12620\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__12638\,
            I => \N__12616\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__12631\,
            I => \N__12609\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__12628\,
            I => \N__12609\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__12625\,
            I => \N__12609\
        );

    \I__2110\ : InMux
    port map (
            O => \N__12624\,
            I => \N__12604\
        );

    \I__2109\ : InMux
    port map (
            O => \N__12623\,
            I => \N__12604\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__12620\,
            I => \N__12601\
        );

    \I__2107\ : InMux
    port map (
            O => \N__12619\,
            I => \N__12595\
        );

    \I__2106\ : InMux
    port map (
            O => \N__12616\,
            I => \N__12595\
        );

    \I__2105\ : Sp12to4
    port map (
            O => \N__12609\,
            I => \N__12592\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__12604\,
            I => \N__12587\
        );

    \I__2103\ : Span12Mux_s2_v
    port map (
            O => \N__12601\,
            I => \N__12587\
        );

    \I__2102\ : InMux
    port map (
            O => \N__12600\,
            I => \N__12584\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__12595\,
            I => \N__12579\
        );

    \I__2100\ : Span12Mux_v
    port map (
            O => \N__12592\,
            I => \N__12579\
        );

    \I__2099\ : Odrv12
    port map (
            O => \N__12587\,
            I => \r_SM_Main_0_adj_954\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__12584\,
            I => \r_SM_Main_0_adj_954\
        );

    \I__2097\ : Odrv12
    port map (
            O => \N__12579\,
            I => \r_SM_Main_0_adj_954\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__12572\,
            I => \N__12566\
        );

    \I__2095\ : InMux
    port map (
            O => \N__12571\,
            I => \N__12562\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__12570\,
            I => \N__12555\
        );

    \I__2093\ : InMux
    port map (
            O => \N__12569\,
            I => \N__12550\
        );

    \I__2092\ : InMux
    port map (
            O => \N__12566\,
            I => \N__12547\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__12565\,
            I => \N__12544\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__12562\,
            I => \N__12541\
        );

    \I__2089\ : InMux
    port map (
            O => \N__12561\,
            I => \N__12534\
        );

    \I__2088\ : InMux
    port map (
            O => \N__12560\,
            I => \N__12534\
        );

    \I__2087\ : InMux
    port map (
            O => \N__12559\,
            I => \N__12534\
        );

    \I__2086\ : InMux
    port map (
            O => \N__12558\,
            I => \N__12529\
        );

    \I__2085\ : InMux
    port map (
            O => \N__12555\,
            I => \N__12529\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__12554\,
            I => \N__12525\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__12553\,
            I => \N__12521\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__12550\,
            I => \N__12518\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__12547\,
            I => \N__12515\
        );

    \I__2080\ : InMux
    port map (
            O => \N__12544\,
            I => \N__12512\
        );

    \I__2079\ : Span12Mux_s5_v
    port map (
            O => \N__12541\,
            I => \N__12509\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__12534\,
            I => \N__12504\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__12529\,
            I => \N__12504\
        );

    \I__2076\ : InMux
    port map (
            O => \N__12528\,
            I => \N__12501\
        );

    \I__2075\ : InMux
    port map (
            O => \N__12525\,
            I => \N__12494\
        );

    \I__2074\ : InMux
    port map (
            O => \N__12524\,
            I => \N__12494\
        );

    \I__2073\ : InMux
    port map (
            O => \N__12521\,
            I => \N__12494\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__12518\,
            I => \N__12489\
        );

    \I__2071\ : Span4Mux_v
    port map (
            O => \N__12515\,
            I => \N__12489\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__12512\,
            I => \r_SM_Main_1_adj_953\
        );

    \I__2069\ : Odrv12
    port map (
            O => \N__12509\,
            I => \r_SM_Main_1_adj_953\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__12504\,
            I => \r_SM_Main_1_adj_953\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__12501\,
            I => \r_SM_Main_1_adj_953\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__12494\,
            I => \r_SM_Main_1_adj_953\
        );

    \I__2065\ : Odrv4
    port map (
            O => \N__12489\,
            I => \r_SM_Main_1_adj_953\
        );

    \I__2064\ : InMux
    port map (
            O => \N__12476\,
            I => \N__12473\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__12473\,
            I => \N__12470\
        );

    \I__2062\ : Span4Mux_v
    port map (
            O => \N__12470\,
            I => \N__12467\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__12467\,
            I => n4780
        );

    \I__2060\ : InMux
    port map (
            O => \N__12464\,
            I => \N__12450\
        );

    \I__2059\ : InMux
    port map (
            O => \N__12463\,
            I => \N__12450\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__12462\,
            I => \N__12445\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__12461\,
            I => \N__12442\
        );

    \I__2056\ : CascadeMux
    port map (
            O => \N__12460\,
            I => \N__12439\
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__12459\,
            I => \N__12436\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__12458\,
            I => \N__12433\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__12457\,
            I => \N__12430\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__12456\,
            I => \N__12427\
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__12455\,
            I => \N__12424\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__12450\,
            I => \N__12421\
        );

    \I__2049\ : InMux
    port map (
            O => \N__12449\,
            I => \N__12418\
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__12448\,
            I => \N__12415\
        );

    \I__2047\ : InMux
    port map (
            O => \N__12445\,
            I => \N__12398\
        );

    \I__2046\ : InMux
    port map (
            O => \N__12442\,
            I => \N__12398\
        );

    \I__2045\ : InMux
    port map (
            O => \N__12439\,
            I => \N__12398\
        );

    \I__2044\ : InMux
    port map (
            O => \N__12436\,
            I => \N__12398\
        );

    \I__2043\ : InMux
    port map (
            O => \N__12433\,
            I => \N__12389\
        );

    \I__2042\ : InMux
    port map (
            O => \N__12430\,
            I => \N__12389\
        );

    \I__2041\ : InMux
    port map (
            O => \N__12427\,
            I => \N__12389\
        );

    \I__2040\ : InMux
    port map (
            O => \N__12424\,
            I => \N__12389\
        );

    \I__2039\ : Sp12to4
    port map (
            O => \N__12421\,
            I => \N__12384\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__12418\,
            I => \N__12384\
        );

    \I__2037\ : InMux
    port map (
            O => \N__12415\,
            I => \N__12381\
        );

    \I__2036\ : InMux
    port map (
            O => \N__12414\,
            I => \N__12378\
        );

    \I__2035\ : InMux
    port map (
            O => \N__12413\,
            I => \N__12371\
        );

    \I__2034\ : InMux
    port map (
            O => \N__12412\,
            I => \N__12371\
        );

    \I__2033\ : InMux
    port map (
            O => \N__12411\,
            I => \N__12371\
        );

    \I__2032\ : InMux
    port map (
            O => \N__12410\,
            I => \N__12368\
        );

    \I__2031\ : InMux
    port map (
            O => \N__12409\,
            I => \N__12361\
        );

    \I__2030\ : InMux
    port map (
            O => \N__12408\,
            I => \N__12361\
        );

    \I__2029\ : InMux
    port map (
            O => \N__12407\,
            I => \N__12361\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__12398\,
            I => \N__12356\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__12389\,
            I => \N__12356\
        );

    \I__2026\ : Odrv12
    port map (
            O => \N__12384\,
            I => \r_SM_Main_2_adj_952\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__12381\,
            I => \r_SM_Main_2_adj_952\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__12378\,
            I => \r_SM_Main_2_adj_952\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__12371\,
            I => \r_SM_Main_2_adj_952\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__12368\,
            I => \r_SM_Main_2_adj_952\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__12361\,
            I => \r_SM_Main_2_adj_952\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__12356\,
            I => \r_SM_Main_2_adj_952\
        );

    \I__2019\ : CascadeMux
    port map (
            O => \N__12341\,
            I => \n3_cascade_\
        );

    \I__2018\ : InMux
    port map (
            O => \N__12338\,
            I => \N__12335\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__12335\,
            I => \N__12331\
        );

    \I__2016\ : InMux
    port map (
            O => \N__12334\,
            I => \N__12328\
        );

    \I__2015\ : Odrv12
    port map (
            O => \N__12331\,
            I => rx_data_6
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__12328\,
            I => rx_data_6
        );

    \I__2013\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12320\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__12320\,
            I => \c0.rx.n4876\
        );

    \I__2011\ : IoInMux
    port map (
            O => \N__12317\,
            I => \N__12314\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__12314\,
            I => tx_enable
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__12311\,
            I => \N__12305\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__12310\,
            I => \N__12302\
        );

    \I__2007\ : InMux
    port map (
            O => \N__12309\,
            I => \N__12299\
        );

    \I__2006\ : InMux
    port map (
            O => \N__12308\,
            I => \N__12296\
        );

    \I__2005\ : InMux
    port map (
            O => \N__12305\,
            I => \N__12291\
        );

    \I__2004\ : InMux
    port map (
            O => \N__12302\,
            I => \N__12291\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__12299\,
            I => data_in_7_5
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__12296\,
            I => data_in_7_5
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__12291\,
            I => data_in_7_5
        );

    \I__2000\ : InMux
    port map (
            O => \N__12284\,
            I => \N__12280\
        );

    \I__1999\ : InMux
    port map (
            O => \N__12283\,
            I => \N__12277\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__12280\,
            I => \N__12274\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__12277\,
            I => \N__12269\
        );

    \I__1996\ : Span4Mux_s3_h
    port map (
            O => \N__12274\,
            I => \N__12266\
        );

    \I__1995\ : InMux
    port map (
            O => \N__12273\,
            I => \N__12263\
        );

    \I__1994\ : InMux
    port map (
            O => \N__12272\,
            I => \N__12260\
        );

    \I__1993\ : Span4Mux_v
    port map (
            O => \N__12269\,
            I => \N__12257\
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__12266\,
            I => data_in_6_5
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__12263\,
            I => data_in_6_5
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__12260\,
            I => data_in_6_5
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__12257\,
            I => data_in_6_5
        );

    \I__1988\ : InMux
    port map (
            O => \N__12248\,
            I => \N__12245\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__12245\,
            I => n4519
        );

    \I__1986\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12239\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__12239\,
            I => n4520
        );

    \I__1984\ : InMux
    port map (
            O => \N__12236\,
            I => \N__12233\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__12233\,
            I => \N__12230\
        );

    \I__1982\ : Span4Mux_v
    port map (
            O => \N__12230\,
            I => \N__12226\
        );

    \I__1981\ : InMux
    port map (
            O => \N__12229\,
            I => \N__12223\
        );

    \I__1980\ : Odrv4
    port map (
            O => \N__12226\,
            I => blink_counter_25
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__12223\,
            I => blink_counter_25
        );

    \I__1978\ : IoInMux
    port map (
            O => \N__12218\,
            I => \N__12215\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__12215\,
            I => \N__12212\
        );

    \I__1976\ : Span12Mux_s9_v
    port map (
            O => \N__12212\,
            I => \N__12209\
        );

    \I__1975\ : Odrv12
    port map (
            O => \N__12209\,
            I => \LED_c\
        );

    \I__1974\ : InMux
    port map (
            O => \N__12206\,
            I => \c0.n3921\
        );

    \I__1973\ : InMux
    port map (
            O => \N__12203\,
            I => \N__12199\
        );

    \I__1972\ : InMux
    port map (
            O => \N__12202\,
            I => \N__12196\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__12199\,
            I => \c0.data_in_frame_6_1\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__12196\,
            I => \c0.data_in_frame_6_1\
        );

    \I__1969\ : InMux
    port map (
            O => \N__12191\,
            I => \N__12187\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__12190\,
            I => \N__12184\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__12187\,
            I => \N__12181\
        );

    \I__1966\ : InMux
    port map (
            O => \N__12184\,
            I => \N__12177\
        );

    \I__1965\ : Span4Mux_v
    port map (
            O => \N__12181\,
            I => \N__12174\
        );

    \I__1964\ : InMux
    port map (
            O => \N__12180\,
            I => \N__12171\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__12177\,
            I => data_in_5_4
        );

    \I__1962\ : Odrv4
    port map (
            O => \N__12174\,
            I => data_in_5_4
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__12171\,
            I => data_in_5_4
        );

    \I__1960\ : InMux
    port map (
            O => \N__12164\,
            I => \N__12160\
        );

    \I__1959\ : InMux
    port map (
            O => \N__12163\,
            I => \N__12156\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__12160\,
            I => \N__12153\
        );

    \I__1957\ : InMux
    port map (
            O => \N__12159\,
            I => \N__12150\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__12156\,
            I => \c0.data_in_field_44\
        );

    \I__1955\ : Odrv12
    port map (
            O => \N__12153\,
            I => \c0.data_in_field_44\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__12150\,
            I => \c0.data_in_field_44\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__12143\,
            I => \N__12140\
        );

    \I__1952\ : InMux
    port map (
            O => \N__12140\,
            I => \N__12134\
        );

    \I__1951\ : InMux
    port map (
            O => \N__12139\,
            I => \N__12131\
        );

    \I__1950\ : InMux
    port map (
            O => \N__12138\,
            I => \N__12128\
        );

    \I__1949\ : InMux
    port map (
            O => \N__12137\,
            I => \N__12125\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__12134\,
            I => \N__12122\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__12131\,
            I => data_in_3_4
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__12128\,
            I => data_in_3_4
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__12125\,
            I => data_in_3_4
        );

    \I__1944\ : Odrv12
    port map (
            O => \N__12122\,
            I => data_in_3_4
        );

    \I__1943\ : InMux
    port map (
            O => \N__12113\,
            I => \N__12109\
        );

    \I__1942\ : InMux
    port map (
            O => \N__12112\,
            I => \N__12106\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__12109\,
            I => \N__12101\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__12106\,
            I => \N__12098\
        );

    \I__1939\ : InMux
    port map (
            O => \N__12105\,
            I => \N__12095\
        );

    \I__1938\ : InMux
    port map (
            O => \N__12104\,
            I => \N__12092\
        );

    \I__1937\ : Span4Mux_s3_h
    port map (
            O => \N__12101\,
            I => \N__12089\
        );

    \I__1936\ : Span4Mux_s1_h
    port map (
            O => \N__12098\,
            I => \N__12084\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__12095\,
            I => \N__12084\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__12092\,
            I => data_in_2_4
        );

    \I__1933\ : Odrv4
    port map (
            O => \N__12089\,
            I => data_in_2_4
        );

    \I__1932\ : Odrv4
    port map (
            O => \N__12084\,
            I => data_in_2_4
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__12077\,
            I => \N__12074\
        );

    \I__1930\ : InMux
    port map (
            O => \N__12074\,
            I => \N__12068\
        );

    \I__1929\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12068\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__12068\,
            I => rx_data_5
        );

    \I__1927\ : InMux
    port map (
            O => \N__12065\,
            I => \N__12061\
        );

    \I__1926\ : CascadeMux
    port map (
            O => \N__12064\,
            I => \N__12058\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__12061\,
            I => \N__12055\
        );

    \I__1924\ : InMux
    port map (
            O => \N__12058\,
            I => \N__12052\
        );

    \I__1923\ : Odrv12
    port map (
            O => \N__12055\,
            I => rx_data_7
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__12052\,
            I => rx_data_7
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__12047\,
            I => \N__12043\
        );

    \I__1920\ : InMux
    port map (
            O => \N__12046\,
            I => \N__12039\
        );

    \I__1919\ : InMux
    port map (
            O => \N__12043\,
            I => \N__12034\
        );

    \I__1918\ : InMux
    port map (
            O => \N__12042\,
            I => \N__12031\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__12039\,
            I => \N__12028\
        );

    \I__1916\ : InMux
    port map (
            O => \N__12038\,
            I => \N__12023\
        );

    \I__1915\ : InMux
    port map (
            O => \N__12037\,
            I => \N__12023\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__12034\,
            I => \N__12020\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__12031\,
            I => \N__12017\
        );

    \I__1912\ : Odrv4
    port map (
            O => \N__12028\,
            I => \c0.data_in_field_39\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__12023\,
            I => \c0.data_in_field_39\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__12020\,
            I => \c0.data_in_field_39\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__12017\,
            I => \c0.data_in_field_39\
        );

    \I__1908\ : InMux
    port map (
            O => \N__12008\,
            I => \N__12004\
        );

    \I__1907\ : InMux
    port map (
            O => \N__12007\,
            I => \N__11999\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__12004\,
            I => \N__11996\
        );

    \I__1905\ : InMux
    port map (
            O => \N__12003\,
            I => \N__11991\
        );

    \I__1904\ : InMux
    port map (
            O => \N__12002\,
            I => \N__11991\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__11999\,
            I => \c0.data_in_field_38\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__11996\,
            I => \c0.data_in_field_38\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__11991\,
            I => \c0.data_in_field_38\
        );

    \I__1900\ : InMux
    port map (
            O => \N__11984\,
            I => \N__11980\
        );

    \I__1899\ : InMux
    port map (
            O => \N__11983\,
            I => \N__11975\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__11980\,
            I => \N__11972\
        );

    \I__1897\ : InMux
    port map (
            O => \N__11979\,
            I => \N__11969\
        );

    \I__1896\ : InMux
    port map (
            O => \N__11978\,
            I => \N__11966\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__11975\,
            I => \N__11963\
        );

    \I__1894\ : Span4Mux_s3_h
    port map (
            O => \N__11972\,
            I => \N__11960\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__11969\,
            I => \N__11957\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__11966\,
            I => data_in_6_4
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__11963\,
            I => data_in_6_4
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__11960\,
            I => data_in_6_4
        );

    \I__1889\ : Odrv12
    port map (
            O => \N__11957\,
            I => data_in_6_4
        );

    \I__1888\ : InMux
    port map (
            O => \N__11948\,
            I => \N__11945\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__11945\,
            I => \N__11940\
        );

    \I__1886\ : InMux
    port map (
            O => \N__11944\,
            I => \N__11935\
        );

    \I__1885\ : InMux
    port map (
            O => \N__11943\,
            I => \N__11935\
        );

    \I__1884\ : Span4Mux_s3_h
    port map (
            O => \N__11940\,
            I => \N__11932\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__11935\,
            I => data_in_4_4
        );

    \I__1882\ : Odrv4
    port map (
            O => \N__11932\,
            I => data_in_4_4
        );

    \I__1881\ : InMux
    port map (
            O => \N__11927\,
            I => \N__11924\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__11924\,
            I => \c0.n8_adj_872\
        );

    \I__1879\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11918\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__11918\,
            I => \N__11914\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__11917\,
            I => \N__11910\
        );

    \I__1876\ : Span4Mux_h
    port map (
            O => \N__11914\,
            I => \N__11907\
        );

    \I__1875\ : InMux
    port map (
            O => \N__11913\,
            I => \N__11902\
        );

    \I__1874\ : InMux
    port map (
            O => \N__11910\,
            I => \N__11902\
        );

    \I__1873\ : Odrv4
    port map (
            O => \N__11907\,
            I => data_in_0_2
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__11902\,
            I => data_in_0_2
        );

    \I__1871\ : InMux
    port map (
            O => \N__11897\,
            I => \N__11893\
        );

    \I__1870\ : InMux
    port map (
            O => \N__11896\,
            I => \N__11888\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__11893\,
            I => \N__11885\
        );

    \I__1868\ : InMux
    port map (
            O => \N__11892\,
            I => \N__11882\
        );

    \I__1867\ : InMux
    port map (
            O => \N__11891\,
            I => \N__11879\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__11888\,
            I => \c0.data_in_field_2\
        );

    \I__1865\ : Odrv12
    port map (
            O => \N__11885\,
            I => \c0.data_in_field_2\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__11882\,
            I => \c0.data_in_field_2\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__11879\,
            I => \c0.data_in_field_2\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__11870\,
            I => \N__11867\
        );

    \I__1861\ : InMux
    port map (
            O => \N__11867\,
            I => \N__11861\
        );

    \I__1860\ : InMux
    port map (
            O => \N__11866\,
            I => \N__11861\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__11861\,
            I => \c0.data_in_frame_7_1\
        );

    \I__1858\ : InMux
    port map (
            O => \N__11858\,
            I => \N__11855\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__11855\,
            I => \N__11852\
        );

    \I__1856\ : Span4Mux_s3_h
    port map (
            O => \N__11852\,
            I => \N__11849\
        );

    \I__1855\ : Span4Mux_v
    port map (
            O => \N__11849\,
            I => \N__11846\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__11846\,
            I => \c0.n4607\
        );

    \I__1853\ : InMux
    port map (
            O => \N__11843\,
            I => \N__11840\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__11840\,
            I => \N__11835\
        );

    \I__1851\ : InMux
    port map (
            O => \N__11839\,
            I => \N__11829\
        );

    \I__1850\ : InMux
    port map (
            O => \N__11838\,
            I => \N__11829\
        );

    \I__1849\ : Span4Mux_v
    port map (
            O => \N__11835\,
            I => \N__11826\
        );

    \I__1848\ : InMux
    port map (
            O => \N__11834\,
            I => \N__11823\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__11829\,
            I => \N__11820\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__11826\,
            I => data_in_3_6
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__11823\,
            I => data_in_3_6
        );

    \I__1844\ : Odrv12
    port map (
            O => \N__11820\,
            I => data_in_3_6
        );

    \I__1843\ : CascadeMux
    port map (
            O => \N__11813\,
            I => \N__11810\
        );

    \I__1842\ : InMux
    port map (
            O => \N__11810\,
            I => \N__11807\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__11807\,
            I => \N__11802\
        );

    \I__1840\ : InMux
    port map (
            O => \N__11806\,
            I => \N__11798\
        );

    \I__1839\ : InMux
    port map (
            O => \N__11805\,
            I => \N__11795\
        );

    \I__1838\ : Span4Mux_h
    port map (
            O => \N__11802\,
            I => \N__11792\
        );

    \I__1837\ : InMux
    port map (
            O => \N__11801\,
            I => \N__11789\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__11798\,
            I => data_in_1_1
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__11795\,
            I => data_in_1_1
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__11792\,
            I => data_in_1_1
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__11789\,
            I => data_in_1_1
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__11780\,
            I => \c0.n8_adj_871_cascade_\
        );

    \I__1831\ : InMux
    port map (
            O => \N__11777\,
            I => \N__11774\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__11774\,
            I => \c0.n12\
        );

    \I__1829\ : InMux
    port map (
            O => \N__11771\,
            I => \N__11768\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__11768\,
            I => \c0.n1418\
        );

    \I__1827\ : InMux
    port map (
            O => \N__11765\,
            I => \N__11762\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__11762\,
            I => \N__11758\
        );

    \I__1825\ : InMux
    port map (
            O => \N__11761\,
            I => \N__11752\
        );

    \I__1824\ : Span4Mux_v
    port map (
            O => \N__11758\,
            I => \N__11749\
        );

    \I__1823\ : InMux
    port map (
            O => \N__11757\,
            I => \N__11746\
        );

    \I__1822\ : InMux
    port map (
            O => \N__11756\,
            I => \N__11743\
        );

    \I__1821\ : InMux
    port map (
            O => \N__11755\,
            I => \N__11740\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__11752\,
            I => \c0.data_in_field_4\
        );

    \I__1819\ : Odrv4
    port map (
            O => \N__11749\,
            I => \c0.data_in_field_4\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__11746\,
            I => \c0.data_in_field_4\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__11743\,
            I => \c0.data_in_field_4\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__11740\,
            I => \c0.data_in_field_4\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__11729\,
            I => \c0.n1418_cascade_\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__11726\,
            I => \c0.n4474_cascade_\
        );

    \I__1813\ : InMux
    port map (
            O => \N__11723\,
            I => \N__11720\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__11720\,
            I => \N__11717\
        );

    \I__1811\ : Span4Mux_h
    port map (
            O => \N__11717\,
            I => \N__11712\
        );

    \I__1810\ : InMux
    port map (
            O => \N__11716\,
            I => \N__11707\
        );

    \I__1809\ : InMux
    port map (
            O => \N__11715\,
            I => \N__11707\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__11712\,
            I => data_in_4_6
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__11707\,
            I => data_in_4_6
        );

    \I__1806\ : InMux
    port map (
            O => \N__11702\,
            I => \N__11699\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__11699\,
            I => \N__11696\
        );

    \I__1804\ : Odrv12
    port map (
            O => \N__11696\,
            I => \c0.n4396\
        );

    \I__1803\ : InMux
    port map (
            O => \N__11693\,
            I => \N__11689\
        );

    \I__1802\ : InMux
    port map (
            O => \N__11692\,
            I => \N__11686\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__11689\,
            I => \N__11681\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__11686\,
            I => \N__11678\
        );

    \I__1799\ : InMux
    port map (
            O => \N__11685\,
            I => \N__11673\
        );

    \I__1798\ : InMux
    port map (
            O => \N__11684\,
            I => \N__11673\
        );

    \I__1797\ : Odrv4
    port map (
            O => \N__11681\,
            I => \c0.data_in_field_21\
        );

    \I__1796\ : Odrv4
    port map (
            O => \N__11678\,
            I => \c0.data_in_field_21\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__11673\,
            I => \c0.data_in_field_21\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__11666\,
            I => \c0.n4396_cascade_\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__11663\,
            I => \N__11658\
        );

    \I__1792\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11655\
        );

    \I__1791\ : InMux
    port map (
            O => \N__11661\,
            I => \N__11649\
        );

    \I__1790\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11649\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__11655\,
            I => \N__11646\
        );

    \I__1788\ : InMux
    port map (
            O => \N__11654\,
            I => \N__11643\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__11649\,
            I => \c0.data_in_field_7\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__11646\,
            I => \c0.data_in_field_7\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__11643\,
            I => \c0.data_in_field_7\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11636\,
            I => \N__11632\
        );

    \I__1783\ : InMux
    port map (
            O => \N__11635\,
            I => \N__11628\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__11632\,
            I => \N__11625\
        );

    \I__1781\ : InMux
    port map (
            O => \N__11631\,
            I => \N__11621\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__11628\,
            I => \N__11618\
        );

    \I__1779\ : Span4Mux_h
    port map (
            O => \N__11625\,
            I => \N__11615\
        );

    \I__1778\ : InMux
    port map (
            O => \N__11624\,
            I => \N__11612\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__11621\,
            I => \c0.data_in_field_0\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__11618\,
            I => \c0.data_in_field_0\
        );

    \I__1775\ : Odrv4
    port map (
            O => \N__11615\,
            I => \c0.data_in_field_0\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__11612\,
            I => \c0.data_in_field_0\
        );

    \I__1773\ : InMux
    port map (
            O => \N__11603\,
            I => \N__11597\
        );

    \I__1772\ : InMux
    port map (
            O => \N__11602\,
            I => \N__11597\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__11597\,
            I => \N__11593\
        );

    \I__1770\ : InMux
    port map (
            O => \N__11596\,
            I => \N__11589\
        );

    \I__1769\ : Span4Mux_v
    port map (
            O => \N__11593\,
            I => \N__11586\
        );

    \I__1768\ : InMux
    port map (
            O => \N__11592\,
            I => \N__11583\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__11589\,
            I => \c0.data_in_field_8\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__11586\,
            I => \c0.data_in_field_8\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__11583\,
            I => \c0.data_in_field_8\
        );

    \I__1764\ : InMux
    port map (
            O => \N__11576\,
            I => \N__11573\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__11573\,
            I => \N__11570\
        );

    \I__1762\ : Span4Mux_v
    port map (
            O => \N__11570\,
            I => \N__11567\
        );

    \I__1761\ : Odrv4
    port map (
            O => \N__11567\,
            I => \c0.n4570\
        );

    \I__1760\ : InMux
    port map (
            O => \N__11564\,
            I => \N__11561\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__11561\,
            I => \c0.n17\
        );

    \I__1758\ : InMux
    port map (
            O => \N__11558\,
            I => \N__11555\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__11555\,
            I => \c0.n4430\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__11552\,
            I => \N__11549\
        );

    \I__1755\ : InMux
    port map (
            O => \N__11549\,
            I => \N__11546\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__11546\,
            I => \c0.n15_adj_885\
        );

    \I__1753\ : InMux
    port map (
            O => \N__11543\,
            I => \N__11540\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__11540\,
            I => \c0.n16_adj_884\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__11537\,
            I => \c0.n17_adj_889_cascade_\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__11534\,
            I => \c0.n4387_cascade_\
        );

    \I__1749\ : InMux
    port map (
            O => \N__11531\,
            I => \N__11527\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__11530\,
            I => \N__11524\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__11527\,
            I => \N__11521\
        );

    \I__1746\ : InMux
    port map (
            O => \N__11524\,
            I => \N__11518\
        );

    \I__1745\ : Span4Mux_s1_v
    port map (
            O => \N__11521\,
            I => \N__11515\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__11518\,
            I => \N__11511\
        );

    \I__1743\ : Span4Mux_v
    port map (
            O => \N__11515\,
            I => \N__11508\
        );

    \I__1742\ : InMux
    port map (
            O => \N__11514\,
            I => \N__11505\
        );

    \I__1741\ : Odrv12
    port map (
            O => \N__11511\,
            I => data_in_4_7
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__11508\,
            I => data_in_4_7
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__11505\,
            I => data_in_4_7
        );

    \I__1738\ : InMux
    port map (
            O => \N__11498\,
            I => \N__11494\
        );

    \I__1737\ : InMux
    port map (
            O => \N__11497\,
            I => \N__11491\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__11494\,
            I => \N__11488\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__11491\,
            I => \N__11482\
        );

    \I__1734\ : Span4Mux_s3_h
    port map (
            O => \N__11488\,
            I => \N__11482\
        );

    \I__1733\ : InMux
    port map (
            O => \N__11487\,
            I => \N__11479\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__11482\,
            I => data_in_5_7
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__11479\,
            I => data_in_5_7
        );

    \I__1730\ : InMux
    port map (
            O => \N__11474\,
            I => \N__11471\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__11471\,
            I => \N__11466\
        );

    \I__1728\ : InMux
    port map (
            O => \N__11470\,
            I => \N__11461\
        );

    \I__1727\ : InMux
    port map (
            O => \N__11469\,
            I => \N__11461\
        );

    \I__1726\ : Span4Mux_s3_h
    port map (
            O => \N__11466\,
            I => \N__11458\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__11461\,
            I => \c0.n1296\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__11458\,
            I => \c0.n1296\
        );

    \I__1723\ : InMux
    port map (
            O => \N__11453\,
            I => \N__11450\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__11450\,
            I => \c0.n11_adj_888\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__11447\,
            I => \N__11444\
        );

    \I__1720\ : InMux
    port map (
            O => \N__11444\,
            I => \N__11441\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__11441\,
            I => \N__11436\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__11440\,
            I => \N__11432\
        );

    \I__1717\ : InMux
    port map (
            O => \N__11439\,
            I => \N__11429\
        );

    \I__1716\ : Span4Mux_h
    port map (
            O => \N__11436\,
            I => \N__11426\
        );

    \I__1715\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11421\
        );

    \I__1714\ : InMux
    port map (
            O => \N__11432\,
            I => \N__11421\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__11429\,
            I => data_in_2_7
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__11426\,
            I => data_in_2_7
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__11421\,
            I => data_in_2_7
        );

    \I__1710\ : InMux
    port map (
            O => \N__11414\,
            I => \N__11404\
        );

    \I__1709\ : InMux
    port map (
            O => \N__11413\,
            I => \N__11404\
        );

    \I__1708\ : InMux
    port map (
            O => \N__11412\,
            I => \N__11404\
        );

    \I__1707\ : InMux
    port map (
            O => \N__11411\,
            I => \N__11400\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__11404\,
            I => \N__11397\
        );

    \I__1705\ : InMux
    port map (
            O => \N__11403\,
            I => \N__11394\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__11400\,
            I => \r_SM_Main_2_N_759_1\
        );

    \I__1703\ : Odrv12
    port map (
            O => \N__11397\,
            I => \r_SM_Main_2_N_759_1\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__11394\,
            I => \r_SM_Main_2_N_759_1\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__11387\,
            I => \n4366_cascade_\
        );

    \I__1700\ : InMux
    port map (
            O => \N__11384\,
            I => \N__11380\
        );

    \I__1699\ : InMux
    port map (
            O => \N__11383\,
            I => \N__11377\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__11380\,
            I => \N__11374\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__11377\,
            I => \N__11370\
        );

    \I__1696\ : Span4Mux_v
    port map (
            O => \N__11374\,
            I => \N__11367\
        );

    \I__1695\ : InMux
    port map (
            O => \N__11373\,
            I => \N__11364\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__11370\,
            I => data_in_4_2
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__11367\,
            I => data_in_4_2
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__11364\,
            I => data_in_4_2
        );

    \I__1691\ : InMux
    port map (
            O => \N__11357\,
            I => \N__11352\
        );

    \I__1690\ : InMux
    port map (
            O => \N__11356\,
            I => \N__11349\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__11355\,
            I => \N__11346\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__11352\,
            I => \N__11343\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__11349\,
            I => \N__11340\
        );

    \I__1686\ : InMux
    port map (
            O => \N__11346\,
            I => \N__11335\
        );

    \I__1685\ : Span4Mux_v
    port map (
            O => \N__11343\,
            I => \N__11332\
        );

    \I__1684\ : Span4Mux_v
    port map (
            O => \N__11340\,
            I => \N__11329\
        );

    \I__1683\ : InMux
    port map (
            O => \N__11339\,
            I => \N__11326\
        );

    \I__1682\ : InMux
    port map (
            O => \N__11338\,
            I => \N__11323\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__11335\,
            I => \c0.data_in_field_11\
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__11332\,
            I => \c0.data_in_field_11\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__11329\,
            I => \c0.data_in_field_11\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__11326\,
            I => \c0.data_in_field_11\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__11323\,
            I => \c0.data_in_field_11\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__11312\,
            I => \c0.n8_adj_879_cascade_\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__11309\,
            I => \c0.n4451_cascade_\
        );

    \I__1674\ : InMux
    port map (
            O => \N__11306\,
            I => \N__11303\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__11303\,
            I => \N__11300\
        );

    \I__1672\ : Odrv4
    port map (
            O => \N__11300\,
            I => \c0.n8_adj_880\
        );

    \I__1671\ : InMux
    port map (
            O => \N__11297\,
            I => \N__11294\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__11294\,
            I => \N__11291\
        );

    \I__1669\ : Odrv12
    port map (
            O => \N__11291\,
            I => \c0.n10_adj_876\
        );

    \I__1668\ : InMux
    port map (
            O => \N__11288\,
            I => \N__11285\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__11285\,
            I => \c0.n4469\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__11282\,
            I => \c0.n1357_cascade_\
        );

    \I__1665\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11276\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__11276\,
            I => \N__11273\
        );

    \I__1663\ : Span4Mux_h
    port map (
            O => \N__11273\,
            I => \N__11269\
        );

    \I__1662\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11266\
        );

    \I__1661\ : Odrv4
    port map (
            O => \N__11269\,
            I => \c0.n4399\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__11266\,
            I => \c0.n4399\
        );

    \I__1659\ : InMux
    port map (
            O => \N__11261\,
            I => \N__11258\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__11258\,
            I => \c0.n4819\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__11255\,
            I => \c0.n4549_cascade_\
        );

    \I__1656\ : InMux
    port map (
            O => \N__11252\,
            I => \N__11249\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__11249\,
            I => \N__11243\
        );

    \I__1654\ : InMux
    port map (
            O => \N__11248\,
            I => \N__11236\
        );

    \I__1653\ : InMux
    port map (
            O => \N__11247\,
            I => \N__11236\
        );

    \I__1652\ : InMux
    port map (
            O => \N__11246\,
            I => \N__11236\
        );

    \I__1651\ : Span4Mux_v
    port map (
            O => \N__11243\,
            I => \N__11231\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__11236\,
            I => \N__11231\
        );

    \I__1649\ : Span4Mux_v
    port map (
            O => \N__11231\,
            I => \N__11224\
        );

    \I__1648\ : InMux
    port map (
            O => \N__11230\,
            I => \N__11219\
        );

    \I__1647\ : InMux
    port map (
            O => \N__11229\,
            I => \N__11219\
        );

    \I__1646\ : InMux
    port map (
            O => \N__11228\,
            I => \N__11216\
        );

    \I__1645\ : InMux
    port map (
            O => \N__11227\,
            I => \N__11213\
        );

    \I__1644\ : Odrv4
    port map (
            O => \N__11224\,
            I => n1030
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__11219\,
            I => n1030
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__11216\,
            I => n1030
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__11213\,
            I => n1030
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__11204\,
            I => \tx2_data_4_keep_cascade_\
        );

    \I__1639\ : InMux
    port map (
            O => \N__11201\,
            I => \N__11197\
        );

    \I__1638\ : InMux
    port map (
            O => \N__11200\,
            I => \N__11194\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__11197\,
            I => \r_Tx_Data_4_adj_960\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__11194\,
            I => \r_Tx_Data_4_adj_960\
        );

    \I__1635\ : InMux
    port map (
            O => \N__11189\,
            I => \N__11186\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__11186\,
            I => \c0.n4597\
        );

    \I__1633\ : InMux
    port map (
            O => \N__11183\,
            I => \N__11179\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__11182\,
            I => \N__11176\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__11179\,
            I => \N__11173\
        );

    \I__1630\ : InMux
    port map (
            O => \N__11176\,
            I => \N__11169\
        );

    \I__1629\ : Span4Mux_h
    port map (
            O => \N__11173\,
            I => \N__11166\
        );

    \I__1628\ : InMux
    port map (
            O => \N__11172\,
            I => \N__11163\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__11169\,
            I => \c0.data_in_field_20\
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__11166\,
            I => \c0.data_in_field_20\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__11163\,
            I => \c0.data_in_field_20\
        );

    \I__1624\ : InMux
    port map (
            O => \N__11156\,
            I => \N__11153\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__11153\,
            I => \c0.n4550\
        );

    \I__1622\ : InMux
    port map (
            O => \N__11150\,
            I => \N__11147\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__11147\,
            I => \c0.tx2.n23\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__11144\,
            I => \n865_cascade_\
        );

    \I__1619\ : InMux
    port map (
            O => \N__11141\,
            I => \N__11138\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__11138\,
            I => \c0.n4543\
        );

    \I__1617\ : InMux
    port map (
            O => \N__11135\,
            I => \N__11129\
        );

    \I__1616\ : InMux
    port map (
            O => \N__11134\,
            I => \N__11129\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__11129\,
            I => \N__11126\
        );

    \I__1614\ : Span4Mux_h
    port map (
            O => \N__11126\,
            I => \N__11122\
        );

    \I__1613\ : InMux
    port map (
            O => \N__11125\,
            I => \N__11119\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__11122\,
            I => blink_counter_22
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__11119\,
            I => blink_counter_22
        );

    \I__1610\ : InMux
    port map (
            O => \N__11114\,
            I => \N__11108\
        );

    \I__1609\ : InMux
    port map (
            O => \N__11113\,
            I => \N__11108\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__11108\,
            I => \N__11105\
        );

    \I__1607\ : Span4Mux_v
    port map (
            O => \N__11105\,
            I => \N__11101\
        );

    \I__1606\ : InMux
    port map (
            O => \N__11104\,
            I => \N__11098\
        );

    \I__1605\ : Odrv4
    port map (
            O => \N__11101\,
            I => blink_counter_24
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__11098\,
            I => blink_counter_24
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__11093\,
            I => \N__11090\
        );

    \I__1602\ : InMux
    port map (
            O => \N__11090\,
            I => \N__11084\
        );

    \I__1601\ : InMux
    port map (
            O => \N__11089\,
            I => \N__11084\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__11084\,
            I => \N__11081\
        );

    \I__1599\ : Span4Mux_h
    port map (
            O => \N__11081\,
            I => \N__11077\
        );

    \I__1598\ : InMux
    port map (
            O => \N__11080\,
            I => \N__11074\
        );

    \I__1597\ : Odrv4
    port map (
            O => \N__11077\,
            I => blink_counter_21
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__11074\,
            I => blink_counter_21
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__11069\,
            I => \N__11065\
        );

    \I__1594\ : InMux
    port map (
            O => \N__11068\,
            I => \N__11060\
        );

    \I__1593\ : InMux
    port map (
            O => \N__11065\,
            I => \N__11060\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__11060\,
            I => \N__11057\
        );

    \I__1591\ : Span4Mux_h
    port map (
            O => \N__11057\,
            I => \N__11053\
        );

    \I__1590\ : InMux
    port map (
            O => \N__11056\,
            I => \N__11050\
        );

    \I__1589\ : Odrv4
    port map (
            O => \N__11053\,
            I => blink_counter_23
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__11050\,
            I => blink_counter_23
        );

    \I__1587\ : InMux
    port map (
            O => \N__11045\,
            I => \N__11042\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__11042\,
            I => \N__11039\
        );

    \I__1585\ : Span4Mux_h
    port map (
            O => \N__11039\,
            I => \N__11036\
        );

    \I__1584\ : Span4Mux_v
    port map (
            O => \N__11036\,
            I => \N__11033\
        );

    \I__1583\ : Odrv4
    port map (
            O => \N__11033\,
            I => \c0.n4580\
        );

    \I__1582\ : InMux
    port map (
            O => \N__11030\,
            I => \N__11027\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__11027\,
            I => \N__11024\
        );

    \I__1580\ : Span4Mux_v
    port map (
            O => \N__11024\,
            I => \N__11021\
        );

    \I__1579\ : Odrv4
    port map (
            O => \N__11021\,
            I => \c0.n4571\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__11018\,
            I => \c0.n4855_cascade_\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__11015\,
            I => \tx2_data_0_keep_cascade_\
        );

    \I__1576\ : InMux
    port map (
            O => \N__11012\,
            I => \N__11008\
        );

    \I__1575\ : InMux
    port map (
            O => \N__11011\,
            I => \N__11005\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__11008\,
            I => \r_Tx_Data_0_adj_964\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__11005\,
            I => \r_Tx_Data_0_adj_964\
        );

    \I__1572\ : InMux
    port map (
            O => \N__11000\,
            I => \N__10996\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__10999\,
            I => \N__10993\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__10996\,
            I => \N__10990\
        );

    \I__1569\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10984\
        );

    \I__1568\ : Span4Mux_v
    port map (
            O => \N__10990\,
            I => \N__10981\
        );

    \I__1567\ : InMux
    port map (
            O => \N__10989\,
            I => \N__10976\
        );

    \I__1566\ : InMux
    port map (
            O => \N__10988\,
            I => \N__10976\
        );

    \I__1565\ : InMux
    port map (
            O => \N__10987\,
            I => \N__10973\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__10984\,
            I => \c0.data_in_field_32\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__10981\,
            I => \c0.data_in_field_32\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__10976\,
            I => \c0.data_in_field_32\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__10973\,
            I => \c0.data_in_field_32\
        );

    \I__1560\ : InMux
    port map (
            O => \N__10964\,
            I => \N__10961\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__10961\,
            I => \c0.n4579\
        );

    \I__1558\ : InMux
    port map (
            O => \N__10958\,
            I => \N__10955\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__10955\,
            I => n1707
        );

    \I__1556\ : InMux
    port map (
            O => \N__10952\,
            I => \N__10949\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__10949\,
            I => n1768
        );

    \I__1554\ : InMux
    port map (
            O => \N__10946\,
            I => \N__10942\
        );

    \I__1553\ : InMux
    port map (
            O => \N__10945\,
            I => \N__10939\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__10942\,
            I => \c0.tx2.r_Clock_Count_0\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__10939\,
            I => \c0.tx2.r_Clock_Count_0\
        );

    \I__1550\ : InMux
    port map (
            O => \N__10934\,
            I => \N__10929\
        );

    \I__1549\ : InMux
    port map (
            O => \N__10933\,
            I => \N__10926\
        );

    \I__1548\ : InMux
    port map (
            O => \N__10932\,
            I => \N__10923\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__10929\,
            I => \c0.tx2.r_Clock_Count_2\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__10926\,
            I => \c0.tx2.r_Clock_Count_2\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__10923\,
            I => \c0.tx2.r_Clock_Count_2\
        );

    \I__1544\ : InMux
    port map (
            O => \N__10916\,
            I => \N__10911\
        );

    \I__1543\ : InMux
    port map (
            O => \N__10915\,
            I => \N__10908\
        );

    \I__1542\ : InMux
    port map (
            O => \N__10914\,
            I => \N__10905\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__10911\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__10908\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__10905\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__10898\,
            I => \N__10893\
        );

    \I__1537\ : InMux
    port map (
            O => \N__10897\,
            I => \N__10890\
        );

    \I__1536\ : InMux
    port map (
            O => \N__10896\,
            I => \N__10887\
        );

    \I__1535\ : InMux
    port map (
            O => \N__10893\,
            I => \N__10884\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__10890\,
            I => \c0.tx2.r_Clock_Count_1\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__10887\,
            I => \c0.tx2.r_Clock_Count_1\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__10884\,
            I => \c0.tx2.r_Clock_Count_1\
        );

    \I__1531\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10872\
        );

    \I__1530\ : InMux
    port map (
            O => \N__10876\,
            I => \N__10869\
        );

    \I__1529\ : InMux
    port map (
            O => \N__10875\,
            I => \N__10866\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__10872\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__10869\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__10866\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__10859\,
            I => \c0.tx2.n5_cascade_\
        );

    \I__1524\ : InMux
    port map (
            O => \N__10856\,
            I => \N__10853\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__10853\,
            I => n1701
        );

    \I__1522\ : InMux
    port map (
            O => \N__10850\,
            I => \N__10845\
        );

    \I__1521\ : InMux
    port map (
            O => \N__10849\,
            I => \N__10842\
        );

    \I__1520\ : InMux
    port map (
            O => \N__10848\,
            I => \N__10839\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__10845\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__10842\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__10839\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__10832\,
            I => \N__10829\
        );

    \I__1515\ : InMux
    port map (
            O => \N__10829\,
            I => \N__10826\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__10826\,
            I => n1692
        );

    \I__1513\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10818\
        );

    \I__1512\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10815\
        );

    \I__1511\ : InMux
    port map (
            O => \N__10821\,
            I => \N__10812\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__10818\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__10815\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__10812\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__10805\,
            I => \r_SM_Main_2_N_759_1_cascade_\
        );

    \I__1506\ : InMux
    port map (
            O => \N__10802\,
            I => \N__10794\
        );

    \I__1505\ : InMux
    port map (
            O => \N__10801\,
            I => \N__10791\
        );

    \I__1504\ : InMux
    port map (
            O => \N__10800\,
            I => \N__10788\
        );

    \I__1503\ : InMux
    port map (
            O => \N__10799\,
            I => \N__10785\
        );

    \I__1502\ : InMux
    port map (
            O => \N__10798\,
            I => \N__10780\
        );

    \I__1501\ : InMux
    port map (
            O => \N__10797\,
            I => \N__10780\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__10794\,
            I => \c0.tx2.r_Clock_Count_8\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__10791\,
            I => \c0.tx2.r_Clock_Count_8\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__10788\,
            I => \c0.tx2.r_Clock_Count_8\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__10785\,
            I => \c0.tx2.r_Clock_Count_8\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__10780\,
            I => \c0.tx2.r_Clock_Count_8\
        );

    \I__1495\ : InMux
    port map (
            O => \N__10769\,
            I => \N__10763\
        );

    \I__1494\ : InMux
    port map (
            O => \N__10768\,
            I => \N__10760\
        );

    \I__1493\ : InMux
    port map (
            O => \N__10767\,
            I => \N__10755\
        );

    \I__1492\ : InMux
    port map (
            O => \N__10766\,
            I => \N__10755\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__10763\,
            I => \c0.tx2.n2902\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__10760\,
            I => \c0.tx2.n2902\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__10755\,
            I => \c0.tx2.n2902\
        );

    \I__1488\ : InMux
    port map (
            O => \N__10748\,
            I => \N__10745\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__10745\,
            I => n4_adj_965
        );

    \I__1486\ : InMux
    port map (
            O => \N__10742\,
            I => \c0.tx2.n3892\
        );

    \I__1485\ : InMux
    port map (
            O => \N__10739\,
            I => \c0.tx2.n3893\
        );

    \I__1484\ : InMux
    port map (
            O => \N__10736\,
            I => \c0.tx2.n3894\
        );

    \I__1483\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10730\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__10730\,
            I => n1698
        );

    \I__1481\ : InMux
    port map (
            O => \N__10727\,
            I => \c0.tx2.n3895\
        );

    \I__1480\ : InMux
    port map (
            O => \N__10724\,
            I => \c0.tx2.n3896\
        );

    \I__1479\ : InMux
    port map (
            O => \N__10721\,
            I => \c0.tx2.n3897\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10718\,
            I => \bfn_4_22_0_\
        );

    \I__1477\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10712\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__10712\,
            I => n1689
        );

    \I__1475\ : InMux
    port map (
            O => \N__10709\,
            I => \N__10706\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__10706\,
            I => \N__10703\
        );

    \I__1473\ : Odrv4
    port map (
            O => \N__10703\,
            I => n1704
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__10700\,
            I => \N__10696\
        );

    \I__1471\ : InMux
    port map (
            O => \N__10699\,
            I => \N__10693\
        );

    \I__1470\ : InMux
    port map (
            O => \N__10696\,
            I => \N__10690\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__10693\,
            I => rx_data_3
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__10690\,
            I => rx_data_3
        );

    \I__1467\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10681\
        );

    \I__1466\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10677\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__10681\,
            I => \N__10674\
        );

    \I__1464\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10671\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__10677\,
            I => data_in_0_1
        );

    \I__1462\ : Odrv4
    port map (
            O => \N__10674\,
            I => data_in_0_1
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__10671\,
            I => data_in_0_1
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__10664\,
            I => \N__10661\
        );

    \I__1459\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10658\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__10658\,
            I => \N__10655\
        );

    \I__1457\ : Span4Mux_s2_h
    port map (
            O => \N__10655\,
            I => \N__10650\
        );

    \I__1456\ : InMux
    port map (
            O => \N__10654\,
            I => \N__10645\
        );

    \I__1455\ : InMux
    port map (
            O => \N__10653\,
            I => \N__10645\
        );

    \I__1454\ : Odrv4
    port map (
            O => \N__10650\,
            I => data_in_5_5
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__10645\,
            I => data_in_5_5
        );

    \I__1452\ : InMux
    port map (
            O => \N__10640\,
            I => \N__10637\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__10637\,
            I => \N__10633\
        );

    \I__1450\ : InMux
    port map (
            O => \N__10636\,
            I => \N__10630\
        );

    \I__1449\ : Span4Mux_v
    port map (
            O => \N__10633\,
            I => \N__10625\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__10630\,
            I => \N__10625\
        );

    \I__1447\ : Span4Mux_v
    port map (
            O => \N__10625\,
            I => \N__10622\
        );

    \I__1446\ : Span4Mux_s1_h
    port map (
            O => \N__10622\,
            I => \N__10618\
        );

    \I__1445\ : InMux
    port map (
            O => \N__10621\,
            I => \N__10615\
        );

    \I__1444\ : Odrv4
    port map (
            O => \N__10618\,
            I => data_in_4_5
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__10615\,
            I => data_in_4_5
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__10610\,
            I => \c0.rx.n4873_cascade_\
        );

    \I__1441\ : InMux
    port map (
            O => \N__10607\,
            I => \N__10604\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__10604\,
            I => \N__10599\
        );

    \I__1439\ : InMux
    port map (
            O => \N__10603\,
            I => \N__10595\
        );

    \I__1438\ : InMux
    port map (
            O => \N__10602\,
            I => \N__10592\
        );

    \I__1437\ : Span4Mux_s3_h
    port map (
            O => \N__10599\,
            I => \N__10589\
        );

    \I__1436\ : InMux
    port map (
            O => \N__10598\,
            I => \N__10586\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__10595\,
            I => data_in_3_7
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__10592\,
            I => data_in_3_7
        );

    \I__1433\ : Odrv4
    port map (
            O => \N__10589\,
            I => data_in_3_7
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__10586\,
            I => data_in_3_7
        );

    \I__1431\ : InMux
    port map (
            O => \N__10577\,
            I => \N__10574\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__10574\,
            I => \N__10569\
        );

    \I__1429\ : InMux
    port map (
            O => \N__10573\,
            I => \N__10566\
        );

    \I__1428\ : InMux
    port map (
            O => \N__10572\,
            I => \N__10563\
        );

    \I__1427\ : Odrv4
    port map (
            O => \N__10569\,
            I => data_in_4_1
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__10566\,
            I => data_in_4_1
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__10563\,
            I => data_in_4_1
        );

    \I__1424\ : InMux
    port map (
            O => \N__10556\,
            I => \N__10553\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__10553\,
            I => \N__10549\
        );

    \I__1422\ : InMux
    port map (
            O => \N__10552\,
            I => \N__10546\
        );

    \I__1421\ : Span4Mux_v
    port map (
            O => \N__10549\,
            I => \N__10542\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__10546\,
            I => \N__10539\
        );

    \I__1419\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10535\
        );

    \I__1418\ : Span4Mux_s0_h
    port map (
            O => \N__10542\,
            I => \N__10532\
        );

    \I__1417\ : Span4Mux_v
    port map (
            O => \N__10539\,
            I => \N__10529\
        );

    \I__1416\ : InMux
    port map (
            O => \N__10538\,
            I => \N__10526\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__10535\,
            I => data_in_3_1
        );

    \I__1414\ : Odrv4
    port map (
            O => \N__10532\,
            I => data_in_3_1
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__10529\,
            I => data_in_3_1
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__10526\,
            I => data_in_3_1
        );

    \I__1411\ : InMux
    port map (
            O => \N__10517\,
            I => \bfn_4_21_0_\
        );

    \I__1410\ : InMux
    port map (
            O => \N__10514\,
            I => \N__10511\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__10511\,
            I => n1710
        );

    \I__1408\ : InMux
    port map (
            O => \N__10508\,
            I => \c0.tx2.n3891\
        );

    \I__1407\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10500\
        );

    \I__1406\ : InMux
    port map (
            O => \N__10504\,
            I => \N__10496\
        );

    \I__1405\ : InMux
    port map (
            O => \N__10503\,
            I => \N__10493\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__10500\,
            I => \N__10490\
        );

    \I__1403\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10487\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__10496\,
            I => data_in_2_1
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__10493\,
            I => data_in_2_1
        );

    \I__1400\ : Odrv4
    port map (
            O => \N__10490\,
            I => data_in_2_1
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__10487\,
            I => data_in_2_1
        );

    \I__1398\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10475\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__10475\,
            I => \N__10471\
        );

    \I__1396\ : InMux
    port map (
            O => \N__10474\,
            I => \N__10467\
        );

    \I__1395\ : Span4Mux_v
    port map (
            O => \N__10471\,
            I => \N__10464\
        );

    \I__1394\ : InMux
    port map (
            O => \N__10470\,
            I => \N__10461\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__10467\,
            I => \c0.data_in_field_17\
        );

    \I__1392\ : Odrv4
    port map (
            O => \N__10464\,
            I => \c0.data_in_field_17\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__10461\,
            I => \c0.data_in_field_17\
        );

    \I__1390\ : InMux
    port map (
            O => \N__10454\,
            I => \N__10451\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__10451\,
            I => \N__10447\
        );

    \I__1388\ : InMux
    port map (
            O => \N__10450\,
            I => \N__10442\
        );

    \I__1387\ : Span4Mux_h
    port map (
            O => \N__10447\,
            I => \N__10439\
        );

    \I__1386\ : InMux
    port map (
            O => \N__10446\,
            I => \N__10436\
        );

    \I__1385\ : InMux
    port map (
            O => \N__10445\,
            I => \N__10433\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__10442\,
            I => \c0.data_in_field_15\
        );

    \I__1383\ : Odrv4
    port map (
            O => \N__10439\,
            I => \c0.data_in_field_15\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__10436\,
            I => \c0.data_in_field_15\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__10433\,
            I => \c0.data_in_field_15\
        );

    \I__1380\ : CascadeMux
    port map (
            O => \N__10424\,
            I => \N__10419\
        );

    \I__1379\ : InMux
    port map (
            O => \N__10423\,
            I => \N__10416\
        );

    \I__1378\ : CascadeMux
    port map (
            O => \N__10422\,
            I => \N__10413\
        );

    \I__1377\ : InMux
    port map (
            O => \N__10419\,
            I => \N__10410\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__10416\,
            I => \N__10407\
        );

    \I__1375\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10404\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__10410\,
            I => \c0.data_in_field_27\
        );

    \I__1373\ : Odrv4
    port map (
            O => \N__10407\,
            I => \c0.data_in_field_27\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__10404\,
            I => \c0.data_in_field_27\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__10397\,
            I => \N__10394\
        );

    \I__1370\ : InMux
    port map (
            O => \N__10394\,
            I => \N__10391\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__10391\,
            I => \N__10388\
        );

    \I__1368\ : Span4Mux_s3_h
    port map (
            O => \N__10388\,
            I => \N__10385\
        );

    \I__1367\ : Odrv4
    port map (
            O => \N__10385\,
            I => \c0.n4547\
        );

    \I__1366\ : InMux
    port map (
            O => \N__10382\,
            I => \N__10379\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__10379\,
            I => \N__10376\
        );

    \I__1364\ : Span4Mux_h
    port map (
            O => \N__10376\,
            I => \N__10371\
        );

    \I__1363\ : InMux
    port map (
            O => \N__10375\,
            I => \N__10368\
        );

    \I__1362\ : InMux
    port map (
            O => \N__10374\,
            I => \N__10365\
        );

    \I__1361\ : Odrv4
    port map (
            O => \N__10371\,
            I => data_in_0_3
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__10368\,
            I => data_in_0_3
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__10365\,
            I => data_in_0_3
        );

    \I__1358\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10354\
        );

    \I__1357\ : InMux
    port map (
            O => \N__10357\,
            I => \N__10351\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__10354\,
            I => \N__10346\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__10351\,
            I => \N__10346\
        );

    \I__1354\ : Odrv4
    port map (
            O => \N__10346\,
            I => \c0.data_in_frame_7_5\
        );

    \I__1353\ : InMux
    port map (
            O => \N__10343\,
            I => \N__10338\
        );

    \I__1352\ : InMux
    port map (
            O => \N__10342\,
            I => \N__10335\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10341\,
            I => \N__10332\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__10338\,
            I => \N__10323\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__10335\,
            I => \N__10323\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__10332\,
            I => \N__10323\
        );

    \I__1347\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10318\
        );

    \I__1346\ : InMux
    port map (
            O => \N__10330\,
            I => \N__10318\
        );

    \I__1345\ : Odrv12
    port map (
            O => \N__10323\,
            I => \c0.data_in_field_34\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__10318\,
            I => \c0.data_in_field_34\
        );

    \I__1343\ : InMux
    port map (
            O => \N__10313\,
            I => \N__10310\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__10310\,
            I => \N__10306\
        );

    \I__1341\ : InMux
    port map (
            O => \N__10309\,
            I => \N__10303\
        );

    \I__1340\ : Span4Mux_v
    port map (
            O => \N__10306\,
            I => \N__10296\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__10303\,
            I => \N__10296\
        );

    \I__1338\ : InMux
    port map (
            O => \N__10302\,
            I => \N__10290\
        );

    \I__1337\ : InMux
    port map (
            O => \N__10301\,
            I => \N__10290\
        );

    \I__1336\ : Span4Mux_v
    port map (
            O => \N__10296\,
            I => \N__10287\
        );

    \I__1335\ : InMux
    port map (
            O => \N__10295\,
            I => \N__10284\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__10290\,
            I => \c0.data_in_field_3\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__10287\,
            I => \c0.data_in_field_3\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__10284\,
            I => \c0.data_in_field_3\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__10277\,
            I => \N__10272\
        );

    \I__1330\ : InMux
    port map (
            O => \N__10276\,
            I => \N__10267\
        );

    \I__1329\ : InMux
    port map (
            O => \N__10275\,
            I => \N__10267\
        );

    \I__1328\ : InMux
    port map (
            O => \N__10272\,
            I => \N__10263\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__10267\,
            I => \N__10260\
        );

    \I__1326\ : InMux
    port map (
            O => \N__10266\,
            I => \N__10257\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__10263\,
            I => \c0.data_in_field_19\
        );

    \I__1324\ : Odrv12
    port map (
            O => \N__10260\,
            I => \c0.data_in_field_19\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__10257\,
            I => \c0.data_in_field_19\
        );

    \I__1322\ : InMux
    port map (
            O => \N__10250\,
            I => \N__10247\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__10247\,
            I => \N__10244\
        );

    \I__1320\ : Odrv12
    port map (
            O => \N__10244\,
            I => \c0.n10\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__10241\,
            I => \N__10237\
        );

    \I__1318\ : InMux
    port map (
            O => \N__10240\,
            I => \N__10234\
        );

    \I__1317\ : InMux
    port map (
            O => \N__10237\,
            I => \N__10229\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__10234\,
            I => \N__10226\
        );

    \I__1315\ : InMux
    port map (
            O => \N__10233\,
            I => \N__10223\
        );

    \I__1314\ : InMux
    port map (
            O => \N__10232\,
            I => \N__10220\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__10229\,
            I => \c0.data_in_field_29\
        );

    \I__1312\ : Odrv12
    port map (
            O => \N__10226\,
            I => \c0.data_in_field_29\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__10223\,
            I => \c0.data_in_field_29\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__10220\,
            I => \c0.data_in_field_29\
        );

    \I__1309\ : InMux
    port map (
            O => \N__10211\,
            I => \N__10208\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__10208\,
            I => \c0.n4411\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__10205\,
            I => \c0.n4411_cascade_\
        );

    \I__1306\ : CascadeMux
    port map (
            O => \N__10202\,
            I => \N__10199\
        );

    \I__1305\ : InMux
    port map (
            O => \N__10199\,
            I => \N__10193\
        );

    \I__1304\ : InMux
    port map (
            O => \N__10198\,
            I => \N__10193\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__10193\,
            I => \c0.data_in_frame_6_5\
        );

    \I__1302\ : InMux
    port map (
            O => \N__10190\,
            I => \N__10187\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__10187\,
            I => \N__10184\
        );

    \I__1300\ : Span4Mux_s3_h
    port map (
            O => \N__10184\,
            I => \N__10181\
        );

    \I__1299\ : Odrv4
    port map (
            O => \N__10181\,
            I => \c0.n4595\
        );

    \I__1298\ : CascadeMux
    port map (
            O => \N__10178\,
            I => \c0.n1340_cascade_\
        );

    \I__1297\ : InMux
    port map (
            O => \N__10175\,
            I => \N__10170\
        );

    \I__1296\ : InMux
    port map (
            O => \N__10174\,
            I => \N__10167\
        );

    \I__1295\ : InMux
    port map (
            O => \N__10173\,
            I => \N__10164\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__10170\,
            I => \N__10160\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__10167\,
            I => \N__10155\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__10164\,
            I => \N__10155\
        );

    \I__1291\ : InMux
    port map (
            O => \N__10163\,
            I => \N__10151\
        );

    \I__1290\ : Span4Mux_v
    port map (
            O => \N__10160\,
            I => \N__10148\
        );

    \I__1289\ : Span4Mux_v
    port map (
            O => \N__10155\,
            I => \N__10145\
        );

    \I__1288\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10142\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__10151\,
            I => \c0.data_in_field_16\
        );

    \I__1286\ : Odrv4
    port map (
            O => \N__10148\,
            I => \c0.data_in_field_16\
        );

    \I__1285\ : Odrv4
    port map (
            O => \N__10145\,
            I => \c0.data_in_field_16\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__10142\,
            I => \c0.data_in_field_16\
        );

    \I__1283\ : CascadeMux
    port map (
            O => \N__10133\,
            I => \N__10127\
        );

    \I__1282\ : InMux
    port map (
            O => \N__10132\,
            I => \N__10124\
        );

    \I__1281\ : InMux
    port map (
            O => \N__10131\,
            I => \N__10121\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__10130\,
            I => \N__10116\
        );

    \I__1279\ : InMux
    port map (
            O => \N__10127\,
            I => \N__10113\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__10124\,
            I => \N__10108\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__10121\,
            I => \N__10108\
        );

    \I__1276\ : InMux
    port map (
            O => \N__10120\,
            I => \N__10105\
        );

    \I__1275\ : InMux
    port map (
            O => \N__10119\,
            I => \N__10100\
        );

    \I__1274\ : InMux
    port map (
            O => \N__10116\,
            I => \N__10100\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__10113\,
            I => \c0.data_in_field_33\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__10108\,
            I => \c0.data_in_field_33\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__10105\,
            I => \c0.data_in_field_33\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__10100\,
            I => \c0.data_in_field_33\
        );

    \I__1269\ : InMux
    port map (
            O => \N__10091\,
            I => \N__10088\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__10088\,
            I => \N__10082\
        );

    \I__1267\ : InMux
    port map (
            O => \N__10087\,
            I => \N__10079\
        );

    \I__1266\ : InMux
    port map (
            O => \N__10086\,
            I => \N__10076\
        );

    \I__1265\ : InMux
    port map (
            O => \N__10085\,
            I => \N__10073\
        );

    \I__1264\ : Span4Mux_h
    port map (
            O => \N__10082\,
            I => \N__10066\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__10079\,
            I => \N__10066\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__10076\,
            I => \N__10066\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__10073\,
            I => data_in_2_2
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__10066\,
            I => data_in_2_2
        );

    \I__1259\ : InMux
    port map (
            O => \N__10061\,
            I => \N__10057\
        );

    \I__1258\ : InMux
    port map (
            O => \N__10060\,
            I => \N__10054\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__10057\,
            I => \N__10049\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__10054\,
            I => \N__10046\
        );

    \I__1255\ : InMux
    port map (
            O => \N__10053\,
            I => \N__10041\
        );

    \I__1254\ : InMux
    port map (
            O => \N__10052\,
            I => \N__10041\
        );

    \I__1253\ : Odrv12
    port map (
            O => \N__10049\,
            I => \c0.data_in_field_18\
        );

    \I__1252\ : Odrv4
    port map (
            O => \N__10046\,
            I => \c0.data_in_field_18\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__10041\,
            I => \c0.data_in_field_18\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__10034\,
            I => \c0.n4429_cascade_\
        );

    \I__1249\ : InMux
    port map (
            O => \N__10031\,
            I => \N__10028\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__10028\,
            I => \c0.n4429\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__10025\,
            I => \N__10022\
        );

    \I__1246\ : InMux
    port map (
            O => \N__10022\,
            I => \N__10015\
        );

    \I__1245\ : InMux
    port map (
            O => \N__10021\,
            I => \N__10012\
        );

    \I__1244\ : InMux
    port map (
            O => \N__10020\,
            I => \N__10009\
        );

    \I__1243\ : InMux
    port map (
            O => \N__10019\,
            I => \N__10006\
        );

    \I__1242\ : InMux
    port map (
            O => \N__10018\,
            I => \N__10003\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__10015\,
            I => \c0.data_in_field_46\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__10012\,
            I => \c0.data_in_field_46\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__10009\,
            I => \c0.data_in_field_46\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__10006\,
            I => \c0.data_in_field_46\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__10003\,
            I => \c0.data_in_field_46\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__9992\,
            I => \N__9989\
        );

    \I__1235\ : InMux
    port map (
            O => \N__9989\,
            I => \N__9986\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__9986\,
            I => \N__9983\
        );

    \I__1233\ : Odrv4
    port map (
            O => \N__9983\,
            I => \c0.n6_adj_877\
        );

    \I__1232\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9974\
        );

    \I__1231\ : InMux
    port map (
            O => \N__9979\,
            I => \N__9971\
        );

    \I__1230\ : InMux
    port map (
            O => \N__9978\,
            I => \N__9968\
        );

    \I__1229\ : InMux
    port map (
            O => \N__9977\,
            I => \N__9965\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__9974\,
            I => \c0.data_in_field_5\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__9971\,
            I => \c0.data_in_field_5\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__9968\,
            I => \c0.data_in_field_5\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__9965\,
            I => \c0.data_in_field_5\
        );

    \I__1224\ : InMux
    port map (
            O => \N__9956\,
            I => \N__9953\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__9953\,
            I => \c0.n4450\
        );

    \I__1222\ : InMux
    port map (
            O => \N__9950\,
            I => \N__9947\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__9947\,
            I => \N__9944\
        );

    \I__1220\ : Span4Mux_v
    port map (
            O => \N__9944\,
            I => \N__9939\
        );

    \I__1219\ : InMux
    port map (
            O => \N__9943\,
            I => \N__9934\
        );

    \I__1218\ : InMux
    port map (
            O => \N__9942\,
            I => \N__9934\
        );

    \I__1217\ : Odrv4
    port map (
            O => \N__9939\,
            I => data_in_0_4
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__9934\,
            I => data_in_0_4
        );

    \I__1215\ : InMux
    port map (
            O => \N__9929\,
            I => \N__9925\
        );

    \I__1214\ : InMux
    port map (
            O => \N__9928\,
            I => \N__9922\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__9925\,
            I => \N__9914\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__9922\,
            I => \N__9914\
        );

    \I__1211\ : InMux
    port map (
            O => \N__9921\,
            I => \N__9909\
        );

    \I__1210\ : InMux
    port map (
            O => \N__9920\,
            I => \N__9909\
        );

    \I__1209\ : InMux
    port map (
            O => \N__9919\,
            I => \N__9906\
        );

    \I__1208\ : Odrv4
    port map (
            O => \N__9914\,
            I => \c0.data_in_field_31\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__9909\,
            I => \c0.data_in_field_31\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__9906\,
            I => \c0.data_in_field_31\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__9899\,
            I => \c0.n1261_cascade_\
        );

    \I__1204\ : InMux
    port map (
            O => \N__9896\,
            I => \N__9891\
        );

    \I__1203\ : InMux
    port map (
            O => \N__9895\,
            I => \N__9888\
        );

    \I__1202\ : InMux
    port map (
            O => \N__9894\,
            I => \N__9884\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__9891\,
            I => \N__9881\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__9888\,
            I => \N__9878\
        );

    \I__1199\ : InMux
    port map (
            O => \N__9887\,
            I => \N__9875\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__9884\,
            I => \c0.data_in_field_6\
        );

    \I__1197\ : Odrv12
    port map (
            O => \N__9881\,
            I => \c0.data_in_field_6\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__9878\,
            I => \c0.data_in_field_6\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__9875\,
            I => \c0.data_in_field_6\
        );

    \I__1194\ : InMux
    port map (
            O => \N__9866\,
            I => \N__9862\
        );

    \I__1193\ : InMux
    port map (
            O => \N__9865\,
            I => \N__9859\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__9862\,
            I => \c0.n1284\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__9859\,
            I => \c0.n1284\
        );

    \I__1190\ : CascadeMux
    port map (
            O => \N__9854\,
            I => \c0.n4408_cascade_\
        );

    \I__1189\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9847\
        );

    \I__1188\ : InMux
    port map (
            O => \N__9850\,
            I => \N__9844\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__9847\,
            I => \c0.n4468\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__9844\,
            I => \c0.n4468\
        );

    \I__1185\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9836\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__9836\,
            I => \N__9833\
        );

    \I__1183\ : Span4Mux_h
    port map (
            O => \N__9833\,
            I => \N__9830\
        );

    \I__1182\ : Span4Mux_v
    port map (
            O => \N__9830\,
            I => \N__9824\
        );

    \I__1181\ : InMux
    port map (
            O => \N__9829\,
            I => \N__9819\
        );

    \I__1180\ : InMux
    port map (
            O => \N__9828\,
            I => \N__9819\
        );

    \I__1179\ : InMux
    port map (
            O => \N__9827\,
            I => \N__9816\
        );

    \I__1178\ : Odrv4
    port map (
            O => \N__9824\,
            I => data_in_2_3
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__9819\,
            I => data_in_2_3
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__9816\,
            I => data_in_2_3
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__9809\,
            I => \N__9805\
        );

    \I__1174\ : InMux
    port map (
            O => \N__9808\,
            I => \N__9802\
        );

    \I__1173\ : InMux
    port map (
            O => \N__9805\,
            I => \N__9797\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__9802\,
            I => \N__9794\
        );

    \I__1171\ : InMux
    port map (
            O => \N__9801\,
            I => \N__9789\
        );

    \I__1170\ : InMux
    port map (
            O => \N__9800\,
            I => \N__9789\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__9797\,
            I => \N__9786\
        );

    \I__1168\ : Span4Mux_h
    port map (
            O => \N__9794\,
            I => \N__9783\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__9789\,
            I => data_in_3_2
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__9786\,
            I => data_in_3_2
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__9783\,
            I => data_in_3_2
        );

    \I__1164\ : InMux
    port map (
            O => \N__9776\,
            I => \N__9773\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__9773\,
            I => \N__9768\
        );

    \I__1162\ : InMux
    port map (
            O => \N__9772\,
            I => \N__9765\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__9771\,
            I => \N__9761\
        );

    \I__1160\ : Span4Mux_h
    port map (
            O => \N__9768\,
            I => \N__9756\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__9765\,
            I => \N__9756\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9764\,
            I => \N__9751\
        );

    \I__1157\ : InMux
    port map (
            O => \N__9761\,
            I => \N__9751\
        );

    \I__1156\ : Odrv4
    port map (
            O => \N__9756\,
            I => data_in_2_5
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__9751\,
            I => data_in_2_5
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__9746\,
            I => \c0.n1271_cascade_\
        );

    \I__1153\ : InMux
    port map (
            O => \N__9743\,
            I => \N__9738\
        );

    \I__1152\ : InMux
    port map (
            O => \N__9742\,
            I => \N__9733\
        );

    \I__1151\ : InMux
    port map (
            O => \N__9741\,
            I => \N__9733\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__9738\,
            I => \c0.data_in_field_22\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__9733\,
            I => \c0.data_in_field_22\
        );

    \I__1148\ : InMux
    port map (
            O => \N__9728\,
            I => \N__9725\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__9725\,
            I => \N__9722\
        );

    \I__1146\ : Span4Mux_v
    port map (
            O => \N__9722\,
            I => \N__9719\
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__9719\,
            I => \c0.n4556\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__9716\,
            I => \c0.n10_adj_874_cascade_\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9713\,
            I => \N__9710\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__9710\,
            I => \N__9707\
        );

    \I__1141\ : Odrv4
    port map (
            O => \N__9707\,
            I => \c0.n4567\
        );

    \I__1140\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9701\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__9701\,
            I => \N__9698\
        );

    \I__1138\ : Span4Mux_v
    port map (
            O => \N__9698\,
            I => \N__9693\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__9697\,
            I => \N__9690\
        );

    \I__1136\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9687\
        );

    \I__1135\ : Span4Mux_h
    port map (
            O => \N__9693\,
            I => \N__9684\
        );

    \I__1134\ : InMux
    port map (
            O => \N__9690\,
            I => \N__9681\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__9687\,
            I => data_in_0_7
        );

    \I__1132\ : Odrv4
    port map (
            O => \N__9684\,
            I => data_in_0_7
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__9681\,
            I => data_in_0_7
        );

    \I__1130\ : InMux
    port map (
            O => \N__9674\,
            I => \N__9671\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__9671\,
            I => \c0.n4541\
        );

    \I__1128\ : InMux
    port map (
            O => \N__9668\,
            I => \N__9665\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__9665\,
            I => \N__9662\
        );

    \I__1126\ : Odrv12
    port map (
            O => \N__9662\,
            I => \c0.n4544\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__9659\,
            I => \n4512_cascade_\
        );

    \I__1124\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9653\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__9653\,
            I => \N__9650\
        );

    \I__1122\ : Span4Mux_v
    port map (
            O => \N__9650\,
            I => \N__9647\
        );

    \I__1121\ : Odrv4
    port map (
            O => \N__9647\,
            I => \c0.n4546\
        );

    \I__1120\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9641\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__9641\,
            I => \c0.n4603\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__9638\,
            I => \N__9634\
        );

    \I__1117\ : InMux
    port map (
            O => \N__9637\,
            I => \N__9626\
        );

    \I__1116\ : InMux
    port map (
            O => \N__9634\,
            I => \N__9626\
        );

    \I__1115\ : InMux
    port map (
            O => \N__9633\,
            I => \N__9626\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__9626\,
            I => n1611
        );

    \I__1113\ : CascadeMux
    port map (
            O => \N__9623\,
            I => \n2326_cascade_\
        );

    \I__1112\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9617\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__9617\,
            I => n4514
        );

    \I__1110\ : InMux
    port map (
            O => \N__9614\,
            I => \N__9605\
        );

    \I__1109\ : InMux
    port map (
            O => \N__9613\,
            I => \N__9605\
        );

    \I__1108\ : InMux
    port map (
            O => \N__9612\,
            I => \N__9605\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__9605\,
            I => n4512
        );

    \I__1106\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9599\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__9599\,
            I => \N__9596\
        );

    \I__1104\ : Span4Mux_v
    port map (
            O => \N__9596\,
            I => \N__9593\
        );

    \I__1103\ : Odrv4
    port map (
            O => \N__9593\,
            I => n4523
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__9590\,
            I => \n4522_cascade_\
        );

    \I__1101\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9584\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__9584\,
            I => n4777
        );

    \I__1099\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9576\
        );

    \I__1098\ : InMux
    port map (
            O => \N__9580\,
            I => \N__9569\
        );

    \I__1097\ : InMux
    port map (
            O => \N__9579\,
            I => \N__9569\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__9576\,
            I => \N__9566\
        );

    \I__1095\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9563\
        );

    \I__1094\ : InMux
    port map (
            O => \N__9574\,
            I => \N__9560\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__9569\,
            I => \r_Bit_Index_1\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__9566\,
            I => \r_Bit_Index_1\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__9563\,
            I => \r_Bit_Index_1\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__9560\,
            I => \r_Bit_Index_1\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__9551\,
            I => \N__9545\
        );

    \I__1088\ : InMux
    port map (
            O => \N__9550\,
            I => \N__9539\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__9549\,
            I => \N__9536\
        );

    \I__1086\ : InMux
    port map (
            O => \N__9548\,
            I => \N__9533\
        );

    \I__1085\ : InMux
    port map (
            O => \N__9545\,
            I => \N__9528\
        );

    \I__1084\ : InMux
    port map (
            O => \N__9544\,
            I => \N__9528\
        );

    \I__1083\ : InMux
    port map (
            O => \N__9543\,
            I => \N__9523\
        );

    \I__1082\ : InMux
    port map (
            O => \N__9542\,
            I => \N__9523\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__9539\,
            I => \N__9520\
        );

    \I__1080\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9517\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__9533\,
            I => \r_Bit_Index_0_adj_956\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__9528\,
            I => \r_Bit_Index_0_adj_956\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__9523\,
            I => \r_Bit_Index_0_adj_956\
        );

    \I__1076\ : Odrv4
    port map (
            O => \N__9520\,
            I => \r_Bit_Index_0_adj_956\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__9517\,
            I => \r_Bit_Index_0_adj_956\
        );

    \I__1074\ : InMux
    port map (
            O => \N__9506\,
            I => \N__9502\
        );

    \I__1073\ : InMux
    port map (
            O => \N__9505\,
            I => \N__9495\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__9502\,
            I => \N__9492\
        );

    \I__1071\ : InMux
    port map (
            O => \N__9501\,
            I => \N__9485\
        );

    \I__1070\ : InMux
    port map (
            O => \N__9500\,
            I => \N__9485\
        );

    \I__1069\ : InMux
    port map (
            O => \N__9499\,
            I => \N__9480\
        );

    \I__1068\ : InMux
    port map (
            O => \N__9498\,
            I => \N__9480\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__9495\,
            I => \N__9475\
        );

    \I__1066\ : Span4Mux_s2_h
    port map (
            O => \N__9492\,
            I => \N__9475\
        );

    \I__1065\ : InMux
    port map (
            O => \N__9491\,
            I => \N__9470\
        );

    \I__1064\ : InMux
    port map (
            O => \N__9490\,
            I => \N__9470\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__9485\,
            I => \r_Bit_Index_2_adj_955\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__9480\,
            I => \r_Bit_Index_2_adj_955\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__9475\,
            I => \r_Bit_Index_2_adj_955\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__9470\,
            I => \r_Bit_Index_2_adj_955\
        );

    \I__1059\ : InMux
    port map (
            O => \N__9461\,
            I => \N__9458\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__9458\,
            I => \N__9455\
        );

    \I__1057\ : Odrv4
    port map (
            O => \N__9455\,
            I => n11_adj_941
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__9452\,
            I => \n4638_cascade_\
        );

    \I__1055\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__9446\,
            I => tx2_done
        );

    \I__1053\ : InMux
    port map (
            O => \N__9443\,
            I => \N__9440\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__9440\,
            I => \c0.n4598\
        );

    \I__1051\ : InMux
    port map (
            O => \N__9437\,
            I => \N__9434\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__9434\,
            I => \c0.n4807\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__9431\,
            I => \tx2_data_2_keep_cascade_\
        );

    \I__1048\ : InMux
    port map (
            O => \N__9428\,
            I => \N__9424\
        );

    \I__1047\ : InMux
    port map (
            O => \N__9427\,
            I => \N__9421\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__9424\,
            I => \r_Tx_Data_2_adj_962\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__9421\,
            I => \r_Tx_Data_2_adj_962\
        );

    \I__1044\ : InMux
    port map (
            O => \N__9416\,
            I => \N__9413\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__9413\,
            I => n9_adj_939
        );

    \I__1042\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9405\
        );

    \I__1041\ : InMux
    port map (
            O => \N__9409\,
            I => \N__9401\
        );

    \I__1040\ : InMux
    port map (
            O => \N__9408\,
            I => \N__9398\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__9405\,
            I => \N__9395\
        );

    \I__1038\ : InMux
    port map (
            O => \N__9404\,
            I => \N__9392\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__9401\,
            I => data_in_2_0
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__9398\,
            I => data_in_2_0
        );

    \I__1035\ : Odrv4
    port map (
            O => \N__9395\,
            I => data_in_2_0
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__9392\,
            I => data_in_2_0
        );

    \I__1033\ : InMux
    port map (
            O => \N__9383\,
            I => \N__9380\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__9380\,
            I => \N__9377\
        );

    \I__1031\ : Odrv4
    port map (
            O => \N__9377\,
            I => \c0.n27\
        );

    \I__1030\ : InMux
    port map (
            O => \N__9374\,
            I => \N__9371\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__9371\,
            I => \c0.rx.r_Rx_Data_R\
        );

    \I__1028\ : InMux
    port map (
            O => \N__9368\,
            I => \N__9363\
        );

    \I__1027\ : InMux
    port map (
            O => \N__9367\,
            I => \N__9360\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__9366\,
            I => \N__9356\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__9363\,
            I => \N__9353\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__9360\,
            I => \N__9350\
        );

    \I__1023\ : InMux
    port map (
            O => \N__9359\,
            I => \N__9345\
        );

    \I__1022\ : InMux
    port map (
            O => \N__9356\,
            I => \N__9345\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__9353\,
            I => data_in_1_4
        );

    \I__1020\ : Odrv4
    port map (
            O => \N__9350\,
            I => data_in_1_4
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__9345\,
            I => data_in_1_4
        );

    \I__1018\ : CascadeMux
    port map (
            O => \N__9338\,
            I => \N__9333\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__9337\,
            I => \N__9329\
        );

    \I__1016\ : InMux
    port map (
            O => \N__9336\,
            I => \N__9326\
        );

    \I__1015\ : InMux
    port map (
            O => \N__9333\,
            I => \N__9323\
        );

    \I__1014\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9320\
        );

    \I__1013\ : InMux
    port map (
            O => \N__9329\,
            I => \N__9317\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__9326\,
            I => \N__9310\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__9323\,
            I => \N__9310\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__9320\,
            I => \N__9310\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__9317\,
            I => data_in_1_7
        );

    \I__1008\ : Odrv4
    port map (
            O => \N__9310\,
            I => data_in_1_7
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__9305\,
            I => \N__9301\
        );

    \I__1006\ : InMux
    port map (
            O => \N__9304\,
            I => \N__9298\
        );

    \I__1005\ : InMux
    port map (
            O => \N__9301\,
            I => \N__9295\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__9298\,
            I => \c0.data_in_frame_7_0\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__9295\,
            I => \c0.data_in_frame_7_0\
        );

    \I__1002\ : CascadeMux
    port map (
            O => \N__9290\,
            I => \N__9286\
        );

    \I__1001\ : InMux
    port map (
            O => \N__9289\,
            I => \N__9283\
        );

    \I__1000\ : InMux
    port map (
            O => \N__9286\,
            I => \N__9280\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__9283\,
            I => \N__9277\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__9280\,
            I => \N__9274\
        );

    \I__997\ : Span4Mux_h
    port map (
            O => \N__9277\,
            I => \N__9269\
        );

    \I__996\ : Span4Mux_v
    port map (
            O => \N__9274\,
            I => \N__9266\
        );

    \I__995\ : InMux
    port map (
            O => \N__9273\,
            I => \N__9261\
        );

    \I__994\ : InMux
    port map (
            O => \N__9272\,
            I => \N__9261\
        );

    \I__993\ : Odrv4
    port map (
            O => \N__9269\,
            I => data_in_2_6
        );

    \I__992\ : Odrv4
    port map (
            O => \N__9266\,
            I => data_in_2_6
        );

    \I__991\ : LocalMux
    port map (
            O => \N__9261\,
            I => data_in_2_6
        );

    \I__990\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9251\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__9251\,
            I => \N__9247\
        );

    \I__988\ : CascadeMux
    port map (
            O => \N__9250\,
            I => \N__9244\
        );

    \I__987\ : Span4Mux_v
    port map (
            O => \N__9247\,
            I => \N__9241\
        );

    \I__986\ : InMux
    port map (
            O => \N__9244\,
            I => \N__9238\
        );

    \I__985\ : Odrv4
    port map (
            O => \N__9241\,
            I => rx_data_2
        );

    \I__984\ : LocalMux
    port map (
            O => \N__9238\,
            I => rx_data_2
        );

    \I__983\ : InMux
    port map (
            O => \N__9233\,
            I => \N__9230\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__9230\,
            I => \PIN_2_c\
        );

    \I__981\ : InMux
    port map (
            O => \N__9227\,
            I => \N__9223\
        );

    \I__980\ : CascadeMux
    port map (
            O => \N__9226\,
            I => \N__9220\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__9223\,
            I => \N__9215\
        );

    \I__978\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9212\
        );

    \I__977\ : InMux
    port map (
            O => \N__9219\,
            I => \N__9209\
        );

    \I__976\ : InMux
    port map (
            O => \N__9218\,
            I => \N__9206\
        );

    \I__975\ : Odrv4
    port map (
            O => \N__9215\,
            I => data_in_1_6
        );

    \I__974\ : LocalMux
    port map (
            O => \N__9212\,
            I => data_in_1_6
        );

    \I__973\ : LocalMux
    port map (
            O => \N__9209\,
            I => data_in_1_6
        );

    \I__972\ : LocalMux
    port map (
            O => \N__9206\,
            I => data_in_1_6
        );

    \I__971\ : InMux
    port map (
            O => \N__9197\,
            I => \N__9194\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__9194\,
            I => \N__9191\
        );

    \I__969\ : Odrv4
    port map (
            O => \N__9191\,
            I => \c0.n26_adj_869\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__9188\,
            I => \N__9185\
        );

    \I__967\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9182\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__9182\,
            I => \N__9177\
        );

    \I__965\ : InMux
    port map (
            O => \N__9181\,
            I => \N__9174\
        );

    \I__964\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9171\
        );

    \I__963\ : Span4Mux_v
    port map (
            O => \N__9177\,
            I => \N__9168\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__9174\,
            I => data_in_0_0
        );

    \I__961\ : LocalMux
    port map (
            O => \N__9171\,
            I => data_in_0_0
        );

    \I__960\ : Odrv4
    port map (
            O => \N__9168\,
            I => data_in_0_0
        );

    \I__959\ : InMux
    port map (
            O => \N__9161\,
            I => \N__9158\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__9158\,
            I => \c0.n30\
        );

    \I__957\ : CascadeMux
    port map (
            O => \N__9155\,
            I => \c0.n25_adj_870_cascade_\
        );

    \I__956\ : InMux
    port map (
            O => \N__9152\,
            I => \N__9149\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__9149\,
            I => \c0.n3933\
        );

    \I__954\ : CascadeMux
    port map (
            O => \N__9146\,
            I => \c0.n1197_cascade_\
        );

    \I__953\ : InMux
    port map (
            O => \N__9143\,
            I => \N__9139\
        );

    \I__952\ : InMux
    port map (
            O => \N__9142\,
            I => \N__9136\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__9139\,
            I => \c0.data_in_frame_6_0\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__9136\,
            I => \c0.data_in_frame_6_0\
        );

    \I__949\ : InMux
    port map (
            O => \N__9131\,
            I => \N__9125\
        );

    \I__948\ : InMux
    port map (
            O => \N__9130\,
            I => \N__9122\
        );

    \I__947\ : InMux
    port map (
            O => \N__9129\,
            I => \N__9119\
        );

    \I__946\ : InMux
    port map (
            O => \N__9128\,
            I => \N__9116\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__9125\,
            I => data_in_3_5
        );

    \I__944\ : LocalMux
    port map (
            O => \N__9122\,
            I => data_in_3_5
        );

    \I__943\ : LocalMux
    port map (
            O => \N__9119\,
            I => data_in_3_5
        );

    \I__942\ : LocalMux
    port map (
            O => \N__9116\,
            I => data_in_3_5
        );

    \I__941\ : InMux
    port map (
            O => \N__9107\,
            I => \N__9104\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__9104\,
            I => \N__9100\
        );

    \I__939\ : InMux
    port map (
            O => \N__9103\,
            I => \N__9096\
        );

    \I__938\ : Span4Mux_v
    port map (
            O => \N__9100\,
            I => \N__9093\
        );

    \I__937\ : InMux
    port map (
            O => \N__9099\,
            I => \N__9090\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__9096\,
            I => data_in_0_6
        );

    \I__935\ : Odrv4
    port map (
            O => \N__9093\,
            I => data_in_0_6
        );

    \I__934\ : LocalMux
    port map (
            O => \N__9090\,
            I => data_in_0_6
        );

    \I__933\ : InMux
    port map (
            O => \N__9083\,
            I => \N__9079\
        );

    \I__932\ : InMux
    port map (
            O => \N__9082\,
            I => \N__9074\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__9079\,
            I => \N__9071\
        );

    \I__930\ : InMux
    port map (
            O => \N__9078\,
            I => \N__9066\
        );

    \I__929\ : InMux
    port map (
            O => \N__9077\,
            I => \N__9066\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__9074\,
            I => \N__9063\
        );

    \I__927\ : Odrv4
    port map (
            O => \N__9071\,
            I => data_in_1_3
        );

    \I__926\ : LocalMux
    port map (
            O => \N__9066\,
            I => data_in_1_3
        );

    \I__925\ : Odrv4
    port map (
            O => \N__9063\,
            I => data_in_1_3
        );

    \I__924\ : InMux
    port map (
            O => \N__9056\,
            I => \N__9051\
        );

    \I__923\ : InMux
    port map (
            O => \N__9055\,
            I => \N__9048\
        );

    \I__922\ : InMux
    port map (
            O => \N__9054\,
            I => \N__9045\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__9051\,
            I => data_in_5_6
        );

    \I__920\ : LocalMux
    port map (
            O => \N__9048\,
            I => data_in_5_6
        );

    \I__919\ : LocalMux
    port map (
            O => \N__9045\,
            I => data_in_5_6
        );

    \I__918\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__9035\,
            I => \c0.n4594\
        );

    \I__916\ : InMux
    port map (
            O => \N__9032\,
            I => \N__9029\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__9029\,
            I => \c0.n4825\
        );

    \I__914\ : InMux
    port map (
            O => \N__9026\,
            I => \N__9023\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__9023\,
            I => \c0.n4813\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__9020\,
            I => \tx2_data_3_keep_cascade_\
        );

    \I__911\ : InMux
    port map (
            O => \N__9017\,
            I => \N__9013\
        );

    \I__910\ : InMux
    port map (
            O => \N__9016\,
            I => \N__9010\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__9013\,
            I => \N__9007\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__9010\,
            I => \r_Tx_Data_3_adj_961\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__9007\,
            I => \r_Tx_Data_3_adj_961\
        );

    \I__906\ : InMux
    port map (
            O => \N__9002\,
            I => \N__8999\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__8999\,
            I => \c0.n4600\
        );

    \I__904\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8993\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__8993\,
            I => \N__8990\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__8990\,
            I => \c0.n4552\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__8987\,
            I => \c0.n4553_cascade_\
        );

    \I__900\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__8981\,
            I => tx2_data_5_keep
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__8978\,
            I => \N__8974\
        );

    \I__897\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8970\
        );

    \I__896\ : InMux
    port map (
            O => \N__8974\,
            I => \N__8967\
        );

    \I__895\ : InMux
    port map (
            O => \N__8973\,
            I => \N__8964\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__8970\,
            I => data_in_0_5
        );

    \I__893\ : LocalMux
    port map (
            O => \N__8967\,
            I => data_in_0_5
        );

    \I__892\ : LocalMux
    port map (
            O => \N__8964\,
            I => data_in_0_5
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__8957\,
            I => \N__8953\
        );

    \I__890\ : InMux
    port map (
            O => \N__8956\,
            I => \N__8949\
        );

    \I__889\ : InMux
    port map (
            O => \N__8953\,
            I => \N__8946\
        );

    \I__888\ : InMux
    port map (
            O => \N__8952\,
            I => \N__8942\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__8949\,
            I => \N__8937\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__8946\,
            I => \N__8937\
        );

    \I__885\ : InMux
    port map (
            O => \N__8945\,
            I => \N__8934\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__8942\,
            I => data_in_1_0
        );

    \I__883\ : Odrv4
    port map (
            O => \N__8937\,
            I => data_in_1_0
        );

    \I__882\ : LocalMux
    port map (
            O => \N__8934\,
            I => data_in_1_0
        );

    \I__881\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8924\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__8924\,
            I => tx2_data_7_keep
        );

    \I__879\ : InMux
    port map (
            O => \N__8921\,
            I => \N__8915\
        );

    \I__878\ : InMux
    port map (
            O => \N__8920\,
            I => \N__8915\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__8915\,
            I => \r_Tx_Data_5_adj_959\
        );

    \I__876\ : InMux
    port map (
            O => \N__8912\,
            I => \N__8909\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__8909\,
            I => n4624
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__8906\,
            I => \c0.n4801_cascade_\
        );

    \I__873\ : CascadeMux
    port map (
            O => \N__8903\,
            I => \tx2_data_1_keep_cascade_\
        );

    \I__872\ : InMux
    port map (
            O => \N__8900\,
            I => \N__8894\
        );

    \I__871\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8894\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__8894\,
            I => \r_Tx_Data_1_adj_963\
        );

    \I__869\ : InMux
    port map (
            O => \N__8891\,
            I => \N__8885\
        );

    \I__868\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8885\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__8885\,
            I => \r_Tx_Data_7_adj_957\
        );

    \I__866\ : InMux
    port map (
            O => \N__8882\,
            I => \N__8879\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__8879\,
            I => n4625
        );

    \I__864\ : InMux
    port map (
            O => \N__8876\,
            I => \N__8873\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__8873\,
            I => \c0.n4540\
        );

    \I__862\ : InMux
    port map (
            O => \N__8870\,
            I => \N__8867\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__8867\,
            I => \c0.n4606\
        );

    \I__860\ : InMux
    port map (
            O => \N__8864\,
            I => \N__8861\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__8861\,
            I => \N__8858\
        );

    \I__858\ : Span4Mux_v
    port map (
            O => \N__8858\,
            I => \N__8854\
        );

    \I__857\ : InMux
    port map (
            O => \N__8857\,
            I => \N__8851\
        );

    \I__856\ : Span4Mux_v
    port map (
            O => \N__8854\,
            I => \N__8848\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__8851\,
            I => \c0.data_in_frame_6_4\
        );

    \I__854\ : Odrv4
    port map (
            O => \N__8848\,
            I => \c0.data_in_frame_6_4\
        );

    \I__853\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8840\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8840\,
            I => \N__8836\
        );

    \I__851\ : InMux
    port map (
            O => \N__8839\,
            I => \N__8833\
        );

    \I__850\ : Span4Mux_h
    port map (
            O => \N__8836\,
            I => \N__8830\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__8833\,
            I => \c0.data_in_frame_7_2\
        );

    \I__848\ : Odrv4
    port map (
            O => \N__8830\,
            I => \c0.data_in_frame_7_2\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__8825\,
            I => \c0.n4604_cascade_\
        );

    \I__846\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8818\
        );

    \I__845\ : InMux
    port map (
            O => \N__8821\,
            I => \N__8815\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__8818\,
            I => \c0.data_in_frame_6_7\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__8815\,
            I => \c0.data_in_frame_6_7\
        );

    \I__842\ : InMux
    port map (
            O => \N__8810\,
            I => \N__8807\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__8807\,
            I => \N__8804\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__8804\,
            I => \c0.n4583\
        );

    \I__839\ : CascadeMux
    port map (
            O => \N__8801\,
            I => \N__8798\
        );

    \I__838\ : InMux
    port map (
            O => \N__8798\,
            I => \N__8792\
        );

    \I__837\ : InMux
    port map (
            O => \N__8797\,
            I => \N__8792\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__8792\,
            I => \N__8789\
        );

    \I__835\ : Odrv4
    port map (
            O => \N__8789\,
            I => \c0.data_in_frame_7_7\
        );

    \I__834\ : InMux
    port map (
            O => \N__8786\,
            I => \N__8782\
        );

    \I__833\ : InMux
    port map (
            O => \N__8785\,
            I => \N__8779\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__8782\,
            I => \c0.data_in_frame_7_4\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__8779\,
            I => \c0.data_in_frame_7_4\
        );

    \I__830\ : InMux
    port map (
            O => \N__8774\,
            I => \N__8771\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__8771\,
            I => \c0.n4555\
        );

    \I__828\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8762\
        );

    \I__827\ : InMux
    port map (
            O => \N__8767\,
            I => \N__8762\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__8762\,
            I => \c0.data_in_frame_6_3\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__8759\,
            I => \N__8755\
        );

    \I__824\ : InMux
    port map (
            O => \N__8758\,
            I => \N__8752\
        );

    \I__823\ : InMux
    port map (
            O => \N__8755\,
            I => \N__8749\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__8752\,
            I => \N__8746\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__8749\,
            I => \c0.data_in_frame_7_6\
        );

    \I__820\ : Odrv12
    port map (
            O => \N__8746\,
            I => \c0.data_in_frame_7_6\
        );

    \I__819\ : InMux
    port map (
            O => \N__8741\,
            I => \N__8738\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__8738\,
            I => \N__8735\
        );

    \I__817\ : Span4Mux_v
    port map (
            O => \N__8735\,
            I => \N__8732\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__8732\,
            I => \c0.n4831\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__8729\,
            I => \tx2_data_6_keep_cascade_\
        );

    \I__814\ : InMux
    port map (
            O => \N__8726\,
            I => \N__8722\
        );

    \I__813\ : InMux
    port map (
            O => \N__8725\,
            I => \N__8719\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__8722\,
            I => \r_Tx_Data_6_adj_958\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__8719\,
            I => \r_Tx_Data_6_adj_958\
        );

    \I__810\ : InMux
    port map (
            O => \N__8714\,
            I => \N__8709\
        );

    \I__809\ : InMux
    port map (
            O => \N__8713\,
            I => \N__8705\
        );

    \I__808\ : InMux
    port map (
            O => \N__8712\,
            I => \N__8702\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__8709\,
            I => \N__8699\
        );

    \I__806\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8696\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__8705\,
            I => data_in_1_5
        );

    \I__804\ : LocalMux
    port map (
            O => \N__8702\,
            I => data_in_1_5
        );

    \I__803\ : Odrv4
    port map (
            O => \N__8699\,
            I => data_in_1_5
        );

    \I__802\ : LocalMux
    port map (
            O => \N__8696\,
            I => data_in_1_5
        );

    \I__801\ : InMux
    port map (
            O => \N__8687\,
            I => \N__8684\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__8684\,
            I => \c0.n28_adj_868\
        );

    \I__799\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8678\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__8678\,
            I => \c0.n26\
        );

    \I__797\ : CascadeMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__796\ : InMux
    port map (
            O => \N__8672\,
            I => \N__8666\
        );

    \I__795\ : InMux
    port map (
            O => \N__8671\,
            I => \N__8666\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__8666\,
            I => \c0.data_in_frame_7_3\
        );

    \I__793\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8660\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__8660\,
            I => \N__8657\
        );

    \I__791\ : Odrv4
    port map (
            O => \N__8657\,
            I => \c0.n4601\
        );

    \I__790\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8648\
        );

    \I__789\ : InMux
    port map (
            O => \N__8653\,
            I => \N__8648\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__8648\,
            I => \c0.data_in_frame_6_6\
        );

    \I__787\ : InMux
    port map (
            O => \N__8645\,
            I => \N__8642\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__8642\,
            I => \c0.n4592\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__8639\,
            I => \c0.n25_cascade_\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__8636\,
            I => \c0.n4591_cascade_\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__8633\,
            I => \c0.n28_cascade_\
        );

    \I__782\ : InMux
    port map (
            O => \N__8630\,
            I => \N__8627\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__8627\,
            I => \c0.n22\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__8624\,
            I => \c0.n4849_cascade_\
        );

    \I__779\ : InMux
    port map (
            O => \N__8621\,
            I => \N__8618\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__8618\,
            I => \c0.n4568\
        );

    \I__777\ : InMux
    port map (
            O => \N__8615\,
            I => \N__8612\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__8612\,
            I => \c0.n4582\
        );

    \I__775\ : InMux
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__8606\,
            I => n6
        );

    \I__773\ : InMux
    port map (
            O => \N__8603\,
            I => n3870
        );

    \I__772\ : InMux
    port map (
            O => \N__8600\,
            I => n3871
        );

    \I__771\ : InMux
    port map (
            O => \N__8597\,
            I => n3872
        );

    \I__770\ : InMux
    port map (
            O => \N__8594\,
            I => n3873
        );

    \I__769\ : InMux
    port map (
            O => \N__8591\,
            I => \bfn_1_25_0_\
        );

    \I__768\ : InMux
    port map (
            O => \N__8588\,
            I => n3875
        );

    \I__767\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8582\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__8582\,
            I => n14
        );

    \I__765\ : InMux
    port map (
            O => \N__8579\,
            I => n3862
        );

    \I__764\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8573\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__8573\,
            I => n13
        );

    \I__762\ : InMux
    port map (
            O => \N__8570\,
            I => n3863
        );

    \I__761\ : InMux
    port map (
            O => \N__8567\,
            I => \N__8564\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__8564\,
            I => n12
        );

    \I__759\ : InMux
    port map (
            O => \N__8561\,
            I => n3864
        );

    \I__758\ : InMux
    port map (
            O => \N__8558\,
            I => \N__8555\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__8555\,
            I => n11
        );

    \I__756\ : InMux
    port map (
            O => \N__8552\,
            I => n3865
        );

    \I__755\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8546\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__8546\,
            I => n10
        );

    \I__753\ : InMux
    port map (
            O => \N__8543\,
            I => \bfn_1_24_0_\
        );

    \I__752\ : InMux
    port map (
            O => \N__8540\,
            I => \N__8537\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__8537\,
            I => n9
        );

    \I__750\ : InMux
    port map (
            O => \N__8534\,
            I => n3867
        );

    \I__749\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8528\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__8528\,
            I => n8
        );

    \I__747\ : InMux
    port map (
            O => \N__8525\,
            I => n3868
        );

    \I__746\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8519\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__8519\,
            I => n7
        );

    \I__744\ : InMux
    port map (
            O => \N__8516\,
            I => n3869
        );

    \I__743\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8510\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__8510\,
            I => n22
        );

    \I__741\ : InMux
    port map (
            O => \N__8507\,
            I => n3854
        );

    \I__740\ : InMux
    port map (
            O => \N__8504\,
            I => \N__8501\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__8501\,
            I => n21
        );

    \I__738\ : InMux
    port map (
            O => \N__8498\,
            I => n3855
        );

    \I__737\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8492\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__8492\,
            I => n20
        );

    \I__735\ : InMux
    port map (
            O => \N__8489\,
            I => n3856
        );

    \I__734\ : InMux
    port map (
            O => \N__8486\,
            I => \N__8483\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__8483\,
            I => n19
        );

    \I__732\ : InMux
    port map (
            O => \N__8480\,
            I => n3857
        );

    \I__731\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8474\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__8474\,
            I => n18
        );

    \I__729\ : InMux
    port map (
            O => \N__8471\,
            I => \bfn_1_23_0_\
        );

    \I__728\ : InMux
    port map (
            O => \N__8468\,
            I => \N__8465\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__8465\,
            I => n17
        );

    \I__726\ : InMux
    port map (
            O => \N__8462\,
            I => n3859
        );

    \I__725\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8456\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__8456\,
            I => n16
        );

    \I__723\ : InMux
    port map (
            O => \N__8453\,
            I => n3860
        );

    \I__722\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8447\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__8447\,
            I => n15
        );

    \I__720\ : InMux
    port map (
            O => \N__8444\,
            I => n3861
        );

    \I__719\ : IoInMux
    port map (
            O => \N__8441\,
            I => \N__8438\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__8438\,
            I => \N__8435\
        );

    \I__717\ : IoSpan4Mux
    port map (
            O => \N__8435\,
            I => \N__8432\
        );

    \I__716\ : IoSpan4Mux
    port map (
            O => \N__8432\,
            I => \N__8429\
        );

    \I__715\ : IoSpan4Mux
    port map (
            O => \N__8429\,
            I => \N__8426\
        );

    \I__714\ : Odrv4
    port map (
            O => \N__8426\,
            I => \CLK_pad_gb_input\
        );

    \I__713\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8420\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__8420\,
            I => n26
        );

    \I__711\ : InMux
    port map (
            O => \N__8417\,
            I => \bfn_1_22_0_\
        );

    \I__710\ : InMux
    port map (
            O => \N__8414\,
            I => \N__8411\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__8411\,
            I => n25
        );

    \I__708\ : InMux
    port map (
            O => \N__8408\,
            I => n3851
        );

    \I__707\ : InMux
    port map (
            O => \N__8405\,
            I => \N__8402\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__8402\,
            I => n24
        );

    \I__705\ : InMux
    port map (
            O => \N__8399\,
            I => n3852
        );

    \I__704\ : InMux
    port map (
            O => \N__8396\,
            I => \N__8393\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__8393\,
            I => n23
        );

    \I__702\ : InMux
    port map (
            O => \N__8390\,
            I => n3853
        );

    \IN_MUX_bfv_4_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_21_0_\
        );

    \IN_MUX_bfv_4_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx2.n3898\,
            carryinitout => \bfn_4_22_0_\
        );

    \IN_MUX_bfv_14_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_27_0_\
        );

    \IN_MUX_bfv_14_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx.n3883\,
            carryinitout => \bfn_14_28_0_\
        );

    \IN_MUX_bfv_5_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_32_0_\
        );

    \IN_MUX_bfv_9_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_25_0_\
        );

    \IN_MUX_bfv_6_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_25_0_\
        );

    \IN_MUX_bfv_6_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n3913\,
            carryinitout => \bfn_6_26_0_\
        );

    \IN_MUX_bfv_5_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_24_0_\
        );

    \IN_MUX_bfv_11_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_27_0_\
        );

    \IN_MUX_bfv_1_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_22_0_\
        );

    \IN_MUX_bfv_1_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n3858,
            carryinitout => \bfn_1_23_0_\
        );

    \IN_MUX_bfv_1_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n3866,
            carryinitout => \bfn_1_24_0_\
        );

    \IN_MUX_bfv_1_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n3874,
            carryinitout => \bfn_1_25_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8441\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \blink_counter_323__i0_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8423\,
            in2 => \_gnd_net_\,
            in3 => \N__8417\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_1_22_0_\,
            carryout => n3851,
            clk => \N__22866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i1_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8414\,
            in2 => \_gnd_net_\,
            in3 => \N__8408\,
            lcout => n25,
            ltout => OPEN,
            carryin => n3851,
            carryout => n3852,
            clk => \N__22866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i2_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8405\,
            in2 => \_gnd_net_\,
            in3 => \N__8399\,
            lcout => n24,
            ltout => OPEN,
            carryin => n3852,
            carryout => n3853,
            clk => \N__22866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i3_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8396\,
            in2 => \_gnd_net_\,
            in3 => \N__8390\,
            lcout => n23,
            ltout => OPEN,
            carryin => n3853,
            carryout => n3854,
            clk => \N__22866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i4_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8513\,
            in2 => \_gnd_net_\,
            in3 => \N__8507\,
            lcout => n22,
            ltout => OPEN,
            carryin => n3854,
            carryout => n3855,
            clk => \N__22866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i5_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8504\,
            in2 => \_gnd_net_\,
            in3 => \N__8498\,
            lcout => n21,
            ltout => OPEN,
            carryin => n3855,
            carryout => n3856,
            clk => \N__22866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i6_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8495\,
            in2 => \_gnd_net_\,
            in3 => \N__8489\,
            lcout => n20,
            ltout => OPEN,
            carryin => n3856,
            carryout => n3857,
            clk => \N__22866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i7_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8486\,
            in2 => \_gnd_net_\,
            in3 => \N__8480\,
            lcout => n19,
            ltout => OPEN,
            carryin => n3857,
            carryout => n3858,
            clk => \N__22866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i8_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8477\,
            in2 => \_gnd_net_\,
            in3 => \N__8471\,
            lcout => n18,
            ltout => OPEN,
            carryin => \bfn_1_23_0_\,
            carryout => n3859,
            clk => \N__22867\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i9_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8468\,
            in2 => \_gnd_net_\,
            in3 => \N__8462\,
            lcout => n17,
            ltout => OPEN,
            carryin => n3859,
            carryout => n3860,
            clk => \N__22867\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i10_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8459\,
            in2 => \_gnd_net_\,
            in3 => \N__8453\,
            lcout => n16,
            ltout => OPEN,
            carryin => n3860,
            carryout => n3861,
            clk => \N__22867\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i11_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8450\,
            in2 => \_gnd_net_\,
            in3 => \N__8444\,
            lcout => n15,
            ltout => OPEN,
            carryin => n3861,
            carryout => n3862,
            clk => \N__22867\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i12_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8585\,
            in2 => \_gnd_net_\,
            in3 => \N__8579\,
            lcout => n14,
            ltout => OPEN,
            carryin => n3862,
            carryout => n3863,
            clk => \N__22867\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i13_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8576\,
            in2 => \_gnd_net_\,
            in3 => \N__8570\,
            lcout => n13,
            ltout => OPEN,
            carryin => n3863,
            carryout => n3864,
            clk => \N__22867\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i14_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8567\,
            in2 => \_gnd_net_\,
            in3 => \N__8561\,
            lcout => n12,
            ltout => OPEN,
            carryin => n3864,
            carryout => n3865,
            clk => \N__22867\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i15_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8558\,
            in2 => \_gnd_net_\,
            in3 => \N__8552\,
            lcout => n11,
            ltout => OPEN,
            carryin => n3865,
            carryout => n3866,
            clk => \N__22867\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i16_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8549\,
            in2 => \_gnd_net_\,
            in3 => \N__8543\,
            lcout => n10,
            ltout => OPEN,
            carryin => \bfn_1_24_0_\,
            carryout => n3867,
            clk => \N__22868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i17_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8540\,
            in2 => \_gnd_net_\,
            in3 => \N__8534\,
            lcout => n9,
            ltout => OPEN,
            carryin => n3867,
            carryout => n3868,
            clk => \N__22868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i18_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8531\,
            in2 => \_gnd_net_\,
            in3 => \N__8525\,
            lcout => n8,
            ltout => OPEN,
            carryin => n3868,
            carryout => n3869,
            clk => \N__22868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i19_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8522\,
            in2 => \_gnd_net_\,
            in3 => \N__8516\,
            lcout => n7,
            ltout => OPEN,
            carryin => n3869,
            carryout => n3870,
            clk => \N__22868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i20_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8609\,
            in2 => \_gnd_net_\,
            in3 => \N__8603\,
            lcout => n6,
            ltout => OPEN,
            carryin => n3870,
            carryout => n3871,
            clk => \N__22868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i21_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11080\,
            in2 => \_gnd_net_\,
            in3 => \N__8600\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n3871,
            carryout => n3872,
            clk => \N__22868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i22_LC_1_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11125\,
            in2 => \_gnd_net_\,
            in3 => \N__8597\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n3872,
            carryout => n3873,
            clk => \N__22868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i23_LC_1_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11056\,
            in2 => \_gnd_net_\,
            in3 => \N__8594\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n3873,
            carryout => n3874,
            clk => \N__22868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i24_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11104\,
            in2 => \_gnd_net_\,
            in3 => \N__8591\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_1_25_0_\,
            carryout => n3875,
            clk => \N__22871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_323__i25_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12229\,
            in2 => \_gnd_net_\,
            in3 => \N__8588\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i55_LC_1_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__8822\,
            in1 => \N__15028\,
            in2 => \N__14589\,
            in3 => \N__13685\,
            lcout => \c0.data_in_frame_6_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i39_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17090\,
            in1 => \N__9055\,
            in2 => \_gnd_net_\,
            in3 => \N__11715\,
            lcout => data_in_4_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i31_LC_1_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11716\,
            in1 => \N__17091\,
            in2 => \_gnd_net_\,
            in3 => \N__11834\,
            lcout => data_in_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_1__bdd_4_lut_4483_LC_1_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__8810\,
            in1 => \N__15638\,
            in2 => \N__15783\,
            in3 => \N__8615\,
            lcout => OPEN,
            ltout => \c0.n4849_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4849_bdd_4_lut_LC_1_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__15761\,
            in1 => \N__9713\,
            in2 => \N__8624\,
            in3 => \N__8621\,
            lcout => tx2_data_7_keep,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4213_3_lut_LC_1_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15517\,
            in1 => \N__9929\,
            in2 => \_gnd_net_\,
            in3 => \N__13376\,
            lcout => \c0.n4568\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4216_3_lut_LC_1_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15516\,
            in1 => \N__13763\,
            in2 => \_gnd_net_\,
            in3 => \N__10175\,
            lcout => \c0.n4571\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i6_LC_1_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8977\,
            in1 => \N__8714\,
            in2 => \_gnd_net_\,
            in3 => \N__17002\,
            lcout => data_in_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i40_LC_1_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17001\,
            in1 => \N__11514\,
            in2 => \_gnd_net_\,
            in3 => \N__11498\,
            lcout => data_in_4_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i27_LC_1_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17000\,
            in1 => \N__11384\,
            in2 => \_gnd_net_\,
            in3 => \N__9801\,
            lcout => data_in_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4227_3_lut_LC_1_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15560\,
            in1 => \N__12046\,
            in2 => \_gnd_net_\,
            in3 => \N__12876\,
            lcout => \c0.n4582\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i19_LC_1_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16999\,
            in1 => \N__9800\,
            in2 => \_gnd_net_\,
            in3 => \N__10085\,
            lcout => data_in_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i58_LC_1_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__8839\,
            in1 => \N__15882\,
            in2 => \N__14715\,
            in3 => \N__14962\,
            lcout => \c0.data_in_frame_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i1_LC_1_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17126\,
            in1 => \N__9180\,
            in2 => \_gnd_net_\,
            in3 => \N__8956\,
            lcout => data_in_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_1__bdd_4_lut_4454_LC_1_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__15646\,
            in1 => \N__8663\,
            in2 => \N__15788\,
            in3 => \N__9002\,
            lcout => \c0.n4813\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i13_LC_1_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__8712\,
            in1 => \N__14961\,
            in2 => \N__14721\,
            in3 => \N__13146\,
            lcout => \c0.data_in_field_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4236_3_lut_LC_1_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15559\,
            in1 => \N__12008\,
            in2 => \_gnd_net_\,
            in3 => \N__10021\,
            lcout => OPEN,
            ltout => \c0.n4591_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_1__bdd_4_lut_4478_LC_1_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__15778\,
            in1 => \N__15647\,
            in2 => \N__8636\,
            in3 => \N__8645\,
            lcout => \c0.n4831\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_LC_1_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8973\,
            in2 => \_gnd_net_\,
            in3 => \N__15078\,
            lcout => \c0.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4197_3_lut_LC_1_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15558\,
            in1 => \N__9979\,
            in2 => \_gnd_net_\,
            in3 => \N__13145\,
            lcout => \c0.n4552\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13784\,
            in1 => \N__9128\,
            in2 => \N__12143\,
            in3 => \N__9272\,
            lcout => OPEN,
            ltout => \c0.n28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_LC_1_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10499\,
            in1 => \N__11838\,
            in2 => \N__8633\,
            in3 => \N__8630\,
            lcout => \c0.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i14_LC_1_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8713\,
            in1 => \N__9772\,
            in2 => \_gnd_net_\,
            in3 => \N__17120\,
            lcout => data_in_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22888\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i11_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17116\,
            in1 => \N__15071\,
            in2 => \_gnd_net_\,
            in3 => \N__10087\,
            lcout => data_in_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22888\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i54_LC_1_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__8654\,
            in1 => \N__14946\,
            in2 => \N__14725\,
            in3 => \N__13939\,
            lcout => \c0.data_in_frame_6_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22888\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i23_LC_1_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__9273\,
            in1 => \_gnd_net_\,
            in2 => \N__17127\,
            in3 => \N__11839\,
            lcout => data_in_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22888\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i41_LC_1_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__14707\,
            in1 => \N__14945\,
            in2 => \N__17468\,
            in3 => \N__13895\,
            lcout => \c0.data_in_field_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22888\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4237_3_lut_LC_1_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__8758\,
            in1 => \N__8653\,
            in2 => \N__15546\,
            in3 => \_gnd_net_\,
            lcout => \c0.n4592\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9082\,
            in1 => \N__10086\,
            in2 => \N__9366\,
            in3 => \N__8945\,
            lcout => OPEN,
            ltout => \c0.n25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8687\,
            in1 => \N__8681\,
            in2 => \N__8639\,
            in3 => \N__9383\,
            lcout => \c0.n3933\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i9_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8952\,
            in1 => \N__16923\,
            in2 => \_gnd_net_\,
            in3 => \N__9410\,
            lcout => data_in_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i30_LC_1_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16920\,
            in1 => \N__10636\,
            in2 => \_gnd_net_\,
            in3 => \N__9129\,
            lcout => data_in_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i18_LC_1_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10556\,
            in1 => \N__16922\,
            in2 => \_gnd_net_\,
            in3 => \N__10503\,
            lcout => data_in_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i13_LC_1_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16919\,
            in1 => \N__12112\,
            in2 => \_gnd_net_\,
            in3 => \N__9359\,
            lcout => data_in_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_291_LC_1_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9332\,
            in1 => \N__9099\,
            in2 => \N__9697\,
            in3 => \N__8708\,
            lcout => \c0.n28_adj_868\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i7_LC_1_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__16921\,
            in1 => \_gnd_net_\,
            in2 => \N__9226\,
            in3 => \N__9103\,
            lcout => data_in_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_LC_1_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10374\,
            in1 => \N__9827\,
            in2 => \N__9771\,
            in3 => \N__9404\,
            lcout => \c0.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i59_LC_1_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__14937\,
            in1 => \N__14716\,
            in2 => \N__8675\,
            in3 => \N__14118\,
            lcout => \c0.data_in_frame_7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22899\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4225_3_lut_LC_1_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__15547\,
            in1 => \_gnd_net_\,
            in2 => \N__9305\,
            in3 => \N__9142\,
            lcout => \c0.n4580\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i63_LC_1_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17020\,
            in1 => \N__12338\,
            in2 => \_gnd_net_\,
            in3 => \N__14084\,
            lcout => data_in_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22899\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i22_LC_1_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9764\,
            in1 => \N__17021\,
            in2 => \_gnd_net_\,
            in3 => \N__9130\,
            lcout => data_in_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22899\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4246_3_lut_LC_1_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8671\,
            in1 => \N__8767\,
            in2 => \_gnd_net_\,
            in3 => \N__15548\,
            lcout => \c0.n4601\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i51_LC_1_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__8768\,
            in1 => \N__14939\,
            in2 => \N__14726\,
            in3 => \N__16595\,
            lcout => \c0.data_in_frame_6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22899\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i62_LC_1_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__14938\,
            in1 => \N__14085\,
            in2 => \N__8759\,
            in3 => \N__14720\,
            lcout => \c0.data_in_frame_7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22899\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i52_LC_1_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__8857\,
            in1 => \N__11984\,
            in2 => \N__14714\,
            in3 => \N__15046\,
            lcout => \c0.data_in_frame_6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22907\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i12_LC_1_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9829\,
            in1 => \N__17094\,
            in2 => \_gnd_net_\,
            in3 => \N__9077\,
            lcout => data_in_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22907\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i20_LC_1_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17093\,
            in1 => \N__14209\,
            in2 => \_gnd_net_\,
            in3 => \N__9828\,
            lcout => data_in_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22907\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i4_LC_1_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17095\,
            in1 => \N__10375\,
            in2 => \_gnd_net_\,
            in3 => \N__9078\,
            lcout => data_in_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22907\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4168_3_lut_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8725\,
            in1 => \N__9427\,
            in2 => \_gnd_net_\,
            in3 => \N__9506\,
            lcout => n4523,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_388_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12569\,
            in2 => \_gnd_net_\,
            in3 => \N__12640\,
            lcout => n11_adj_941,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4831_bdd_4_lut_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001010"
        )
    port map (
            in0 => \N__8774\,
            in1 => \N__9728\,
            in2 => \N__15787\,
            in3 => \N__8741\,
            lcout => OPEN,
            ltout => \tx2_data_6_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i6_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11228\,
            in2 => \N__8729\,
            in3 => \N__8726\,
            lcout => \r_Tx_Data_6_adj_958\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4243_3_lut_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8785\,
            in1 => \N__8864\,
            in2 => \_gnd_net_\,
            in3 => \N__15518\,
            lcout => \c0.n4598\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4249_3_lut_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8843\,
            in1 => \N__12932\,
            in2 => \_gnd_net_\,
            in3 => \N__15467\,
            lcout => OPEN,
            ltout => \c0.n4604_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_1__bdd_4_lut_4449_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__15731\,
            in1 => \N__15635\,
            in2 => \N__8825\,
            in3 => \N__9644\,
            lcout => \c0.n4807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4228_3_lut_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8797\,
            in1 => \N__15466\,
            in2 => \_gnd_net_\,
            in3 => \N__8821\,
            lcout => \c0.n4583\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i63_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__14963\,
            in1 => \N__14574\,
            in2 => \N__8801\,
            in3 => \N__13723\,
            lcout => \c0.data_in_frame_7_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22872\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i60_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__8786\,
            in1 => \N__13835\,
            in2 => \N__14670\,
            in3 => \N__14964\,
            lcout => \c0.data_in_frame_7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22872\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4200_3_lut_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15471\,
            in1 => \N__12790\,
            in2 => \_gnd_net_\,
            in3 => \N__9896\,
            lcout => \c0.n4555\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1384_2_lut_4_lut_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__9550\,
            in1 => \N__9575\,
            in2 => \N__12572\,
            in3 => \N__9505\,
            lcout => n1611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Bit_Index_1__bdd_4_lut_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__9574\,
            in1 => \N__8882\,
            in2 => \N__9549\,
            in3 => \N__8912\,
            lcout => n4777,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i5_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11247\,
            in1 => \N__8984\,
            in2 => \_gnd_net_\,
            in3 => \N__8921\,
            lcout => \r_Tx_Data_5_adj_959\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i7_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8891\,
            in1 => \N__11248\,
            in2 => \_gnd_net_\,
            in3 => \N__8927\,
            lcout => \r_Tx_Data_7_adj_957\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4269_3_lut_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9490\,
            in1 => \N__8920\,
            in2 => \_gnd_net_\,
            in3 => \N__8899\,
            lcout => n4624,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_1__bdd_4_lut_4444_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__15639\,
            in1 => \N__8870\,
            in2 => \N__15784\,
            in3 => \N__11858\,
            lcout => OPEN,
            ltout => \c0.n4801_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4801_bdd_4_lut_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__8876\,
            in1 => \N__15765\,
            in2 => \N__8906\,
            in3 => \N__9674\,
            lcout => OPEN,
            ltout => \tx2_data_1_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i1_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__8900\,
            in1 => \_gnd_net_\,
            in2 => \N__8903\,
            in3 => \N__11246\,
            lcout => \r_Tx_Data_1_adj_963\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4270_3_lut_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9491\,
            in1 => \N__8890\,
            in2 => \_gnd_net_\,
            in3 => \N__9017\,
            lcout => n4625,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4185_3_lut_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15512\,
            in1 => \N__12836\,
            in2 => \_gnd_net_\,
            in3 => \N__13496\,
            lcout => \c0.n4540\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4251_3_lut_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15525\,
            in1 => \N__13906\,
            in2 => \_gnd_net_\,
            in3 => \N__10132\,
            lcout => \c0.n4606\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i22_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__9742\,
            in1 => \N__14646\,
            in2 => \N__9290\,
            in3 => \N__15033\,
            lcout => \c0.data_in_field_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4239_3_lut_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13044\,
            in1 => \N__15511\,
            in2 => \_gnd_net_\,
            in3 => \N__13328\,
            lcout => \c0.n4594\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4198_3_lut_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11693\,
            in1 => \N__15526\,
            in2 => \_gnd_net_\,
            in3 => \N__10240\,
            lcout => OPEN,
            ltout => \c0.n4553_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4825_bdd_4_lut_LC_2_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__15760\,
            in1 => \N__8996\,
            in2 => \N__8987\,
            in3 => \N__9032\,
            lcout => tx2_data_5_keep,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_321_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10174\,
            in1 => \N__9928\,
            in2 => \N__15883\,
            in3 => \N__10019\,
            lcout => \c0.n10_adj_876\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13597\,
            in1 => \N__9741\,
            in2 => \_gnd_net_\,
            in3 => \N__13327\,
            lcout => \c0.n1284\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i5_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__14958\,
            in1 => \N__14641\,
            in2 => \N__8978\,
            in3 => \N__9980\,
            lcout => \c0.data_in_field_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i59_LC_2_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17129\,
            in1 => \N__9254\,
            in2 => \_gnd_net_\,
            in3 => \N__15878\,
            lcout => data_in_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i8_LC_2_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__14959\,
            in1 => \N__14644\,
            in2 => \N__8957\,
            in3 => \N__11596\,
            lcout => \c0.data_in_field_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i47_LC_2_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17128\,
            in1 => \N__9054\,
            in2 => \_gnd_net_\,
            in3 => \N__13940\,
            lcout => data_in_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i46_LC_2_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__14957\,
            in1 => \N__9056\,
            in2 => \N__10025\,
            in3 => \N__14643\,
            lcout => \c0.data_in_field_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i36_LC_2_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__14645\,
            in1 => \N__14960\,
            in2 => \N__13612\,
            in3 => \N__11948\,
            lcout => \c0.data_in_field_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i37_LC_2_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__14956\,
            in1 => \N__10640\,
            in2 => \N__13342\,
            in3 => \N__14642\,
            lcout => \c0.data_in_field_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_1__bdd_4_lut_4464_LC_2_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__10190\,
            in1 => \N__15640\,
            in2 => \N__15782\,
            in3 => \N__9038\,
            lcout => \c0.n4825\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4813_bdd_4_lut_LC_2_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000100010"
        )
    port map (
            in0 => \N__9656\,
            in1 => \N__15766\,
            in2 => \N__10397\,
            in3 => \N__9026\,
            lcout => OPEN,
            ltout => \tx2_data_3_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i3_LC_2_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11252\,
            in2 => \N__9020\,
            in3 => \N__9016\,
            lcout => \r_Tx_Data_3_adj_961\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22889\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i20_LC_2_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__15021\,
            in1 => \N__12113\,
            in2 => \N__11182\,
            in3 => \N__14628\,
            lcout => \c0.data_in_field_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22889\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i35_LC_2_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__13644\,
            in1 => \N__14234\,
            in2 => \N__14702\,
            in3 => \N__15024\,
            lcout => \c0.data_in_field_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22889\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4245_3_lut_LC_2_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15520\,
            in1 => \N__13558\,
            in2 => \_gnd_net_\,
            in3 => \N__13643\,
            lcout => \c0.n4600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i6_LC_2_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__9107\,
            in1 => \N__15023\,
            in2 => \N__14703\,
            in3 => \N__9894\,
            lcout => \c0.data_in_field_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22889\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_296_LC_2_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13886\,
            in2 => \_gnd_net_\,
            in3 => \N__11338\,
            lcout => \c0.n4450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i45_LC_2_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__14621\,
            in1 => \N__15022\,
            in2 => \N__10664\,
            in3 => \N__13031\,
            lcout => \c0.data_in_field_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22889\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_323_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14086\,
            in2 => \_gnd_net_\,
            in3 => \N__10988\,
            lcout => \c0.n6_adj_877\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i33_LC_2_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__14629\,
            in1 => \N__14932\,
            in2 => \N__10133\,
            in3 => \N__10577\,
            lcout => \c0.data_in_field_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22894\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_rep_38_2_lut_LC_2_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10989\,
            in2 => \_gnd_net_\,
            in3 => \N__9920\,
            lcout => \c0.n4927\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i31_LC_2_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__9921\,
            in1 => \N__10607\,
            in2 => \N__14706\,
            in3 => \N__14933\,
            lcout => \c0.data_in_field_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22894\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i11_LC_2_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__14928\,
            in1 => \N__9083\,
            in2 => \N__11355\,
            in3 => \N__14639\,
            lcout => \c0.data_in_field_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22894\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i0_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__9181\,
            in1 => \N__14930\,
            in2 => \N__14704\,
            in3 => \N__11631\,
            lcout => \c0.data_in_field_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22894\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i27_LC_2_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__14929\,
            in1 => \N__14210\,
            in2 => \N__10424\,
            in3 => \N__14640\,
            lcout => \c0.data_in_field_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22894\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i12_LC_2_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__9368\,
            in1 => \N__14931\,
            in2 => \N__14705\,
            in3 => \N__14012\,
            lcout => \c0.data_in_field_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22894\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_293_LC_2_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12105\,
            in1 => \N__14202\,
            in2 => \N__9188\,
            in3 => \N__9808\,
            lcout => OPEN,
            ltout => \c0.n25_adj_870_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__9161\,
            in1 => \N__9197\,
            in2 => \N__9155\,
            in3 => \N__9152\,
            lcout => \c0.n1197\,
            ltout => \c0.n1197_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i48_LC_2_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__14687\,
            in1 => \N__9143\,
            in2 => \N__9146\,
            in3 => \N__16088\,
            lcout => \c0.data_in_frame_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22900\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i8_LC_2_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9336\,
            in1 => \N__9696\,
            in2 => \_gnd_net_\,
            in3 => \N__16918\,
            lcout => data_in_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22900\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i15_LC_2_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__14686\,
            in1 => \N__14940\,
            in2 => \N__9338\,
            in3 => \N__10450\,
            lcout => \c0.data_in_field_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22900\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i14_LC_2_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__9227\,
            in1 => \N__12786\,
            in2 => \N__15025\,
            in3 => \N__14688\,
            lcout => \c0.data_in_field_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22900\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i25_LC_2_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16917\,
            in1 => \N__14254\,
            in2 => \_gnd_net_\,
            in3 => \N__13785\,
            lcout => data_in_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22900\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i29_LC_2_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__9131\,
            in1 => \N__14944\,
            in2 => \N__10241\,
            in3 => \N__14689\,
            lcout => \c0.data_in_field_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22900\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i60_LC_2_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__10699\,
            in1 => \_gnd_net_\,
            in2 => \N__17098\,
            in3 => \N__14114\,
            lcout => data_in_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i56_LC_2_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__15019\,
            in1 => \N__9304\,
            in2 => \N__16132\,
            in3 => \N__14693\,
            lcout => \c0.data_in_frame_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i10_LC_2_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17064\,
            in1 => \N__10504\,
            in2 => \_gnd_net_\,
            in3 => \N__11806\,
            lcout => data_in_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i24_LC_2_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11439\,
            in1 => \N__17069\,
            in2 => \_gnd_net_\,
            in3 => \N__10602\,
            lcout => data_in_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i16_LC_2_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__9408\,
            in1 => \N__15020\,
            in2 => \N__14722\,
            in3 => \N__10163\,
            lcout => \c0.data_in_field_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i34_LC_2_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17019\,
            in1 => \N__10572\,
            in2 => \_gnd_net_\,
            in3 => \N__17458\,
            lcout => data_in_4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i15_LC_2_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17065\,
            in1 => \N__9219\,
            in2 => \_gnd_net_\,
            in3 => \N__9289\,
            lcout => data_in_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i2_LC_2_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__14150\,
            in1 => \N__15143\,
            in2 => \N__9250\,
            in3 => \N__17683\,
            lcout => rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_R_49_LC_2_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9233\,
            lcout => \c0.rx.r_Rx_Data_R\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_292_LC_2_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10598\,
            in1 => \N__9218\,
            in2 => \N__11917\,
            in3 => \N__10538\,
            lcout => \c0.n26_adj_869\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i17_LC_2_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17101\,
            in1 => \N__13792\,
            in2 => \_gnd_net_\,
            in3 => \N__9409\,
            lcout => data_in_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_LC_2_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11801\,
            in1 => \N__9942\,
            in2 => \N__11440\,
            in3 => \N__10680\,
            lcout => \c0.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_50_LC_2_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9374\,
            lcout => \r_Rx_Data\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i5_LC_2_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17100\,
            in1 => \N__9367\,
            in2 => \_gnd_net_\,
            in3 => \N__9943\,
            lcout => data_in_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i16_LC_2_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17099\,
            in2 => \N__9337\,
            in3 => \N__11435\,
            lcout => data_in_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i3_LC_2_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11913\,
            in1 => \N__17102\,
            in2 => \_gnd_net_\,
            in3 => \N__15079\,
            lcout => data_in_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_4_lut_4_lut_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__12410\,
            in1 => \N__10799\,
            in2 => \N__12649\,
            in3 => \N__10768\,
            lcout => n9_adj_939,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i5_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15223\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10733\,
            lcout => \c0.tx2.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i8_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15224\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10715\,
            lcout => \c0.tx2.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i1_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10514\,
            in2 => \_gnd_net_\,
            in3 => \N__15222\,
            lcout => \c0.tx2.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i4362_2_lut_3_lut_4_lut_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__12648\,
            in1 => \N__10802\,
            in2 => \N__12565\,
            in3 => \N__10769\,
            lcout => OPEN,
            ltout => \n4638_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Done_44_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111111000"
        )
    port map (
            in0 => \N__9449\,
            in1 => \N__9461\,
            in2 => \N__9452\,
            in3 => \N__12413\,
            lcout => tx2_done,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_1__bdd_4_lut_4459_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__9443\,
            in1 => \N__15636\,
            in2 => \N__15785\,
            in3 => \N__11189\,
            lcout => \c0.n4819\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_2_lut_3_lut_4_lut_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__12528\,
            in1 => \N__12644\,
            in2 => \N__12701\,
            in3 => \N__12411\,
            lcout => n1030,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4807_bdd_4_lut_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001010"
        )
    port map (
            in0 => \N__11141\,
            in1 => \N__9668\,
            in2 => \N__15786\,
            in3 => \N__9437\,
            lcout => OPEN,
            ltout => \tx2_data_2_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i2_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11227\,
            in2 => \N__9431\,
            in3 => \N__9428\,
            lcout => \r_Tx_Data_2_adj_962\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__12412\,
            in1 => \N__10748\,
            in2 => \N__12650\,
            in3 => \N__9416\,
            lcout => n6_adj_940,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i1_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001110010001000"
        )
    port map (
            in0 => \N__9614\,
            in1 => \N__9580\,
            in2 => \N__9551\,
            in3 => \N__9637\,
            lcout => \r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22877\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i4157_4_lut_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__12414\,
            in1 => \N__11403\,
            in2 => \N__12570\,
            in3 => \N__12600\,
            lcout => n4512,
            ltout => \n4512_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4159_2_lut_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9659\,
            in3 => \N__9633\,
            lcout => n4514,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4191_3_lut_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15470\,
            in1 => \N__11357\,
            in2 => \_gnd_net_\,
            in3 => \N__10313\,
            lcout => \c0.n4546\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4248_3_lut_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15519\,
            in1 => \N__13193\,
            in2 => \_gnd_net_\,
            in3 => \N__10343\,
            lcout => \c0.n4603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2099_4_lut_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001100000"
        )
    port map (
            in0 => \N__9579\,
            in1 => \N__9500\,
            in2 => \N__9638\,
            in3 => \N__9612\,
            lcout => OPEN,
            ltout => \n2326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i2_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__9501\,
            in1 => \N__9548\,
            in2 => \N__9623\,
            in3 => \N__9620\,
            lcout => \r_Bit_Index_2_adj_955\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22877\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i0_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000100010"
        )
    port map (
            in0 => \N__12558\,
            in1 => \N__9544\,
            in2 => \_gnd_net_\,
            in3 => \N__9613\,
            lcout => \r_Bit_Index_0_adj_956\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22877\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4167_3_lut_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11200\,
            in1 => \N__11011\,
            in2 => \_gnd_net_\,
            in3 => \N__9498\,
            lcout => OPEN,
            ltout => \n4522_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n4777_bdd_4_lut_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__9542\,
            in1 => \N__9602\,
            in2 => \N__9590\,
            in3 => \N__9587\,
            lcout => n4780,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_3_lut_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9581\,
            in1 => \N__9543\,
            in2 => \_gnd_net_\,
            in3 => \N__9499\,
            lcout => \c0.tx2.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_330_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13495\,
            in1 => \N__13759\,
            in2 => \N__12047\,
            in3 => \N__9866\,
            lcout => \c0.n8_adj_880\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4201_3_lut_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15521\,
            in1 => \N__13448\,
            in2 => \_gnd_net_\,
            in3 => \N__9743\,
            lcout => \c0.n4556\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_320_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10131\,
            in1 => \N__9895\,
            in2 => \N__13722\,
            in3 => \N__13598\,
            lcout => OPEN,
            ltout => \c0.n10_adj_874_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_322_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13645\,
            in1 => \N__10341\,
            in2 => \N__9716\,
            in3 => \N__9851\,
            lcout => \c0.n4469\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4212_3_lut_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__15513\,
            in1 => \N__10454\,
            in2 => \N__11663\,
            in3 => \_gnd_net_\,
            lcout => \c0.n4567\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i7_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__9704\,
            in1 => \N__11661\,
            in2 => \N__14501\,
            in3 => \N__15027\,
            lcout => \c0.data_in_field_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_338_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11474\,
            in1 => \N__10173\,
            in2 => \N__13265\,
            in3 => \N__10309\,
            lcout => \c0.n15_adj_885\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4186_3_lut_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10478\,
            in1 => \N__13297\,
            in2 => \_gnd_net_\,
            in3 => \N__15515\,
            lcout => \c0.n4541\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4189_3_lut_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15514\,
            in1 => \N__13530\,
            in2 => \_gnd_net_\,
            in3 => \N__10061\,
            lcout => \c0.n4544\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_303_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__11654\,
            in1 => \N__9887\,
            in2 => \_gnd_net_\,
            in3 => \N__9865\,
            lcout => \c0.n4408\,
            ltout => \c0.n4408_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_LC_3_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11592\,
            in1 => \N__10018\,
            in2 => \N__9854\,
            in3 => \N__9850\,
            lcout => \c0.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_337_LC_3_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11636\,
            in1 => \N__13151\,
            in2 => \N__16133\,
            in3 => \N__11771\,
            lcout => \c0.n16_adj_884\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_302_LC_3_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9977\,
            in1 => \N__10266\,
            in2 => \N__12878\,
            in3 => \N__11684\,
            lcout => \c0.n4468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i19_LC_3_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__9839\,
            in1 => \N__15042\,
            in2 => \N__10277\,
            in3 => \N__14653\,
            lcout => \c0.data_in_field_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22890\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i26_LC_3_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__14652\,
            in1 => \N__15038\,
            in2 => \N__9809\,
            in3 => \N__13531\,
            lcout => \c0.data_in_field_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22890\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i21_LC_3_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__9776\,
            in1 => \N__11685\,
            in2 => \N__15047\,
            in3 => \N__14654\,
            lcout => \c0.data_in_field_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22890\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_308_LC_3_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13636\,
            in1 => \N__10330\,
            in2 => \_gnd_net_\,
            in3 => \N__11172\,
            lcout => \c0.n1271\,
            ltout => \c0.n1271_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_357_LC_3_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11756\,
            in1 => \N__10120\,
            in2 => \N__9746\,
            in3 => \N__10060\,
            lcout => \c0.n4429\,
            ltout => \c0.n4429_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_341_LC_3_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13022\,
            in1 => \N__10211\,
            in2 => \N__10034\,
            in3 => \N__12895\,
            lcout => \c0.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_339_LC_3_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10031\,
            in1 => \N__10020\,
            in2 => \N__9992\,
            in3 => \N__9978\,
            lcout => \c0.n4430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i25_LC_3_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__10552\,
            in1 => \N__14997\,
            in2 => \N__14713\,
            in3 => \N__13284\,
            lcout => \c0.data_in_field_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_297_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14005\,
            in1 => \N__13283\,
            in2 => \N__10422\,
            in3 => \N__9956\,
            lcout => \c0.n1296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i34_LC_3_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__10331\,
            in1 => \N__11383\,
            in2 => \N__15043\,
            in3 => \N__14665\,
            lcout => \c0.data_in_field_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i4_LC_3_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__9950\,
            in1 => \N__14935\,
            in2 => \N__14712\,
            in3 => \N__11761\,
            lcout => \c0.data_in_field_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22901\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_310_LC_3_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__10987\,
            in1 => \N__9919\,
            in2 => \_gnd_net_\,
            in3 => \N__10470\,
            lcout => \c0.n1261\,
            ltout => \c0.n1261_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_312_LC_3_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13553\,
            in1 => \N__10445\,
            in2 => \N__9899\,
            in3 => \N__11892\,
            lcout => \c0.n4390\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i53_LC_3_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__14934\,
            in1 => \N__14655\,
            in2 => \N__10202\,
            in3 => \N__12284\,
            lcout => \c0.data_in_frame_6_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22901\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i43_LC_3_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__13554\,
            in1 => \N__16562\,
            in2 => \N__14711\,
            in3 => \N__14936\,
            lcout => \c0.data_in_field_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22901\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_294_LC_3_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12817\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13432\,
            lcout => \c0.n4411\,
            ltout => \c0.n4411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_354_LC_3_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11624\,
            in1 => \N__10233\,
            in2 => \N__10205\,
            in3 => \N__12779\,
            lcout => \c0.n4399\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4240_3_lut_LC_3_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10198\,
            in1 => \N__15528\,
            in2 => \_gnd_net_\,
            in3 => \N__10357\,
            lcout => \c0.n4595\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_298_LC_3_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__10119\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11757\,
            lcout => OPEN,
            ltout => \c0.n1340_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_324_LC_3_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13045\,
            in1 => \N__10250\,
            in2 => \N__10178\,
            in3 => \N__13068\,
            lcout => \c0.n4445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_306_LC_3_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10154\,
            in1 => \N__10295\,
            in2 => \N__10130\,
            in3 => \N__10052\,
            lcout => \c0.n8_adj_872\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i1_LC_3_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__15009\,
            in1 => \N__14694\,
            in2 => \N__12834\,
            in3 => \N__10685\,
            lcout => \c0.data_in_field_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22909\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i18_LC_3_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__10091\,
            in1 => \N__15012\,
            in2 => \N__14724\,
            in3 => \N__10053\,
            lcout => \c0.data_in_field_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22909\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i32_LC_3_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__15010\,
            in1 => \N__14255\,
            in2 => \N__10999\,
            in3 => \N__14695\,
            lcout => \c0.data_in_field_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22909\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i17_LC_3_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__10505\,
            in1 => \N__15011\,
            in2 => \N__14723\,
            in3 => \N__10474\,
            lcout => \c0.data_in_field_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22909\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_317_LC_3_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11339\,
            in1 => \N__10446\,
            in2 => \N__14014\,
            in3 => \N__11272\,
            lcout => \c0.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4192_3_lut_LC_3_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15545\,
            in1 => \N__10423\,
            in2 => \_gnd_net_\,
            in3 => \N__10276\,
            lcout => \c0.n4547\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i3_LC_3_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__10302\,
            in1 => \N__10382\,
            in2 => \N__14669\,
            in3 => \N__14978\,
            lcout => \c0.data_in_field_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22916\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i61_LC_3_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__14977\,
            in1 => \N__14570\,
            in2 => \N__12311\,
            in3 => \N__10358\,
            lcout => \c0.data_in_frame_7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22916\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_314_LC_3_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10342\,
            in1 => \N__10301\,
            in2 => \N__12310\,
            in3 => \N__10275\,
            lcout => \c0.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i45_LC_3_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11983\,
            in1 => \N__17024\,
            in2 => \_gnd_net_\,
            in3 => \N__12180\,
            lcout => data_in_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22916\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_349_LC_3_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13433\,
            in1 => \N__10232\,
            in2 => \_gnd_net_\,
            in3 => \N__12818\,
            lcout => \c0.n1280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i3_LC_3_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__15142\,
            in1 => \N__15110\,
            in2 => \N__10700\,
            in3 => \N__17711\,
            lcout => rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22916\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i46_LC_3_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17058\,
            in1 => \N__10653\,
            in2 => \_gnd_net_\,
            in3 => \N__12273\,
            lcout => data_in_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22923\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i2_LC_3_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11805\,
            in1 => \N__17059\,
            in2 => \_gnd_net_\,
            in3 => \N__10684\,
            lcout => data_in_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22923\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i38_LC_3_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17057\,
            in1 => \N__10654\,
            in2 => \_gnd_net_\,
            in3 => \N__10621\,
            lcout => data_in_4_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22923\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_3_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101001110000"
        )
    port map (
            in0 => \N__17555\,
            in1 => \N__17378\,
            in2 => \N__17778\,
            in3 => \N__16046\,
            lcout => OPEN,
            ltout => \c0.rx.n4873_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.n4873_bdd_4_lut_4_lut_LC_3_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111000001"
        )
    port map (
            in0 => \N__17686\,
            in1 => \N__17556\,
            in2 => \N__10610\,
            in3 => \N__17816\,
            lcout => \c0.rx.n4876\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i32_LC_3_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10603\,
            in1 => \N__11531\,
            in2 => \_gnd_net_\,
            in3 => \N__17060\,
            lcout => data_in_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22923\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i26_LC_3_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17056\,
            in1 => \N__10573\,
            in2 => \_gnd_net_\,
            in3 => \N__10545\,
            lcout => data_in_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22923\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_2_lut_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__10946\,
            in1 => \N__10945\,
            in2 => \N__12455\,
            in3 => \N__10517\,
            lcout => n1768,
            ltout => OPEN,
            carryin => \bfn_4_21_0_\,
            carryout => \c0.tx2.n3891\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_3_lut_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__10897\,
            in1 => \N__10896\,
            in2 => \N__12459\,
            in3 => \N__10508\,
            lcout => n1710,
            ltout => OPEN,
            carryin => \c0.tx2.n3891\,
            carryout => \c0.tx2.n3892\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_4_lut_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__10934\,
            in1 => \N__10933\,
            in2 => \N__12456\,
            in3 => \N__10742\,
            lcout => n1707,
            ltout => OPEN,
            carryin => \c0.tx2.n3892\,
            carryout => \c0.tx2.n3893\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_5_lut_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__10877\,
            in1 => \N__10876\,
            in2 => \N__12460\,
            in3 => \N__10739\,
            lcout => n1704,
            ltout => OPEN,
            carryin => \c0.tx2.n3893\,
            carryout => \c0.tx2.n3894\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_6_lut_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__10850\,
            in1 => \N__10849\,
            in2 => \N__12457\,
            in3 => \N__10736\,
            lcout => n1701,
            ltout => OPEN,
            carryin => \c0.tx2.n3894\,
            carryout => \c0.tx2.n3895\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_7_lut_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__10916\,
            in1 => \N__10915\,
            in2 => \N__12461\,
            in3 => \N__10727\,
            lcout => n1698,
            ltout => OPEN,
            carryin => \c0.tx2.n3895\,
            carryout => \c0.tx2.n3896\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_8_lut_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__15194\,
            in1 => \N__15193\,
            in2 => \N__12458\,
            in3 => \N__10724\,
            lcout => n1695,
            ltout => OPEN,
            carryin => \c0.tx2.n3896\,
            carryout => \c0.tx2.n3897\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_9_lut_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__10823\,
            in1 => \N__10822\,
            in2 => \N__12462\,
            in3 => \N__10721\,
            lcout => n1692,
            ltout => OPEN,
            carryin => \c0.tx2.n3897\,
            carryout => \c0.tx2.n3898\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_10_lut_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__10800\,
            in1 => \N__10801\,
            in2 => \N__12448\,
            in3 => \N__10718\,
            lcout => n1689,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i3_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15227\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10709\,
            lcout => \c0.tx2.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i2_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10958\,
            in2 => \_gnd_net_\,
            in3 => \N__15226\,
            lcout => \c0.tx2.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i0_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__15225\,
            in1 => \N__10952\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx2.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_4_lut_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__10932\,
            in1 => \N__10914\,
            in2 => \N__10898\,
            in3 => \N__10875\,
            lcout => OPEN,
            ltout => \c0.tx2.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2675_4_lut_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__15192\,
            in1 => \N__10848\,
            in2 => \N__10859\,
            in3 => \N__10821\,
            lcout => \c0.tx2.n2902\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i4_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10856\,
            in2 => \_gnd_net_\,
            in3 => \N__15228\,
            lcout => \c0.tx2.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i7_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__15229\,
            in1 => \_gnd_net_\,
            in2 => \N__10832\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx2.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2677_2_lut_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10797\,
            in2 => \_gnd_net_\,
            in3 => \N__10766\,
            lcout => \r_SM_Main_2_N_759_1\,
            ltout => \r_SM_Main_2_N_759_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i2_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__12623\,
            in1 => \N__12524\,
            in2 => \N__10805\,
            in3 => \N__12409\,
            lcout => \r_SM_Main_2_adj_952\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22878\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_3_lut_4_lut_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__12407\,
            in1 => \N__10798\,
            in2 => \N__12553\,
            in3 => \N__10767\,
            lcout => n4_adj_965,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4188_3_lut_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15430\,
            in1 => \N__14315\,
            in2 => \_gnd_net_\,
            in3 => \N__11897\,
            lcout => \c0.n4543\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i1_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__12408\,
            in1 => \N__12624\,
            in2 => \N__12554\,
            in3 => \N__11411\,
            lcout => \r_SM_Main_1_adj_953\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22878\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4164_4_lut_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000000"
        )
    port map (
            in0 => \N__11113\,
            in1 => \N__11134\,
            in2 => \N__11069\,
            in3 => \N__11089\,
            lcout => n4519,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4165_4_lut_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111100000"
        )
    port map (
            in0 => \N__11135\,
            in1 => \N__11114\,
            in2 => \N__11093\,
            in3 => \N__11068\,
            lcout => n4520,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_1__bdd_4_lut_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__15604\,
            in1 => \N__11045\,
            in2 => \N__15777\,
            in3 => \N__10964\,
            lcout => OPEN,
            ltout => \c0.n4855_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4855_bdd_4_lut_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__11030\,
            in1 => \N__15747\,
            in2 => \N__11018\,
            in3 => \N__11576\,
            lcout => OPEN,
            ltout => \tx2_data_0_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i0_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11229\,
            in2 => \N__11015\,
            in3 => \N__11012\,
            lcout => \r_Tx_Data_0_adj_964\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4224_3_lut_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15469\,
            in1 => \N__13976\,
            in2 => \_gnd_net_\,
            in3 => \N__11000\,
            lcout => \c0.n4579\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4194_3_lut_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15432\,
            in1 => \N__14018\,
            in2 => \_gnd_net_\,
            in3 => \N__11765\,
            lcout => OPEN,
            ltout => \c0.n4549_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4819_bdd_4_lut_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010011000"
        )
    port map (
            in0 => \N__11261\,
            in1 => \N__15746\,
            in2 => \N__11255\,
            in3 => \N__11156\,
            lcout => OPEN,
            ltout => \tx2_data_4_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i4_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11230\,
            in2 => \N__11204\,
            in3 => \N__11201\,
            lcout => \r_Tx_Data_4_adj_960\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4242_3_lut_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15468\,
            in1 => \N__12164\,
            in2 => \_gnd_net_\,
            in3 => \N__13613\,
            lcout => \c0.n4597\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4397_2_lut_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14405\,
            in2 => \_gnd_net_\,
            in3 => \N__13091\,
            lcout => \c0.n1675\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i48_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17087\,
            in1 => \N__11487\,
            in2 => \_gnd_net_\,
            in3 => \N__13681\,
            lcout => data_in_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4195_3_lut_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15431\,
            in1 => \N__13223\,
            in2 => \_gnd_net_\,
            in3 => \N__11183\,
            lcout => \c0.n4550\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_wait_for_transmission_621_LC_4_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110001101"
        )
    port map (
            in0 => \N__14406\,
            in1 => \N__12710\,
            in2 => \N__13099\,
            in3 => \N__15332\,
            lcout => \c0.FRAME_MATCHER_wait_for_transmission\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i639_4_lut_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__11150\,
            in1 => \N__12559\,
            in2 => \N__12694\,
            in3 => \N__11412\,
            lcout => OPEN,
            ltout => \n865_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i0_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001110100"
        )
    port map (
            in0 => \N__11414\,
            in1 => \N__12619\,
            in2 => \N__11144\,
            in3 => \N__12463\,
            lcout => \r_SM_Main_0_adj_954\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i4383_3_lut_4_lut_4_lut_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001000000010"
        )
    port map (
            in0 => \N__12688\,
            in1 => \N__12560\,
            in2 => \N__12638\,
            in3 => \N__11413\,
            lcout => OPEN,
            ltout => \n4366_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Active_47_LC_4_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011100"
        )
    port map (
            in0 => \N__12561\,
            in1 => \N__12725\,
            in2 => \N__11387\,
            in3 => \N__12464\,
            lcout => tx2_active,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i64_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13712\,
            in1 => \N__12065\,
            in2 => \_gnd_net_\,
            in3 => \N__17089\,
            lcout => data_in_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22891\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i35_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17088\,
            in1 => \N__14173\,
            in2 => \_gnd_net_\,
            in3 => \N__11373\,
            lcout => data_in_4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22891\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_329_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13752\,
            in1 => \N__11356\,
            in2 => \N__13907\,
            in3 => \N__13526\,
            lcout => OPEN,
            ltout => \c0.n8_adj_879_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_3_lut_adj_331_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11979\,
            in2 => \N__11312\,
            in3 => \N__13263\,
            lcout => OPEN,
            ltout => \c0.n4451_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_336_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__15853\,
            in1 => \N__11702\,
            in2 => \N__11309\,
            in3 => \N__11306\,
            lcout => \c0.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_295_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13184\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13222\,
            lcout => OPEN,
            ltout => \c0.n1357_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_333_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011101111011"
        )
    port map (
            in0 => \N__11297\,
            in1 => \N__11288\,
            in2 => \N__11282\,
            in3 => \N__11279\,
            lcout => \c0.n22_adj_881\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_346_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011101111011"
        )
    port map (
            in0 => \N__11564\,
            in1 => \N__11558\,
            in2 => \N__11552\,
            in3 => \N__11543\,
            lcout => OPEN,
            ltout => \c0.n17_adj_889_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_352_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111101"
        )
    port map (
            in0 => \N__13382\,
            in1 => \N__11453\,
            in2 => \N__11537\,
            in3 => \N__12752\,
            lcout => \c0.n25_adj_893\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_300_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13972\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12037\,
            lcout => OPEN,
            ltout => \c0.n4387_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_325_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13185\,
            in1 => \N__12283\,
            in2 => \N__11534\,
            in3 => \N__11470\,
            lcout => \c0.n4388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i39_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__14464\,
            in1 => \N__15035\,
            in2 => \N__11530\,
            in3 => \N__12038\,
            lcout => \c0.data_in_field_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i47_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__15034\,
            in1 => \N__14465\,
            in2 => \N__12877\,
            in3 => \N__11497\,
            lcout => \c0.data_in_field_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_345_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13076\,
            in1 => \N__13264\,
            in2 => \N__17276\,
            in3 => \N__11469\,
            lcout => \c0.n11_adj_888\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i23_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__13367\,
            in1 => \N__15031\,
            in2 => \N__11447\,
            in3 => \N__14472\,
            lcout => \c0.data_in_field_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22902\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i28_LC_4_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__15029\,
            in1 => \N__12139\,
            in2 => \N__14578\,
            in3 => \N__13221\,
            lcout => \c0.data_in_field_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22902\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i9_LC_4_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__13481\,
            in1 => \N__15032\,
            in2 => \N__11813\,
            in3 => \N__14473\,
            lcout => \c0.data_in_field_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22902\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_304_LC_4_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13525\,
            in2 => \_gnd_net_\,
            in3 => \N__13366\,
            lcout => OPEN,
            ltout => \c0.n8_adj_871_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_LC_4_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13480\,
            in1 => \N__13742\,
            in2 => \N__11780\,
            in3 => \N__11777\,
            lcout => \c0.n1418\,
            ltout => \c0.n1418_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_309_LC_4_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11755\,
            in1 => \N__15943\,
            in2 => \N__11729\,
            in3 => \N__13393\,
            lcout => \c0.n4474\,
            ltout => \c0.n4474_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_LC_4_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13673\,
            in2 => \N__11726\,
            in3 => \N__13183\,
            lcout => \c0.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i38_LC_4_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__15030\,
            in1 => \N__11723\,
            in2 => \N__14579\,
            in3 => \N__12007\,
            lcout => \c0.data_in_field_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22902\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_299_LC_4_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12003\,
            in2 => \_gnd_net_\,
            in3 => \N__11602\,
            lcout => \c0.n4396\,
            ltout => \c0.n4396_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_316_LC_4_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16751\,
            in1 => \N__11692\,
            in2 => \N__11666\,
            in3 => \N__11662\,
            lcout => \c0.n12_adj_873\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4215_3_lut_LC_4_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15510\,
            in1 => \N__11635\,
            in2 => \_gnd_net_\,
            in3 => \N__11603\,
            lcout => \c0.n4570\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i29_LC_4_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11943\,
            in1 => \N__17062\,
            in2 => \_gnd_net_\,
            in3 => \N__12137\,
            lcout => data_in_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_353_LC_4_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12042\,
            in1 => \N__12002\,
            in2 => \N__14311\,
            in3 => \N__13963\,
            lcout => \c0.n1290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i53_LC_4_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11978\,
            in1 => \N__13821\,
            in2 => \_gnd_net_\,
            in3 => \N__17063\,
            lcout => data_in_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i37_LC_4_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17061\,
            in1 => \N__12191\,
            in2 => \_gnd_net_\,
            in3 => \N__11944\,
            lcout => data_in_4_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_3_lut_LC_4_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__11891\,
            in1 => \N__12159\,
            in2 => \_gnd_net_\,
            in3 => \N__11927\,
            lcout => \c0.n1267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i2_LC_4_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__11921\,
            in1 => \N__15016\,
            in2 => \N__14590\,
            in3 => \N__11896\,
            lcout => \c0.data_in_field_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i57_LC_4_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__15015\,
            in1 => \N__14486\,
            in2 => \N__11870\,
            in3 => \N__17272\,
            lcout => \c0.data_in_frame_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4252_3_lut_LC_4_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15544\,
            in1 => \N__11866\,
            in2 => \_gnd_net_\,
            in3 => \N__12202\,
            lcout => \c0.n4607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i30_LC_4_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__15013\,
            in1 => \N__11843\,
            in2 => \N__13447\,
            in3 => \N__14493\,
            lcout => \c0.data_in_field_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i49_LC_4_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__12203\,
            in1 => \N__16762\,
            in2 => \N__14591\,
            in3 => \N__15018\,
            lcout => \c0.data_in_frame_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i44_LC_4_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__15014\,
            in1 => \N__14485\,
            in2 => \N__12190\,
            in3 => \N__12163\,
            lcout => \c0.data_in_field_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i40_LC_4_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__14484\,
            in1 => \N__15017\,
            in2 => \N__14276\,
            in3 => \N__13971\,
            lcout => \c0.data_in_field_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i21_LC_4_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12138\,
            in1 => \N__16996\,
            in2 => \_gnd_net_\,
            in3 => \N__12104\,
            lcout => data_in_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i4_LC_4_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__15127\,
            in1 => \N__14142\,
            in2 => \N__13852\,
            in3 => \N__17707\,
            lcout => rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22924\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i5_LC_4_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__17705\,
            in1 => \N__15128\,
            in2 => \N__12077\,
            in3 => \N__15105\,
            lcout => rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22924\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i62_LC_4_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17023\,
            in1 => \N__12073\,
            in2 => \_gnd_net_\,
            in3 => \N__12308\,
            lcout => data_in_7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22924\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i57_LC_4_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17022\,
            in1 => \N__15155\,
            in2 => \_gnd_net_\,
            in3 => \N__16118\,
            lcout => data_in_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22924\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i7_LC_4_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__15106\,
            in1 => \N__14288\,
            in2 => \N__12064\,
            in3 => \N__17708\,
            lcout => rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22924\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_4_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110011001"
        )
    port map (
            in0 => \N__12639\,
            in1 => \N__12571\,
            in2 => \_gnd_net_\,
            in3 => \N__12476\,
            lcout => OPEN,
            ltout => \n3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_45_LC_4_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__12449\,
            in1 => \_gnd_net_\,
            in2 => \N__12341\,
            in3 => \N__14049\,
            lcout => tx2_o_adj_949,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22924\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i6_LC_4_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__17706\,
            in1 => \N__12334\,
            in2 => \N__14149\,
            in3 => \N__14287\,
            lcout => rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22924\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i0_LC_4_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17639\,
            in2 => \_gnd_net_\,
            in3 => \N__12323\,
            lcout => \c0.rx.r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22931\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17158\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => tx_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i54_LC_4_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17049\,
            in1 => \N__12272\,
            in2 => \_gnd_net_\,
            in3 => \N__12309\,
            lcout => data_in_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22931\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4166_3_lut_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__12248\,
            in1 => \N__12242\,
            in2 => \_gnd_net_\,
            in3 => \N__12236\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_325_326__i1_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15327\,
            in2 => \N__15495\,
            in3 => \_gnd_net_\,
            lcout => \c0.byte_transmit_counter2_0\,
            ltout => OPEN,
            carryin => \bfn_5_24_0_\,
            carryout => \c0.n3921\,
            clk => \N__22886\,
            ce => \N__12734\,
            sr => \N__12743\
        );

    \c0.byte_transmit_counter2_325_326__i2_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15608\,
            in2 => \_gnd_net_\,
            in3 => \N__12206\,
            lcout => \c0.byte_transmit_counter2_1\,
            ltout => OPEN,
            carryin => \c0.n3921\,
            carryout => \c0.n3922\,
            clk => \N__22886\,
            ce => \N__12734\,
            sr => \N__12743\
        );

    \c0.byte_transmit_counter2_325_326__i3_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15705\,
            in2 => \_gnd_net_\,
            in3 => \N__12746\,
            lcout => \c0.byte_transmit_counter2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22886\,
            ce => \N__12734\,
            sr => \N__12743\
        );

    \c0.i288_3_lut_4_lut_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100100111"
        )
    port map (
            in0 => \N__14404\,
            in1 => \N__12724\,
            in2 => \N__13100\,
            in3 => \N__12693\,
            lcout => \c0.n688\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i4_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21520\,
            in2 => \_gnd_net_\,
            in3 => \N__19457\,
            lcout => \c0.byte_transmit_counter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22892\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i7_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21519\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19847\,
            lcout => \c0.byte_transmit_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22892\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i6_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21521\,
            in2 => \_gnd_net_\,
            in3 => \N__19379\,
            lcout => \c0.byte_transmit_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22892\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i5_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21518\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19418\,
            lcout => \c0.byte_transmit_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22892\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2421_2_lut_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12723\,
            in2 => \_gnd_net_\,
            in3 => \N__12692\,
            lcout => \c0.n2643\,
            ltout => \c0.n2643_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_transmit_619_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100001011101"
        )
    port map (
            in0 => \N__14428\,
            in1 => \N__15328\,
            in2 => \N__12704\,
            in3 => \N__13098\,
            lcout => \c0.tx2_transmit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22892\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_351_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12665\,
            in1 => \N__13457\,
            in2 => \N__12659\,
            in3 => \N__12965\,
            lcout => OPEN,
            ltout => \c0.n30_adj_892_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2415_4_lut_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15026\,
            in1 => \N__12938\,
            in2 => \N__13109\,
            in3 => \N__13106\,
            lcout => \c0.n2637\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13075\,
            in1 => \N__13232\,
            in2 => \N__13046\,
            in3 => \N__13004\,
            lcout => OPEN,
            ltout => \c0.n16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__13571\,
            in1 => \N__12995\,
            in2 => \N__12983\,
            in3 => \N__12980\,
            lcout => \c0.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_348_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__12842\,
            in1 => \N__12959\,
            in2 => \N__12953\,
            in3 => \N__15932\,
            lcout => \c0.n26_adj_890\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i50_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__15037\,
            in1 => \N__12928\,
            in2 => \N__15852\,
            in3 => \N__14495\,
            lcout => \c0.data_in_frame_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22903\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_326_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12914\,
            in1 => \N__12899\,
            in2 => \N__14129\,
            in3 => \N__12866\,
            lcout => \c0.n4391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i42_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__15036\,
            in1 => \N__14494\,
            in2 => \N__14177\,
            in3 => \N__13189\,
            lcout => \c0.data_in_field_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22903\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_342_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13121\,
            in1 => \N__12835\,
            in2 => \N__12794\,
            in3 => \N__12758\,
            lcout => \c0.n12_adj_887\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i56_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13724\,
            in1 => \N__16998\,
            in2 => \_gnd_net_\,
            in3 => \N__13674\,
            lcout => data_in_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22903\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_319_LC_5_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13369\,
            in1 => \N__13341\,
            in2 => \N__13652\,
            in3 => \N__13608\,
            lcout => \c0.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_332_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13865\,
            in1 => \N__13120\,
            in2 => \N__13565\,
            in3 => \N__13535\,
            lcout => OPEN,
            ltout => \c0.n4415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_335_LC_5_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__16577\,
            in1 => \N__13304\,
            in2 => \N__13499\,
            in3 => \N__13485\,
            lcout => \c0.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_344_LC_5_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13443\,
            in1 => \N__13406\,
            in2 => \N__13831\,
            in3 => \N__13394\,
            lcout => \c0.n4421\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_adj_334_LC_5_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13250\,
            in1 => \N__13368\,
            in2 => \N__13298\,
            in3 => \N__13343\,
            lcout => \c0.n8_adj_883\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_301_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13293\,
            in2 => \_gnd_net_\,
            in3 => \N__13249\,
            lcout => \c0.n4441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_355_LC_5_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13214\,
            in1 => \N__13182\,
            in2 => \_gnd_net_\,
            in3 => \N__13147\,
            lcout => \c0.n4414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i52_LC_5_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16578\,
            in1 => \N__17096\,
            in2 => \_gnd_net_\,
            in3 => \N__14128\,
            lcout => data_in_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i55_LC_5_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16986\,
            in1 => \N__13928\,
            in2 => \_gnd_net_\,
            in3 => \N__14090\,
            lcout => data_in_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22918\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i41_LC_5_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16086\,
            in1 => \N__14271\,
            in2 => \_gnd_net_\,
            in3 => \N__16988\,
            lcout => data_in_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22918\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14056\,
            lcout => tx2_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_328_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14013\,
            in1 => \N__13964\,
            in2 => \N__13935\,
            in3 => \N__13896\,
            lcout => \c0.n12_adj_878\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i61_LC_5_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16987\,
            in1 => \N__13856\,
            in2 => \_gnd_net_\,
            in3 => \N__13820\,
            lcout => data_in_7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22918\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i24_LC_5_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__13796\,
            in1 => \N__15045\,
            in2 => \N__14685\,
            in3 => \N__13751\,
            lcout => \c0.data_in_field_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22918\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i36_LC_5_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16985\,
            in1 => \N__16561\,
            in2 => \_gnd_net_\,
            in3 => \N__14226\,
            lcout => data_in_4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22918\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i10_LC_5_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__15080\,
            in1 => \N__15044\,
            in2 => \N__14684\,
            in3 => \N__14310\,
            lcout => \c0.data_in_field_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22918\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i50_LC_5_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17265\,
            in1 => \N__16973\,
            in2 => \_gnd_net_\,
            in3 => \N__16752\,
            lcout => data_in_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2429_2_lut_LC_5_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16360\,
            in2 => \_gnd_net_\,
            in3 => \N__16393\,
            lcout => n2651,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i0_LC_5_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__16032\,
            in1 => \N__16158\,
            in2 => \_gnd_net_\,
            in3 => \N__16143\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i1_LC_5_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010001000"
        )
    port map (
            in0 => \N__16144\,
            in1 => \N__16361\,
            in2 => \N__16163\,
            in3 => \N__16033\,
            lcout => \c0.rx.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i33_LC_5_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17097\,
            in1 => \N__14272\,
            in2 => \_gnd_net_\,
            in3 => \N__14247\,
            lcout => data_in_4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i28_LC_5_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16971\,
            in1 => \N__14227\,
            in2 => \_gnd_net_\,
            in3 => \N__14201\,
            lcout => data_in_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i2_LC_5_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101000000000"
        )
    port map (
            in0 => \N__16394\,
            in1 => \N__16162\,
            in2 => \N__16004\,
            in3 => \N__16145\,
            lcout => \r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i43_LC_5_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16972\,
            in1 => \N__14161\,
            in2 => \_gnd_net_\,
            in3 => \N__15854\,
            lcout => data_in_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_4_lut_LC_5_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__15119\,
            in1 => \N__17557\,
            in2 => \N__16034\,
            in3 => \N__17637\,
            lcout => n1222,
            ltout => \n1222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i0_LC_5_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__15154\,
            in1 => \N__16327\,
            in2 => \N__15158\,
            in3 => \N__17709\,
            lcout => rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_27_i4_2_lut_LC_5_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__16396\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16363\,
            lcout => n4_adj_950,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_25_i4_2_lut_LC_5_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16362\,
            in2 => \_gnd_net_\,
            in3 => \N__16395\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_LC_5_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17756\,
            in2 => \_gnd_net_\,
            in3 => \N__17372\,
            lcout => \c0.rx.n2269\,
            ltout => \c0.rx.n2269_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_4_lut_adj_279_LC_5_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__16031\,
            in1 => \N__17558\,
            in2 => \N__15113\,
            in3 => \N__17638\,
            lcout => n1227,
            ltout => \n1227_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i1_LC_5_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__17287\,
            in1 => \N__16328\,
            in2 => \N__15092\,
            in3 => \N__17710\,
            lcout => rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_2_lut_LC_5_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16226\,
            in3 => \N__15089\,
            lcout => n226,
            ltout => OPEN,
            carryin => \bfn_5_32_0_\,
            carryout => \c0.rx.n3884\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_3_lut_LC_5_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16517\,
            in1 => \N__16306\,
            in2 => \_gnd_net_\,
            in3 => \N__15086\,
            lcout => \c0.rx.n4679\,
            ltout => OPEN,
            carryin => \c0.rx.n3884\,
            carryout => \c0.rx.n3885\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_4_lut_LC_5_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17423\,
            in2 => \_gnd_net_\,
            in3 => \N__15083\,
            lcout => n224,
            ltout => OPEN,
            carryin => \c0.rx.n3885\,
            carryout => \c0.rx.n3886\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_5_lut_LC_5_32_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16428\,
            in2 => \_gnd_net_\,
            in3 => \N__15260\,
            lcout => n223,
            ltout => OPEN,
            carryin => \c0.rx.n3886\,
            carryout => \c0.rx.n3887\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_6_lut_LC_5_32_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16180\,
            in2 => \_gnd_net_\,
            in3 => \N__15257\,
            lcout => n222,
            ltout => OPEN,
            carryin => \c0.rx.n3887\,
            carryout => \c0.rx.n3888\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_7_lut_LC_5_32_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16474\,
            in2 => \_gnd_net_\,
            in3 => \N__15254\,
            lcout => n221,
            ltout => OPEN,
            carryin => \c0.rx.n3888\,
            carryout => \c0.rx.n3889\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_8_lut_LC_5_32_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17855\,
            in2 => \_gnd_net_\,
            in3 => \N__15251\,
            lcout => n220,
            ltout => OPEN,
            carryin => \c0.rx.n3889\,
            carryout => \c0.rx.n3890\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_9_lut_LC_5_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16273\,
            in2 => \_gnd_net_\,
            in3 => \N__15248\,
            lcout => n219,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i1_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__22427\,
            in1 => \N__21540\,
            in2 => \_gnd_net_\,
            in3 => \N__21257\,
            lcout => data_out_field_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22887\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i6_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15245\,
            in2 => \_gnd_net_\,
            in3 => \N__15233\,
            lcout => \c0.tx2.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22887\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i0_LC_6_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18277\,
            in2 => \_gnd_net_\,
            in3 => \N__15164\,
            lcout => \c0.data_0\,
            ltout => OPEN,
            carryin => \bfn_6_25_0_\,
            carryout => \c0.n3906\,
            clk => \N__22897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i1_LC_6_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15898\,
            in2 => \_gnd_net_\,
            in3 => \N__15161\,
            lcout => \c0.data_1\,
            ltout => OPEN,
            carryin => \c0.n3906\,
            carryout => \c0.n3907\,
            clk => \N__22897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i2_LC_6_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19060\,
            in2 => \_gnd_net_\,
            in3 => \N__15287\,
            lcout => \c0.data_2\,
            ltout => OPEN,
            carryin => \c0.n3907\,
            carryout => \c0.n3908\,
            clk => \N__22897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i3_LC_6_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18613\,
            in2 => \_gnd_net_\,
            in3 => \N__15284\,
            lcout => \c0.data_3\,
            ltout => OPEN,
            carryin => \c0.n3908\,
            carryout => \c0.n3909\,
            clk => \N__22897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i4_LC_6_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18658\,
            in2 => \_gnd_net_\,
            in3 => \N__15281\,
            lcout => \c0.data_4\,
            ltout => OPEN,
            carryin => \c0.n3909\,
            carryout => \c0.n3910\,
            clk => \N__22897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i5_LC_6_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18814\,
            in2 => \_gnd_net_\,
            in3 => \N__15278\,
            lcout => \c0.data_5\,
            ltout => OPEN,
            carryin => \c0.n3910\,
            carryout => \c0.n3911\,
            clk => \N__22897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i6_LC_6_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18106\,
            in2 => \_gnd_net_\,
            in3 => \N__15275\,
            lcout => \c0.data_6\,
            ltout => OPEN,
            carryin => \c0.n3911\,
            carryout => \c0.n3912\,
            clk => \N__22897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i7_LC_6_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18088\,
            in2 => \_gnd_net_\,
            in3 => \N__15272\,
            lcout => \c0.data_7\,
            ltout => OPEN,
            carryin => \c0.n3912\,
            carryout => \c0.n3913\,
            clk => \N__22897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i8_LC_6_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18028\,
            in2 => \_gnd_net_\,
            in3 => \N__15269\,
            lcout => \c0.data_8\,
            ltout => OPEN,
            carryin => \bfn_6_26_0_\,
            carryout => \c0.n3914\,
            clk => \N__22904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i9_LC_6_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15301\,
            in2 => \_gnd_net_\,
            in3 => \N__15266\,
            lcout => \c0.data_9\,
            ltout => OPEN,
            carryin => \c0.n3914\,
            carryout => \c0.n3915\,
            clk => \N__22904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i10_LC_6_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18184\,
            in2 => \_gnd_net_\,
            in3 => \N__15263\,
            lcout => \c0.data_10\,
            ltout => OPEN,
            carryin => \c0.n3915\,
            carryout => \c0.n3916\,
            clk => \N__22904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i11_LC_6_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18634\,
            in2 => \_gnd_net_\,
            in3 => \N__15803\,
            lcout => \c0.data_11\,
            ltout => OPEN,
            carryin => \c0.n3916\,
            carryout => \c0.n3917\,
            clk => \N__22904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i12_LC_6_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19297\,
            in2 => \_gnd_net_\,
            in3 => \N__15800\,
            lcout => \c0.data_12\,
            ltout => OPEN,
            carryin => \c0.n3917\,
            carryout => \c0.n3918\,
            clk => \N__22904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i13_LC_6_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21619\,
            in2 => \_gnd_net_\,
            in3 => \N__15797\,
            lcout => \c0.data_13\,
            ltout => OPEN,
            carryin => \c0.n3918\,
            carryout => \c0.n3919\,
            clk => \N__22904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i14_LC_6_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18067\,
            in2 => \_gnd_net_\,
            in3 => \N__15794\,
            lcout => \c0.data_14\,
            ltout => OPEN,
            carryin => \c0.n3919\,
            carryout => \c0.n3920\,
            clk => \N__22904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_327__i15_LC_6_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17977\,
            in2 => \_gnd_net_\,
            in3 => \N__15791\,
            lcout => \c0.data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4401_3_lut_LC_6_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__15767\,
            in1 => \N__15637\,
            in2 => \_gnd_net_\,
            in3 => \N__15527\,
            lcout => \c0.FRAME_MATCHER_wait_for_transmission_N_423\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i34_LC_6_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__18894\,
            in1 => \N__21562\,
            in2 => \N__15305\,
            in3 => \N__21255\,
            lcout => \c0.data_out_field_47_N_682_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4264_3_lut_LC_6_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18383\,
            in1 => \N__20288\,
            in2 => \_gnd_net_\,
            in3 => \N__20551\,
            lcout => OPEN,
            ltout => \c0.n4619_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_4435_LC_6_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__20783\,
            in1 => \N__20693\,
            in2 => \N__15290\,
            in3 => \N__19565\,
            lcout => \c0.n4789\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i0_LC_6_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010000110000"
        )
    port map (
            in0 => \N__23249\,
            in1 => \N__21852\,
            in2 => \N__19210\,
            in3 => \N__23207\,
            lcout => \c0.tx.r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_318_LC_6_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18558\,
            in1 => \N__18172\,
            in2 => \_gnd_net_\,
            in3 => \N__18888\,
            lcout => \c0.n4380\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i42_LC_6_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__21256\,
            in1 => \N__18585\,
            in2 => \N__15905\,
            in3 => \N__21554\,
            lcout => \c0.data_out_field_47_N_682_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i51_LC_6_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16997\,
            in1 => \N__15845\,
            in2 => \_gnd_net_\,
            in3 => \N__15887\,
            lcout => data_in_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22919\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4162_3_lut_LC_6_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20550\,
            in1 => \N__18137\,
            in2 => \_gnd_net_\,
            in3 => \N__18233\,
            lcout => OPEN,
            ltout => \c0.n4517_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_LC_6_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__19589\,
            in1 => \N__15917\,
            in2 => \N__15818\,
            in3 => \N__20706\,
            lcout => OPEN,
            ltout => \c0.n4867_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4867_bdd_4_lut_LC_6_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__15809\,
            in1 => \N__18395\,
            in2 => \N__15815\,
            in3 => \N__19590\,
            lcout => OPEN,
            ltout => \tx_data_2_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i2_LC_6_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22116\,
            in2 => \N__15812\,
            in3 => \N__17191\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22919\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4209_3_lut_LC_6_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20549\,
            in1 => \N__22001\,
            in2 => \_gnd_net_\,
            in3 => \N__21680\,
            lcout => \c0.n4564\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_327_LC_6_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16087\,
            in1 => \N__15962\,
            in2 => \_gnd_net_\,
            in3 => \N__15950\,
            lcout => \c0.n4409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i4354_2_lut_LC_6_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__17363\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17618\,
            lcout => \c0.rx.n4677\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_2_lut_LC_6_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16225\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17856\,
            lcout => \c0.rx.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i223_3_lut_LC_6_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001000"
        )
    port map (
            in0 => \N__17419\,
            in1 => \N__16430\,
            in2 => \N__16310\,
            in3 => \_gnd_net_\,
            lcout => \c0.rx.n232\,
            ltout => \c0.rx.n232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i2_LC_6_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__15977\,
            in1 => \N__17857\,
            in2 => \N__15920\,
            in3 => \N__16277\,
            lcout => \c0.rx.r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22926\,
            ce => 'H',
            sr => \N__17330\
        );

    \c0.i4161_3_lut_LC_6_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20341\,
            in1 => \N__18563\,
            in2 => \_gnd_net_\,
            in3 => \N__20519\,
            lcout => \c0.n4516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4171_3_lut_LC_6_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18173\,
            in1 => \N__19772\,
            in2 => \_gnd_net_\,
            in3 => \N__20518\,
            lcout => \c0.n4526\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i13_4_lut_4_lut_LC_6_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100000101"
        )
    port map (
            in0 => \N__17553\,
            in1 => \N__17620\,
            in2 => \N__17789\,
            in3 => \N__17368\,
            lcout => OPEN,
            ltout => \c0.rx.n1464_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_52_LC_6_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__17621\,
            in1 => \N__16906\,
            in2 => \N__15908\,
            in3 => \N__17554\,
            lcout => rx_data_ready_keep,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22933\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_4_lut_4_lut_LC_6_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__17551\,
            in1 => \N__17619\,
            in2 => \N__17788\,
            in3 => \N__17367\,
            lcout => n1527,
            ltout => \n1527_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_3_lut_4_lut_LC_6_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100001111"
        )
    port map (
            in0 => \N__16392\,
            in1 => \N__16000\,
            in2 => \N__16148\,
            in3 => \N__17552\,
            lcout => n2142,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i49_LC_6_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16905\,
            in1 => \N__16085\,
            in2 => \_gnd_net_\,
            in3 => \N__16131\,
            lcout => data_in_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22933\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_adj_276_LC_6_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__17858\,
            in1 => \N__15973\,
            in2 => \N__16058\,
            in3 => \N__16272\,
            lcout => \c0.rx.r_SM_Main_2_N_816_2\,
            ltout => \c0.rx.r_SM_Main_2_N_816_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i4336_2_lut_3_lut_4_lut_LC_6_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16358\,
            in1 => \N__16026\,
            in2 => \N__16049\,
            in3 => \N__16391\,
            lcout => \c0.rx.n4678\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_274_LC_6_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16027\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16359\,
            lcout => n4_adj_943,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i3_LC_6_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__16429\,
            in1 => \N__17925\,
            in2 => \N__15989\,
            in3 => \N__17888\,
            lcout => \r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_289_LC_6_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18562\,
            in2 => \_gnd_net_\,
            in3 => \N__20198\,
            lcout => n4_adj_942,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_275_LC_6_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16473\,
            in2 => \_gnd_net_\,
            in3 => \N__16179\,
            lcout => \c0.rx.n214\,
            ltout => \c0.rx.n214_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_adj_268_LC_6_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16424\,
            in1 => \N__16270\,
            in2 => \N__16403\,
            in3 => \N__16304\,
            lcout => \c0.rx.n4\,
            ltout => \c0.rx.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_4_lut_LC_6_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__17837\,
            in1 => \N__16217\,
            in2 => \N__16400\,
            in3 => \N__17416\,
            lcout => \c0.rx.n2179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_28_i4_2_lut_LC_6_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__16397\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16364\,
            lcout => n4_adj_951,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i1_LC_6_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16305\,
            in1 => \N__16316\,
            in2 => \_gnd_net_\,
            in3 => \N__17924\,
            lcout => \c0.rx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i7_LC_6_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__17889\,
            in1 => \N__16283\,
            in2 => \N__17933\,
            in3 => \N__16271\,
            lcout => \r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2038_4_lut_LC_6_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__17306\,
            in1 => \N__16247\,
            in2 => \N__17550\,
            in3 => \N__16490\,
            lcout => n573,
            ltout => \n573_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i0_LC_6_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__16238\,
            in1 => \N__16224\,
            in2 => \N__16229\,
            in3 => \N__17929\,
            lcout => \r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i4_LC_6_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__17930\,
            in1 => \N__16184\,
            in2 => \N__16196\,
            in3 => \N__17886\,
            lcout => \r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i4353_3_lut_LC_6_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__17766\,
            in1 => \N__17685\,
            in2 => \_gnd_net_\,
            in3 => \N__17809\,
            lcout => OPEN,
            ltout => \c0.rx.n4641_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_adj_269_LC_6_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011111110"
        )
    port map (
            in0 => \N__17524\,
            in1 => \N__17632\,
            in2 => \N__16520\,
            in3 => \N__17374\,
            lcout => \c0.rx.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i4_4_lut_LC_6_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__16511\,
            in1 => \N__17417\,
            in2 => \N__16505\,
            in3 => \N__17304\,
            lcout => \c0.rx.n4093\,
            ltout => \c0.rx.n4093_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i82_3_lut_4_lut_LC_6_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111010001"
        )
    port map (
            in0 => \N__17305\,
            in1 => \N__17767\,
            in2 => \N__16493\,
            in3 => \N__17631\,
            lcout => \c0.rx.n2246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i5_LC_6_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__17887\,
            in1 => \N__17931\,
            in2 => \N__16484\,
            in3 => \N__16475\,
            lcout => \r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i25_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__21525\,
            in1 => \N__18314\,
            in2 => \_gnd_net_\,
            in3 => \N__21249\,
            lcout => data_out_field_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22898\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_4430_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__16607\,
            in1 => \N__19602\,
            in2 => \N__16439\,
            in3 => \N__20705\,
            lcout => OPEN,
            ltout => \c0.n4783_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4783_bdd_4_lut_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__19603\,
            in1 => \N__16601\,
            in2 => \N__16457\,
            in3 => \N__16454\,
            lcout => OPEN,
            ltout => \tx_data_3_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i3_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22151\,
            in2 => \N__16442\,
            in3 => \N__17206\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22905\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4267_3_lut_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20546\,
            in1 => \N__18056\,
            in2 => \_gnd_net_\,
            in3 => \N__18793\,
            lcout => \c0.n4622\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4266_3_lut_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21957\,
            in1 => \N__19822\,
            in2 => \_gnd_net_\,
            in3 => \N__20547\,
            lcout => \c0.n4621\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4170_3_lut_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20548\,
            in1 => \N__18479\,
            in2 => \_gnd_net_\,
            in3 => \N__18364\,
            lcout => \c0.n4525\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i44_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16548\,
            in1 => \N__17092\,
            in2 => \_gnd_net_\,
            in3 => \N__16591\,
            lcout => data_in_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4765_bdd_4_lut_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__20369\,
            in1 => \N__19286\,
            in2 => \N__21931\,
            in3 => \N__20708\,
            lcout => OPEN,
            ltout => \c0.n4768_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i277446_i1_3_lut_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17963\,
            in2 => \N__16532\,
            in3 => \N__19585\,
            lcout => OPEN,
            ltout => \tx_data_7_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i7_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22150\,
            in2 => \N__16529\,
            in3 => \N__16658\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_4488_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__16646\,
            in1 => \N__19566\,
            in2 => \N__16625\,
            in3 => \N__20694\,
            lcout => OPEN,
            ltout => \c0.n4843_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4843_bdd_4_lut_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__19567\,
            in1 => \N__19082\,
            in2 => \N__16526\,
            in3 => \N__18245\,
            lcout => OPEN,
            ltout => \tx_data_1_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i1_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22141\,
            in2 => \N__16523\,
            in3 => \N__17236\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22920\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4234_3_lut_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19185\,
            in1 => \N__16657\,
            in2 => \_gnd_net_\,
            in3 => \N__16639\,
            lcout => \c0.tx.n4589\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4230_3_lut_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18887\,
            in1 => \N__18584\,
            in2 => \_gnd_net_\,
            in3 => \N__20554\,
            lcout => \c0.n4585\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1361_2_lut_LC_7_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__23244\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23205\,
            lcout => \c0.tx.n1588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i6_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16640\,
            in1 => \N__22142\,
            in2 => \_gnd_net_\,
            in3 => \N__19334\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22920\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_4493_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__16712\,
            in1 => \N__19596\,
            in2 => \N__19676\,
            in3 => \N__20701\,
            lcout => OPEN,
            ltout => \c0.n4861_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4861_bdd_4_lut_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__19597\,
            in1 => \N__16616\,
            in2 => \N__16631\,
            in3 => \N__18200\,
            lcout => OPEN,
            ltout => \tx_data_0_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i0_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22114\,
            in2 => \N__16628\,
            in3 => \N__17221\,
            lcout => \r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22927\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4231_3_lut_LC_7_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18214\,
            in1 => \N__17999\,
            in2 => \_gnd_net_\,
            in3 => \N__20553\,
            lcout => \c0.n4586\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4233_3_lut_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19199\,
            in1 => \N__16687\,
            in2 => \_gnd_net_\,
            in3 => \N__16723\,
            lcout => \c0.tx.n4588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4218_3_lut_LC_7_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22431\,
            in1 => \N__22232\,
            in2 => \_gnd_net_\,
            in3 => \N__20552\,
            lcout => \c0.n4573\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4789_bdd_4_lut_LC_7_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101111001000"
        )
    port map (
            in0 => \N__18419\,
            in1 => \N__16733\,
            in2 => \N__19604\,
            in3 => \N__17387\,
            lcout => OPEN,
            ltout => \tx_data_4_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i4_LC_7_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__22115\,
            in1 => \_gnd_net_\,
            in2 => \N__16727\,
            in3 => \N__16724\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22927\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4221_3_lut_LC_7_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19112\,
            in1 => \N__18515\,
            in2 => \_gnd_net_\,
            in3 => \N__20516\,
            lcout => \c0.n4576\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_1__bdd_4_lut_LC_7_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__19226\,
            in1 => \N__16706\,
            in2 => \N__19261\,
            in3 => \N__16697\,
            lcout => \c0.tx.n4837\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4795_bdd_4_lut_LC_7_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__20084\,
            in1 => \N__18998\,
            in2 => \N__19721\,
            in3 => \N__19601\,
            lcout => OPEN,
            ltout => \tx_data_5_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i5_LC_7_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__22143\,
            in1 => \_gnd_net_\,
            in2 => \N__16691\,
            in3 => \N__16688\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i1_LC_7_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001110000000"
        )
    port map (
            in0 => \N__19209\,
            in1 => \N__21853\,
            in2 => \N__16676\,
            in3 => \N__19228\,
            lcout => \c0.tx.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4360_2_lut_LC_7_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19227\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19208\,
            lcout => OPEN,
            ltout => \c0.tx.n4715_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i2_LC_7_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101110000000"
        )
    port map (
            in0 => \N__16675\,
            in1 => \N__21854\,
            in2 => \N__16661\,
            in3 => \N__19256\,
            lcout => \c0.tx.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i58_LC_7_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16970\,
            in1 => \N__17294\,
            in2 => \_gnd_net_\,
            in3 => \N__17261\,
            lcout => data_in_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22939\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_375_LC_7_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19139\,
            in1 => \N__18365\,
            in2 => \N__21740\,
            in3 => \N__19768\,
            lcout => n4_adj_970,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4203_3_lut_LC_7_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17237\,
            in1 => \N__17222\,
            in2 => \_gnd_net_\,
            in3 => \N__19206\,
            lcout => \c0.tx.n4558\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_LC_7_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19767\,
            in2 => \_gnd_net_\,
            in3 => \N__19132\,
            lcout => \c0.n1333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4204_3_lut_LC_7_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17207\,
            in1 => \N__17192\,
            in2 => \_gnd_net_\,
            in3 => \N__19207\,
            lcout => OPEN,
            ltout => \c0.tx.n4559_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.n4837_bdd_4_lut_LC_7_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__19257\,
            in1 => \N__17177\,
            in2 => \N__17171\,
            in3 => \N__17168\,
            lcout => \c0.tx.o_Tx_Serial_N_790\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i26_LC_7_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__21560\,
            in1 => \N__19140\,
            in2 => \_gnd_net_\,
            in3 => \N__21259\,
            lcout => data_out_field_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22939\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_45_LC_7_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__17145\,
            in1 => \N__23501\,
            in2 => \_gnd_net_\,
            in3 => \N__17315\,
            lcout => tx_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i42_LC_7_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16907\,
            in1 => \N__17451\,
            in2 => \_gnd_net_\,
            in3 => \N__16763\,
            lcout => data_in_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i2_LC_7_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__17418\,
            in1 => \N__17932\,
            in2 => \N__17438\,
            in3 => \N__17891\,
            lcout => \r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4173_3_lut_LC_7_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20150\,
            in1 => \N__18452\,
            in2 => \_gnd_net_\,
            in3 => \N__20555\,
            lcout => \c0.n4528\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i4346_2_lut_LC_7_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17780\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17373\,
            lcout => \c0.rx.n4667\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i13_LC_7_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__20151\,
            in1 => \N__21561\,
            in2 => \_gnd_net_\,
            in3 => \N__21260\,
            lcout => data_out_field_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i4404_2_lut_3_lut_LC_7_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__17781\,
            in1 => \N__17633\,
            in2 => \_gnd_net_\,
            in3 => \N__17542\,
            lcout => \c0.rx.n1024\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i26_3_lut_LC_7_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001100110"
        )
    port map (
            in0 => \N__23206\,
            in1 => \N__23018\,
            in2 => \_gnd_net_\,
            in3 => \N__17321\,
            lcout => \c0.tx.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_277_LC_7_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__17762\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17517\,
            lcout => \c0.rx.n4378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_2_lut_adj_271_LC_7_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17684\,
            in2 => \_gnd_net_\,
            in3 => \N__17807\,
            lcout => \c0.rx.n6\,
            ltout => \c0.rx.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_adj_272_LC_7_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__17760\,
            in1 => \N__17516\,
            in2 => \N__17309\,
            in3 => \N__17627\,
            lcout => \c0.rx.n357\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_4_lut_adj_278_LC_7_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__17628\,
            in1 => \N__17761\,
            in2 => \N__17544\,
            in3 => \N__17954\,
            lcout => OPEN,
            ltout => \c0.rx.n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_adj_273_LC_7_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110011"
        )
    port map (
            in0 => \N__17948\,
            in1 => \N__17629\,
            in2 => \N__17942\,
            in3 => \N__17939\,
            lcout => n1554,
            ltout => \n1554_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i6_LC_7_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__17900\,
            in1 => \N__17890\,
            in2 => \N__17861\,
            in3 => \N__17846\,
            lcout => \r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22951\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i4356_3_lut_LC_7_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101111"
        )
    port map (
            in0 => \N__17808\,
            in1 => \_gnd_net_\,
            in2 => \N__17779\,
            in3 => \N__17687\,
            lcout => OPEN,
            ltout => \c0.rx.n4666_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i1_LC_7_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000101000101"
        )
    port map (
            in0 => \N__17630\,
            in1 => \N__17543\,
            in2 => \N__17567\,
            in3 => \N__17564\,
            lcout => \c0.rx.r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22951\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_328__i0_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18122\,
            in2 => \N__18764\,
            in3 => \_gnd_net_\,
            lcout => \c0.delay_counter_0\,
            ltout => OPEN,
            carryin => \bfn_9_25_0_\,
            carryout => \c0.n3899\,
            clk => \N__22921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_328__i1_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18710\,
            in2 => \_gnd_net_\,
            in3 => \N__17474\,
            lcout => \c0.delay_counter_1\,
            ltout => OPEN,
            carryin => \c0.n3899\,
            carryout => \c0.n3900\,
            clk => \N__22921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_328__i2_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18748\,
            in2 => \_gnd_net_\,
            in3 => \N__17471\,
            lcout => \c0.delay_counter_2\,
            ltout => OPEN,
            carryin => \c0.n3900\,
            carryout => \c0.n3901\,
            clk => \N__22921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_328__i3_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18683\,
            in2 => \_gnd_net_\,
            in3 => \N__18014\,
            lcout => \c0.delay_counter_3\,
            ltout => OPEN,
            carryin => \c0.n3901\,
            carryout => \c0.n3902\,
            clk => \N__22921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_328__i4_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18734\,
            in2 => \_gnd_net_\,
            in3 => \N__18011\,
            lcout => \c0.delay_counter_4\,
            ltout => OPEN,
            carryin => \c0.n3902\,
            carryout => \c0.n3903\,
            clk => \N__22921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_328__i5_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18722\,
            in2 => \_gnd_net_\,
            in3 => \N__18008\,
            lcout => \c0.delay_counter_5\,
            ltout => OPEN,
            carryin => \c0.n3903\,
            carryout => \c0.n3904\,
            clk => \N__22921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_328__i6_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18776\,
            in2 => \_gnd_net_\,
            in3 => \N__18005\,
            lcout => \c0.delay_counter_6\,
            ltout => OPEN,
            carryin => \c0.n3904\,
            carryout => \c0.n3905\,
            clk => \N__22921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_328__i7_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18697\,
            in2 => \_gnd_net_\,
            in3 => \N__18002\,
            lcout => \c0.delay_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i50_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__21577\,
            in1 => \N__17995\,
            in2 => \N__20723\,
            in3 => \N__21136\,
            lcout => data_out_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i40_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__21133\,
            in1 => \N__17981\,
            in2 => \N__21735\,
            in3 => \N__21583\,
            lcout => \c0.data_out_field_47_N_682_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4885_bdd_4_lut_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__22324\,
            in1 => \N__21724\,
            in2 => \N__18830\,
            in3 => \N__20707\,
            lcout => \c0.n4888\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_transmit_612_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__22270\,
            in1 => \N__22458\,
            in2 => \_gnd_net_\,
            in3 => \N__21213\,
            lcout => \c0.tx_transmit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_340_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__22457\,
            in1 => \N__21131\,
            in2 => \_gnd_net_\,
            in3 => \N__22269\,
            lcout => \c0.n2429\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i47_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__21134\,
            in1 => \N__21579\,
            in2 => \N__18116\,
            in3 => \N__19877\,
            lcout => \c0.data_out_field_47_N_682_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i48_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__22325\,
            in1 => \N__18095\,
            in2 => \N__21584\,
            in3 => \N__21135\,
            lcout => \c0.data_out_field_47_N_682_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i39_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__21132\,
            in1 => \N__21578\,
            in2 => \N__18077\,
            in3 => \N__21814\,
            lcout => data_out_field_38,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i27_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__21542\,
            in1 => \N__22042\,
            in2 => \_gnd_net_\,
            in3 => \N__21145\,
            lcout => data_out_field_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22935\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i60_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001001110"
        )
    port map (
            in0 => \N__21148\,
            in1 => \N__18055\,
            in2 => \N__22301\,
            in3 => \N__21545\,
            lcout => data_out_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22935\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i12_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__21541\,
            in1 => \N__18356\,
            in2 => \_gnd_net_\,
            in3 => \N__21144\,
            lcout => data_out_field_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22935\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i33_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__21147\,
            in1 => \N__18508\,
            in2 => \N__18038\,
            in3 => \N__21544\,
            lcout => \c0.data_out_field_47_N_682_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22935\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_adj_359_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20583\,
            in1 => \N__20882\,
            in2 => \_gnd_net_\,
            in3 => \N__22547\,
            lcout => OPEN,
            ltout => \n8_adj_932_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i59_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011010"
        )
    port map (
            in0 => \N__18602\,
            in1 => \N__18229\,
            in2 => \N__18017\,
            in3 => \N__20070\,
            lcout => data_out_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22935\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i5_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__21543\,
            in1 => \N__18450\,
            in2 => \_gnd_net_\,
            in3 => \N__21146\,
            lcout => data_out_field_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22935\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21692\,
            in1 => \N__18328\,
            in2 => \_gnd_net_\,
            in3 => \N__20816\,
            lcout => n8_adj_936,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i32_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__21537\,
            in1 => \_gnd_net_\,
            in2 => \N__20590\,
            in3 => \N__21178\,
            lcout => data_out_field_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i58_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__20056\,
            in1 => \N__18215\,
            in2 => \N__19322\,
            in3 => \N__19004\,
            lcout => data_out_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i18_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__21536\,
            in1 => \N__18265\,
            in2 => \_gnd_net_\,
            in3 => \N__21176\,
            lcout => data_out_field_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4219_3_lut_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18327\,
            in1 => \N__18964\,
            in2 => \_gnd_net_\,
            in3 => \N__20495\,
            lcout => \c0.n4574\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i35_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__21538\,
            in1 => \N__18191\,
            in2 => \N__18557\,
            in3 => \N__21179\,
            lcout => \c0.data_out_field_47_N_682_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i20_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__21177\,
            in1 => \N__18165\,
            in2 => \_gnd_net_\,
            in3 => \N__21539\,
            lcout => data_out_field_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i51_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__18143\,
            in1 => \N__18136\,
            in2 => \N__20075\,
            in3 => \N__18407\,
            lcout => data_out_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4210_3_lut_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22031\,
            in1 => \N__20235\,
            in2 => \_gnd_net_\,
            in3 => \N__20496\,
            lcout => \c0.n4565\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_385_LC_9_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20578\,
            in1 => \N__18261\,
            in2 => \_gnd_net_\,
            in3 => \N__18509\,
            lcout => \c0.n1312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_3_lut_4_lut_adj_384_LC_9_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18510\,
            in1 => \N__20579\,
            in2 => \N__20237\,
            in3 => \N__18475\,
            lcout => OPEN,
            ltout => \n11_adj_967_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i61_LC_9_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110100100001"
        )
    port map (
            in0 => \N__18857\,
            in1 => \N__20062\,
            in2 => \N__18386\,
            in3 => \N__18379\,
            lcout => data_out_7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22946\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_LC_9_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21815\,
            in1 => \N__18357\,
            in2 => \_gnd_net_\,
            in3 => \N__21728\,
            lcout => OPEN,
            ltout => \c0.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_LC_9_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21672\,
            in1 => \N__22038\,
            in2 => \N__18332\,
            in3 => \N__18329\,
            lcout => \c0.n4456\,
            ltout => \c0.n4456_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_386_LC_9_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18592\,
            in2 => \N__18290\,
            in3 => \N__19105\,
            lcout => n1255,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i41_LC_9_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__19106\,
            in1 => \N__21576\,
            in2 => \N__18287\,
            in3 => \N__21246\,
            lcout => \c0.data_out_field_47_N_682_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22946\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4207_3_lut_LC_9_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20494\,
            in1 => \N__18266\,
            in2 => \_gnd_net_\,
            in3 => \N__19142\,
            lcout => \c0.n4562\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_LC_9_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18596\,
            in1 => \N__19110\,
            in2 => \N__20345\,
            in3 => \N__20162\,
            lcout => n4462,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i4_LC_9_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__21242\,
            in1 => \N__18471\,
            in2 => \_gnd_net_\,
            in3 => \N__21524\,
            lcout => data_out_field_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22952\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_364_LC_9_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18556\,
            in2 => \_gnd_net_\,
            in3 => \N__18901\,
            lcout => OPEN,
            ltout => \c0.n1384_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_350_LC_9_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19886\,
            in1 => \N__18446\,
            in2 => \N__18518\,
            in3 => \N__18511\,
            lcout => n10_adj_947,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_365_LC_9_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18470\,
            in1 => \N__18926\,
            in2 => \N__18451\,
            in3 => \N__22348\,
            lcout => \c0.n4465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4174_3_lut_LC_9_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20891\,
            in1 => \N__20194\,
            in2 => \_gnd_net_\,
            in3 => \N__20493\,
            lcout => \c0.n4529\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i14_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__20913\,
            in1 => \N__21522\,
            in2 => \_gnd_net_\,
            in3 => \N__21258\,
            lcout => data_out_field_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22906\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i10_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__21433\,
            in1 => \N__21768\,
            in2 => \_gnd_net_\,
            in3 => \N__21234\,
            lcout => data_out_field_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19632\,
            in2 => \_gnd_net_\,
            in3 => \N__22231\,
            lcout => n7_adj_937,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i16_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__21917\,
            in1 => \N__21444\,
            in2 => \_gnd_net_\,
            in3 => \N__21214\,
            lcout => data_out_field_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22922\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_374_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18775\,
            in1 => \N__18760\,
            in2 => \N__18749\,
            in3 => \N__18733\,
            lcout => \c0.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_373_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18721\,
            in1 => \N__18709\,
            in2 => \N__18698\,
            in3 => \N__18682\,
            lcout => OPEN,
            ltout => \c0.n14_adj_902_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22459\,
            in1 => \N__18671\,
            in2 => \N__18665\,
            in3 => \N__22271\,
            lcout => n3580,
            ltout => \n3580_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i45_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__20849\,
            in1 => \N__18662\,
            in2 => \N__18647\,
            in3 => \N__21215\,
            lcout => \c0.data_out_field_47_N_682_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22922\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i36_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__21436\,
            in1 => \N__19821\,
            in2 => \N__18644\,
            in3 => \N__21152\,
            lcout => \c0.data_out_field_47_N_682_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i44_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__21153\,
            in1 => \N__21956\,
            in2 => \N__18623\,
            in3 => \N__21438\,
            lcout => data_out_field_43,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21891\,
            in1 => \N__18966\,
            in2 => \_gnd_net_\,
            in3 => \N__19876\,
            lcout => n7_adj_933,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_363_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21992\,
            in2 => \_gnd_net_\,
            in3 => \N__21890\,
            lcout => \c0.n4393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i23_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__21434\,
            in1 => \N__19633\,
            in2 => \_gnd_net_\,
            in3 => \N__21149\,
            lcout => data_out_field_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__18845\,
            in1 => \N__20644\,
            in2 => \N__19037\,
            in3 => \N__20438\,
            lcout => \c0.n4885\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i29_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__21435\,
            in1 => \N__20883\,
            in2 => \_gnd_net_\,
            in3 => \N__21150\,
            lcout => data_out_field_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i31_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__21151\,
            in1 => \N__21892\,
            in2 => \_gnd_net_\,
            in3 => \N__21437\,
            lcout => data_out_field_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i46_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__21143\,
            in1 => \N__18821\,
            in2 => \N__21526\,
            in3 => \N__19945\,
            lcout => \c0.data_out_field_47_N_682_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i17_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__18967\,
            in1 => \N__21464\,
            in2 => \_gnd_net_\,
            in3 => \N__21142\,
            lcout => data_out_field_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_376_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19483\,
            in2 => \_gnd_net_\,
            in3 => \N__19837\,
            lcout => OPEN,
            ltout => \c0.n6_adj_904_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_377_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19447\,
            in1 => \N__19408\,
            in2 => \N__18803\,
            in3 => \N__19369\,
            lcout => n7_adj_938,
            ltout => \n7_adj_938_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i52_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__21462\,
            in1 => \N__21644\,
            in2 => \N__18800\,
            in3 => \N__18797\,
            lcout => data_out_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i11_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__21671\,
            in1 => \N__21463\,
            in2 => \_gnd_net_\,
            in3 => \N__21141\,
            lcout => data_out_field_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_370_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18925\,
            in1 => \N__19817\,
            in2 => \_gnd_net_\,
            in3 => \N__20809\,
            lcout => n7_adj_935,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_356_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20856\,
            in1 => \N__18905\,
            in2 => \N__18866\,
            in3 => \N__18965\,
            lcout => n12_adj_966,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_379_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21448\,
            in2 => \_gnd_net_\,
            in3 => \N__21137\,
            lcout => n1677,
            ltout => \n1677_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i56_LC_10_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__22490\,
            in1 => \N__18844\,
            in2 => \N__18848\,
            in3 => \N__18989\,
            lcout => data_out_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i22_LC_10_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__20759\,
            in1 => \N__21449\,
            in2 => \_gnd_net_\,
            in3 => \N__21139\,
            lcout => data_out_field_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i21_LC_10_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__21138\,
            in1 => \N__21466\,
            in2 => \_gnd_net_\,
            in3 => \N__20193\,
            lcout => data_out_field_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i6_LC_10_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__21465\,
            in1 => \N__20263\,
            in2 => \_gnd_net_\,
            in3 => \N__21140\,
            lcout => data_out_field_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_366_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20755\,
            in2 => \_gnd_net_\,
            in3 => \N__22329\,
            lcout => \c0.n4483\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_LC_10_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22330\,
            in1 => \N__19664\,
            in2 => \N__20764\,
            in3 => \N__20262\,
            lcout => OPEN,
            ltout => \n8_adj_934_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i64_LC_10_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100101"
        )
    port map (
            in0 => \N__19046\,
            in1 => \N__19033\,
            in2 => \N__19040\,
            in3 => \N__20063\,
            lcout => data_out_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_361_LC_10_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19019\,
            in1 => \N__20299\,
            in2 => \N__20990\,
            in3 => \N__20092\,
            lcout => \c0.n4447\,
            ltout => \c0.n4447_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_LC_10_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19007\,
            in3 => \N__19982\,
            lcout => n9_adj_972,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_4473_LC_10_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__20689\,
            in1 => \N__19148\,
            in2 => \N__19568\,
            in3 => \N__19922\,
            lcout => \c0.n4795\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_3_lut_4_lut_LC_10_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20093\,
            in1 => \N__20858\,
            in2 => \N__19955\,
            in3 => \N__19983\,
            lcout => n11_adj_945,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i54_LC_10_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011000000110"
        )
    port map (
            in0 => \N__22063\,
            in1 => \N__18980\,
            in2 => \N__20074\,
            in3 => \N__19160\,
            lcout => data_out_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22947\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_368_LC_10_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19878\,
            in2 => \_gnd_net_\,
            in3 => \N__18968\,
            lcout => \c0.n4417\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_383_LC_10_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19984\,
            in1 => \N__19953\,
            in2 => \_gnd_net_\,
            in3 => \N__18935\,
            lcout => OPEN,
            ltout => \n7_adj_969_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i57_LC_10_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111000010100"
        )
    port map (
            in0 => \N__20055\,
            in1 => \N__19706\,
            in2 => \N__18929\,
            in3 => \N__19697\,
            lcout => data_out_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22947\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i19_LC_10_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__21523\,
            in1 => \N__20234\,
            in2 => \_gnd_net_\,
            in3 => \N__21238\,
            lcout => data_out_field_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22953\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_3_lut_LC_10_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19265\,
            in1 => \N__19235\,
            in2 => \_gnd_net_\,
            in3 => \N__19211\,
            lcout => \c0.tx.n84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4261_3_lut_LC_10_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19966\,
            in1 => \N__19159\,
            in2 => \_gnd_net_\,
            in3 => \N__20479\,
            lcout => \c0.n4616\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_287_LC_10_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19141\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19111\,
            lcout => n4480,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4206_3_lut_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20989\,
            in1 => \N__21767\,
            in2 => \_gnd_net_\,
            in3 => \N__20478\,
            lcout => \c0.n4561\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i43_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__21248\,
            in1 => \N__20328\,
            in2 => \N__19067\,
            in3 => \N__21447\,
            lcout => \c0.data_out_field_47_N_682_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i3_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__21996\,
            in1 => \N__21445\,
            in2 => \_gnd_net_\,
            in3 => \N__21247\,
            lcout => data_out_field_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_4502_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__20477\,
            in1 => \N__21872\,
            in2 => \N__19634\,
            in3 => \N__20681\,
            lcout => OPEN,
            ltout => \c0.n4771_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4771_bdd_4_lut_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__20682\,
            in1 => \N__20360\,
            in2 => \N__19049\,
            in3 => \N__19657\,
            lcout => OPEN,
            ltout => \c0.n4774_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i276843_i1_3_lut_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20930\,
            in2 => \N__19337\,
            in3 => \N__19561\,
            lcout => tx_data_6_keep,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_360_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22081\,
            in1 => \N__22391\,
            in2 => \N__22000\,
            in3 => \N__20845\,
            lcout => n10_adj_971,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i8_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__19281\,
            in1 => \N__21446\,
            in2 => \_gnd_net_\,
            in3 => \N__21184\,
            lcout => data_out_field_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i7_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__21183\,
            in1 => \N__21442\,
            in2 => \_gnd_net_\,
            in3 => \N__19656\,
            lcout => data_out_field_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i37_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__21440\,
            in1 => \N__20807\,
            in2 => \N__19307\,
            in3 => \N__21185\,
            lcout => \c0.data_out_field_47_N_682_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i3_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21441\,
            in2 => \_gnd_net_\,
            in3 => \N__19484\,
            lcout => \c0.byte_transmit_counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i2_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__21439\,
            in1 => \N__20984\,
            in2 => \_gnd_net_\,
            in3 => \N__21182\,
            lcout => data_out_field_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i55_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__21186\,
            in1 => \N__19916\,
            in2 => \N__22010\,
            in3 => \N__21443\,
            lcout => data_out_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_380_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21602\,
            in1 => \N__19813\,
            in2 => \N__19285\,
            in3 => \N__20806\,
            lcout => n1246,
            ltout => \n1246_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19655\,
            in2 => \N__19637\,
            in3 => \N__19628\,
            lcout => n4438,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i0_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22283\,
            in2 => \N__20453\,
            in3 => \N__20054\,
            lcout => \c0.byte_transmit_counter_0\,
            ltout => OPEN,
            carryin => \bfn_11_27_0_\,
            carryout => \c0.n3844\,
            clk => \N__22942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i1_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20053\,
            in1 => \N__20643\,
            in2 => \_gnd_net_\,
            in3 => \N__19607\,
            lcout => \c0.byte_transmit_counter_1\,
            ltout => OPEN,
            carryin => \c0.n3844\,
            carryout => \c0.n3845\,
            clk => \N__22942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i2_LC_11_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20061\,
            in1 => \N__19522\,
            in2 => \_gnd_net_\,
            in3 => \N__19493\,
            lcout => \c0.byte_transmit_counter_2\,
            ltout => OPEN,
            carryin => \c0.n3845\,
            carryout => \c0.n3846\,
            clk => \N__22942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_637_5_lut_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19490\,
            in2 => \_gnd_net_\,
            in3 => \N__19472\,
            lcout => \c0.tx_transmit_N_274_3\,
            ltout => OPEN,
            carryin => \c0.n3846\,
            carryout => \c0.n3847\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_637_6_lut_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19469\,
            in2 => \_gnd_net_\,
            in3 => \N__19436\,
            lcout => \c0.tx_transmit_N_274_4\,
            ltout => OPEN,
            carryin => \c0.n3847\,
            carryout => \c0.n3848\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_637_7_lut_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19433\,
            in2 => \_gnd_net_\,
            in3 => \N__19397\,
            lcout => \c0.tx_transmit_N_274_5\,
            ltout => OPEN,
            carryin => \c0.n3848\,
            carryout => \c0.n3849\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_637_8_lut_LC_11_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19394\,
            in2 => \_gnd_net_\,
            in3 => \N__19358\,
            lcout => \c0.tx_transmit_N_274_6\,
            ltout => OPEN,
            carryin => \c0.n3849\,
            carryout => \c0.n3850\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_637_9_lut_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19355\,
            in2 => \_gnd_net_\,
            in3 => \N__19340\,
            lcout => \c0.tx_transmit_N_274_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_4_lut_LC_11_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20236\,
            in1 => \N__20192\,
            in2 => \N__20264\,
            in3 => \N__19826\,
            lcout => OPEN,
            ltout => \n9_adj_948_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i63_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101101000001"
        )
    port map (
            in0 => \N__20057\,
            in1 => \N__19787\,
            in2 => \N__19775\,
            in3 => \N__19903\,
            lcout => data_out_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i24_LC_11_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__21485\,
            in1 => \N__22192\,
            in2 => \_gnd_net_\,
            in3 => \N__21180\,
            lcout => data_out_field_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i28_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__21181\,
            in1 => \N__19758\,
            in2 => \_gnd_net_\,
            in3 => \N__21486\,
            lcout => data_out_field_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i49_LC_11_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111100"
        )
    port map (
            in0 => \N__19685\,
            in1 => \N__20108\,
            in2 => \N__19736\,
            in3 => \N__20058\,
            lcout => data_out_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4176_3_lut_LC_11_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20923\,
            in1 => \N__20452\,
            in2 => \_gnd_net_\,
            in3 => \N__20258\,
            lcout => \c0.n4531\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_adj_362_LC_11_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22373\,
            in1 => \N__22439\,
            in2 => \_gnd_net_\,
            in3 => \N__20924\,
            lcout => n8_adj_968,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4222_3_lut_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19696\,
            in1 => \N__20451\,
            in2 => \_gnd_net_\,
            in3 => \N__19684\,
            lcout => \c0.n4577\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i53_LC_11_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__20284\,
            in1 => \_gnd_net_\,
            in2 => \N__20306\,
            in3 => \N__20060\,
            lcout => data_out_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22954\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_367_LC_11_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20257\,
            in1 => \N__20224\,
            in2 => \_gnd_net_\,
            in3 => \N__20185\,
            lcout => OPEN,
            ltout => \c0.n4432_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_369_LC_11_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21775\,
            in1 => \N__20161\,
            in2 => \N__20129\,
            in3 => \N__20126\,
            lcout => OPEN,
            ltout => \c0.n10_adj_900_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_371_LC_11_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20120\,
            in1 => \N__22162\,
            in2 => \N__20111\,
            in3 => \N__20107\,
            lcout => \c0.n4489\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4177_3_lut_LC_11_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20954\,
            in1 => \N__20760\,
            in2 => \_gnd_net_\,
            in3 => \N__20466\,
            lcout => \c0.n4532\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i62_LC_11_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__20059\,
            in1 => \N__19967\,
            in2 => \N__19954\,
            in3 => \N__19991\,
            lcout => \c0.data_out_7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22954\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4260_3_lut_LC_11_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21608\,
            in1 => \N__19946\,
            in2 => \_gnd_net_\,
            in3 => \N__20465\,
            lcout => \c0.n4615\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_4507_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__19915\,
            in1 => \N__20679\,
            in2 => \N__20517\,
            in3 => \N__19904\,
            lcout => OPEN,
            ltout => \c0.n4879_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n4879_bdd_4_lut_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__20680\,
            in1 => \N__21823\,
            in2 => \N__19889\,
            in3 => \N__19885\,
            lcout => \c0.n4882\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_290_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21918\,
            in1 => \N__21990\,
            in2 => \_gnd_net_\,
            in3 => \N__21893\,
            lcout => \c0.n1378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_387_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20922\,
            in2 => \_gnd_net_\,
            in3 => \N__20890\,
            lcout => n4423,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i15_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__20359\,
            in1 => \N__21555\,
            in2 => \_gnd_net_\,
            in3 => \N__21250\,
            lcout => data_out_field_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22943\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4263_3_lut_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20423\,
            in1 => \N__20857\,
            in2 => \_gnd_net_\,
            in3 => \N__20808\,
            lcout => \c0.n4618\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4368_4_lut_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20768\,
            in1 => \N__22166\,
            in2 => \N__20735\,
            in3 => \N__21822\,
            lcout => n4663,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i30_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__21251\,
            in1 => \N__20950\,
            in2 => \_gnd_net_\,
            in3 => \N__21559\,
            lcout => data_out_field_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22943\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_4417_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__22193\,
            in1 => \N__20660\,
            in2 => \N__20594\,
            in3 => \N__20424\,
            lcout => \c0.n4765\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_372_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20358\,
            in2 => \_gnd_net_\,
            in3 => \N__20327\,
            lcout => \c0.n1421\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4372_4_lut_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21959\,
            in1 => \N__22082\,
            in2 => \N__22067\,
            in3 => \N__22043\,
            lcout => n4655,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21991\,
            in1 => \N__21958\,
            in2 => \N__21935\,
            in3 => \N__21889\,
            lcout => \c0.n4453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__23014\,
            in1 => \N__23453\,
            in2 => \N__23201\,
            in3 => \N__23069\,
            lcout => \c0.tx.n1514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21824\,
            in1 => \N__21606\,
            in2 => \N__21779\,
            in3 => \N__21736\,
            lcout => n4426,
            ltout => \n4426_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4370_4_lut_LC_12_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22191\,
            in1 => \N__22525\,
            in2 => \N__21683\,
            in3 => \N__21676\,
            lcout => n4659,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i38_LC_12_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__21220\,
            in1 => \N__21564\,
            in2 => \N__21632\,
            in3 => \N__21607\,
            lcout => \c0.data_out_field_47_N_682_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__i9_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__21563\,
            in1 => \N__22221\,
            in2 => \_gnd_net_\,
            in3 => \N__21219\,
            lcout => data_out_field_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_378_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20985\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20946\,
            lcout => \c0.n1306\,
            ltout => \c0.n1306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_358_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22369\,
            in1 => \N__22355\,
            in2 => \N__22337\,
            in3 => \N__22334\,
            lcout => n4454,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_active_prev_611_LC_12_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22254\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx_active_prev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22955\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_343_LC_12_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22289\,
            in2 => \_gnd_net_\,
            in3 => \N__22252\,
            lcout => \c0.n50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22992\,
            in2 => \_gnd_net_\,
            in3 => \N__23072\,
            lcout => OPEN,
            ltout => \c0.tx.n2908_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_4_lut_LC_12_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__23161\,
            in1 => \N__22088\,
            in2 => \N__22277\,
            in3 => \N__23472\,
            lcout => OPEN,
            ltout => \c0.tx.n1457_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Active_47_LC_12_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011111010"
        )
    port map (
            in0 => \N__22253\,
            in1 => \_gnd_net_\,
            in2 => \N__22274\,
            in3 => \N__23162\,
            lcout => \c0.tx_active\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22955\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_288_LC_12_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22214\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22187\,
            lcout => n1325,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_3_lut_4_lut_LC_12_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__23471\,
            in1 => \N__23160\,
            in2 => \N__22481\,
            in3 => \N__22993\,
            lcout => n1025,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_adj_280_LC_12_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__22991\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22477\,
            lcout => \c0.tx.n752\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_adj_284_LC_12_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22471\,
            in2 => \_gnd_net_\,
            in3 => \N__23473\,
            lcout => \c0.tx.n3643\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_2_lut_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23574\,
            in2 => \_gnd_net_\,
            in3 => \N__23631\,
            lcout => \c0.tx.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i2_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000001000"
        )
    port map (
            in0 => \N__22604\,
            in1 => \N__23315\,
            in2 => \N__23100\,
            in3 => \N__23463\,
            lcout => \c0.tx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i2_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23080\,
            in1 => \N__23189\,
            in2 => \N__23493\,
            in3 => \N__23013\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i6_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000001000"
        )
    port map (
            in0 => \N__23558\,
            in1 => \N__23317\,
            in2 => \N__23102\,
            in3 => \N__23465\,
            lcout => \c0.tx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i4_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000001000"
        )
    port map (
            in0 => \N__23615\,
            in1 => \N__23316\,
            in2 => \N__23101\,
            in3 => \N__23464\,
            lcout => \c0.tx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_381_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22438\,
            in1 => \N__22390\,
            in2 => \_gnd_net_\,
            in3 => \N__22379\,
            lcout => \c0.n4477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i1_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__23309\,
            in1 => \N__22634\,
            in2 => \N__23099\,
            in3 => \N__23469\,
            lcout => \c0.tx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22956\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_adj_283_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__22593\,
            in1 => \N__23604\,
            in2 => \N__22625\,
            in3 => \N__22650\,
            lcout => OPEN,
            ltout => \c0.tx.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_adj_285_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__23522\,
            in1 => \N__22568\,
            in2 => \N__22562\,
            in3 => \N__23547\,
            lcout => \c0.tx.n17\,
            ltout => \c0.tx.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i7_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010001000"
        )
    port map (
            in0 => \N__23466\,
            in1 => \N__23531\,
            in2 => \N__22559\,
            in3 => \N__23314\,
            lcout => \c0.tx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22956\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i0_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__23308\,
            in1 => \N__22661\,
            in2 => \N__23098\,
            in3 => \N__23468\,
            lcout => \c0.tx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22956\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i5_LC_13_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000000"
        )
    port map (
            in0 => \N__23078\,
            in1 => \N__23313\,
            in2 => \N__23588\,
            in3 => \N__23470\,
            lcout => \c0.tx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22956\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i3_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101000"
        )
    port map (
            in0 => \N__22577\,
            in1 => \N__23467\,
            in2 => \N__23318\,
            in3 => \N__23079\,
            lcout => \c0.tx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22956\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_adj_281_LC_13_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23474\,
            in2 => \_gnd_net_\,
            in3 => \N__23070\,
            lcout => n4375,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i8_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011001000"
        )
    port map (
            in0 => \N__23475\,
            in1 => \N__23327\,
            in2 => \N__23307\,
            in3 => \N__23071\,
            lcout => \c0.tx.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22957\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_382_LC_13_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22556\,
            in1 => \N__22540\,
            in2 => \N__22529\,
            in3 => \N__22502\,
            lcout => n12_adj_944,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i1_LC_13_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__23002\,
            in1 => \N__23478\,
            in2 => \N__23200\,
            in3 => \N__23096\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22958\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i605_2_lut_LC_13_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23182\,
            in2 => \_gnd_net_\,
            in3 => \N__23000\,
            lcout => n88,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_LC_13_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011100000"
        )
    port map (
            in0 => \N__23172\,
            in1 => \N__23001\,
            in2 => \N__23264\,
            in3 => \N__23114\,
            lcout => OPEN,
            ltout => \n4_adj_946_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Done_44_LC_13_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011111100"
        )
    port map (
            in0 => \N__23263\,
            in1 => \N__23476\,
            in2 => \N__23321\,
            in3 => \N__23306\,
            lcout => tx_done,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22958\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i25_4_lut_LC_13_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__23245\,
            in1 => \N__23213\,
            in2 => \N__23193\,
            in3 => \N__23113\,
            lcout => OPEN,
            ltout => \c0.tx.n25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i0_LC_13_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__23003\,
            in1 => \N__23477\,
            in2 => \N__23105\,
            in3 => \N__23097\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22958\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_2_lut_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22673\,
            in1 => \N__22672\,
            in2 => \N__23479\,
            in3 => \N__22655\,
            lcout => \c0.tx.n1979\,
            ltout => OPEN,
            carryin => \bfn_14_27_0_\,
            carryout => \c0.tx.n3876\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_3_lut_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22652\,
            in1 => \N__22651\,
            in2 => \N__23483\,
            in3 => \N__22628\,
            lcout => \c0.tx.n1754\,
            ltout => OPEN,
            carryin => \c0.tx.n3876\,
            carryout => \c0.tx.n3877\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_4_lut_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22624\,
            in1 => \N__22623\,
            in2 => \N__23480\,
            in3 => \N__22598\,
            lcout => \c0.tx.n1751\,
            ltout => OPEN,
            carryin => \c0.tx.n3877\,
            carryout => \c0.tx.n3878\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_5_lut_LC_14_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22595\,
            in1 => \N__22594\,
            in2 => \N__23484\,
            in3 => \N__22571\,
            lcout => \c0.tx.n1748\,
            ltout => OPEN,
            carryin => \c0.tx.n3878\,
            carryout => \c0.tx.n3879\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_6_lut_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__23633\,
            in1 => \N__23632\,
            in2 => \N__23481\,
            in3 => \N__23609\,
            lcout => \c0.tx.n1745\,
            ltout => OPEN,
            carryin => \c0.tx.n3879\,
            carryout => \c0.tx.n3880\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_7_lut_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__23606\,
            in1 => \N__23605\,
            in2 => \N__23485\,
            in3 => \N__23579\,
            lcout => \c0.tx.n1742\,
            ltout => OPEN,
            carryin => \c0.tx.n3880\,
            carryout => \c0.tx.n3881\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_8_lut_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__23576\,
            in1 => \N__23575\,
            in2 => \N__23482\,
            in3 => \N__23552\,
            lcout => \c0.tx.n1739\,
            ltout => OPEN,
            carryin => \c0.tx.n3881\,
            carryout => \c0.tx.n3882\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_9_lut_LC_14_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__23549\,
            in1 => \N__23548\,
            in2 => \N__23486\,
            in3 => \N__23525\,
            lcout => \c0.tx.n1736\,
            ltout => OPEN,
            carryin => \c0.tx.n3882\,
            carryout => \c0.tx.n3883\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_10_lut_LC_14_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__23520\,
            in1 => \N__23521\,
            in2 => \N__23494\,
            in3 => \N__23330\,
            lcout => \c0.tx.n1733\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
