// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Sep 12 2019 19:18:20

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    output USBPU;
    input PIN_9;
    input PIN_8;
    input PIN_7;
    input PIN_6;
    input PIN_5;
    input PIN_4;
    inout PIN_3;
    input PIN_24;
    input PIN_23;
    input PIN_22;
    input PIN_21;
    input PIN_20;
    inout PIN_2;
    input PIN_19;
    input PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    input PIN_13;
    input PIN_12;
    input PIN_11;
    input PIN_10;
    inout PIN_1;
    output LED;
    input CLK;

    wire N__52613;
    wire N__52612;
    wire N__52611;
    wire N__52604;
    wire N__52603;
    wire N__52602;
    wire N__52595;
    wire N__52594;
    wire N__52593;
    wire N__52586;
    wire N__52585;
    wire N__52584;
    wire N__52577;
    wire N__52576;
    wire N__52575;
    wire N__52568;
    wire N__52567;
    wire N__52566;
    wire N__52549;
    wire N__52548;
    wire N__52545;
    wire N__52544;
    wire N__52541;
    wire N__52538;
    wire N__52535;
    wire N__52532;
    wire N__52527;
    wire N__52524;
    wire N__52521;
    wire N__52518;
    wire N__52513;
    wire N__52512;
    wire N__52511;
    wire N__52508;
    wire N__52505;
    wire N__52502;
    wire N__52499;
    wire N__52498;
    wire N__52497;
    wire N__52494;
    wire N__52491;
    wire N__52488;
    wire N__52483;
    wire N__52480;
    wire N__52477;
    wire N__52474;
    wire N__52465;
    wire N__52464;
    wire N__52463;
    wire N__52462;
    wire N__52461;
    wire N__52460;
    wire N__52459;
    wire N__52458;
    wire N__52457;
    wire N__52456;
    wire N__52455;
    wire N__52454;
    wire N__52453;
    wire N__52452;
    wire N__52451;
    wire N__52448;
    wire N__52445;
    wire N__52438;
    wire N__52437;
    wire N__52434;
    wire N__52429;
    wire N__52426;
    wire N__52419;
    wire N__52416;
    wire N__52415;
    wire N__52410;
    wire N__52409;
    wire N__52408;
    wire N__52407;
    wire N__52406;
    wire N__52405;
    wire N__52404;
    wire N__52399;
    wire N__52396;
    wire N__52393;
    wire N__52388;
    wire N__52385;
    wire N__52380;
    wire N__52377;
    wire N__52374;
    wire N__52369;
    wire N__52364;
    wire N__52361;
    wire N__52358;
    wire N__52355;
    wire N__52352;
    wire N__52351;
    wire N__52348;
    wire N__52345;
    wire N__52338;
    wire N__52335;
    wire N__52322;
    wire N__52319;
    wire N__52306;
    wire N__52303;
    wire N__52302;
    wire N__52301;
    wire N__52300;
    wire N__52297;
    wire N__52296;
    wire N__52295;
    wire N__52294;
    wire N__52291;
    wire N__52290;
    wire N__52289;
    wire N__52288;
    wire N__52285;
    wire N__52282;
    wire N__52279;
    wire N__52272;
    wire N__52269;
    wire N__52266;
    wire N__52265;
    wire N__52264;
    wire N__52261;
    wire N__52258;
    wire N__52257;
    wire N__52254;
    wire N__52251;
    wire N__52246;
    wire N__52243;
    wire N__52240;
    wire N__52237;
    wire N__52236;
    wire N__52233;
    wire N__52232;
    wire N__52231;
    wire N__52230;
    wire N__52227;
    wire N__52224;
    wire N__52221;
    wire N__52216;
    wire N__52213;
    wire N__52208;
    wire N__52205;
    wire N__52202;
    wire N__52197;
    wire N__52192;
    wire N__52187;
    wire N__52176;
    wire N__52175;
    wire N__52172;
    wire N__52165;
    wire N__52162;
    wire N__52159;
    wire N__52150;
    wire N__52147;
    wire N__52144;
    wire N__52141;
    wire N__52140;
    wire N__52137;
    wire N__52136;
    wire N__52135;
    wire N__52132;
    wire N__52131;
    wire N__52128;
    wire N__52125;
    wire N__52122;
    wire N__52119;
    wire N__52116;
    wire N__52113;
    wire N__52110;
    wire N__52099;
    wire N__52098;
    wire N__52097;
    wire N__52096;
    wire N__52093;
    wire N__52092;
    wire N__52091;
    wire N__52090;
    wire N__52089;
    wire N__52088;
    wire N__52087;
    wire N__52086;
    wire N__52085;
    wire N__52084;
    wire N__52083;
    wire N__52082;
    wire N__52081;
    wire N__52080;
    wire N__52077;
    wire N__52076;
    wire N__52073;
    wire N__52072;
    wire N__52071;
    wire N__52070;
    wire N__52067;
    wire N__52066;
    wire N__52065;
    wire N__52064;
    wire N__52063;
    wire N__52062;
    wire N__52061;
    wire N__52060;
    wire N__52057;
    wire N__52056;
    wire N__52055;
    wire N__52054;
    wire N__52045;
    wire N__52044;
    wire N__52043;
    wire N__52042;
    wire N__52041;
    wire N__52040;
    wire N__52039;
    wire N__52038;
    wire N__52035;
    wire N__52030;
    wire N__52025;
    wire N__52022;
    wire N__52019;
    wire N__52016;
    wire N__52013;
    wire N__52010;
    wire N__52005;
    wire N__51998;
    wire N__51997;
    wire N__51996;
    wire N__51995;
    wire N__51994;
    wire N__51993;
    wire N__51990;
    wire N__51987;
    wire N__51984;
    wire N__51979;
    wire N__51976;
    wire N__51973;
    wire N__51972;
    wire N__51971;
    wire N__51970;
    wire N__51967;
    wire N__51964;
    wire N__51957;
    wire N__51954;
    wire N__51951;
    wire N__51948;
    wire N__51939;
    wire N__51938;
    wire N__51935;
    wire N__51924;
    wire N__51921;
    wire N__51918;
    wire N__51913;
    wire N__51910;
    wire N__51905;
    wire N__51898;
    wire N__51893;
    wire N__51888;
    wire N__51887;
    wire N__51882;
    wire N__51879;
    wire N__51874;
    wire N__51871;
    wire N__51864;
    wire N__51857;
    wire N__51854;
    wire N__51851;
    wire N__51846;
    wire N__51843;
    wire N__51836;
    wire N__51829;
    wire N__51826;
    wire N__51823;
    wire N__51812;
    wire N__51809;
    wire N__51802;
    wire N__51797;
    wire N__51794;
    wire N__51781;
    wire N__51778;
    wire N__51775;
    wire N__51774;
    wire N__51771;
    wire N__51770;
    wire N__51767;
    wire N__51764;
    wire N__51763;
    wire N__51762;
    wire N__51761;
    wire N__51758;
    wire N__51755;
    wire N__51752;
    wire N__51749;
    wire N__51746;
    wire N__51743;
    wire N__51740;
    wire N__51739;
    wire N__51738;
    wire N__51733;
    wire N__51730;
    wire N__51727;
    wire N__51724;
    wire N__51721;
    wire N__51718;
    wire N__51715;
    wire N__51714;
    wire N__51711;
    wire N__51702;
    wire N__51701;
    wire N__51698;
    wire N__51695;
    wire N__51692;
    wire N__51689;
    wire N__51686;
    wire N__51683;
    wire N__51670;
    wire N__51667;
    wire N__51664;
    wire N__51661;
    wire N__51658;
    wire N__51655;
    wire N__51652;
    wire N__51651;
    wire N__51648;
    wire N__51647;
    wire N__51646;
    wire N__51645;
    wire N__51644;
    wire N__51643;
    wire N__51640;
    wire N__51637;
    wire N__51634;
    wire N__51633;
    wire N__51632;
    wire N__51631;
    wire N__51626;
    wire N__51623;
    wire N__51622;
    wire N__51621;
    wire N__51620;
    wire N__51619;
    wire N__51618;
    wire N__51617;
    wire N__51616;
    wire N__51615;
    wire N__51614;
    wire N__51613;
    wire N__51610;
    wire N__51609;
    wire N__51608;
    wire N__51601;
    wire N__51594;
    wire N__51589;
    wire N__51586;
    wire N__51583;
    wire N__51580;
    wire N__51577;
    wire N__51576;
    wire N__51571;
    wire N__51564;
    wire N__51561;
    wire N__51558;
    wire N__51553;
    wire N__51550;
    wire N__51545;
    wire N__51536;
    wire N__51535;
    wire N__51532;
    wire N__51525;
    wire N__51522;
    wire N__51515;
    wire N__51512;
    wire N__51509;
    wire N__51496;
    wire N__51493;
    wire N__51490;
    wire N__51487;
    wire N__51484;
    wire N__51481;
    wire N__51478;
    wire N__51475;
    wire N__51472;
    wire N__51469;
    wire N__51466;
    wire N__51463;
    wire N__51462;
    wire N__51459;
    wire N__51456;
    wire N__51453;
    wire N__51452;
    wire N__51451;
    wire N__51448;
    wire N__51447;
    wire N__51446;
    wire N__51443;
    wire N__51440;
    wire N__51437;
    wire N__51434;
    wire N__51431;
    wire N__51428;
    wire N__51423;
    wire N__51420;
    wire N__51415;
    wire N__51412;
    wire N__51411;
    wire N__51408;
    wire N__51405;
    wire N__51404;
    wire N__51401;
    wire N__51398;
    wire N__51395;
    wire N__51390;
    wire N__51387;
    wire N__51384;
    wire N__51381;
    wire N__51378;
    wire N__51373;
    wire N__51370;
    wire N__51365;
    wire N__51362;
    wire N__51359;
    wire N__51356;
    wire N__51353;
    wire N__51346;
    wire N__51343;
    wire N__51340;
    wire N__51339;
    wire N__51338;
    wire N__51335;
    wire N__51332;
    wire N__51329;
    wire N__51328;
    wire N__51327;
    wire N__51322;
    wire N__51319;
    wire N__51316;
    wire N__51313;
    wire N__51310;
    wire N__51305;
    wire N__51304;
    wire N__51301;
    wire N__51298;
    wire N__51295;
    wire N__51292;
    wire N__51289;
    wire N__51280;
    wire N__51279;
    wire N__51278;
    wire N__51277;
    wire N__51276;
    wire N__51275;
    wire N__51274;
    wire N__51273;
    wire N__51272;
    wire N__51271;
    wire N__51266;
    wire N__51261;
    wire N__51256;
    wire N__51251;
    wire N__51250;
    wire N__51249;
    wire N__51248;
    wire N__51247;
    wire N__51246;
    wire N__51245;
    wire N__51244;
    wire N__51243;
    wire N__51240;
    wire N__51237;
    wire N__51228;
    wire N__51225;
    wire N__51224;
    wire N__51223;
    wire N__51222;
    wire N__51221;
    wire N__51220;
    wire N__51219;
    wire N__51218;
    wire N__51217;
    wire N__51216;
    wire N__51215;
    wire N__51214;
    wire N__51213;
    wire N__51212;
    wire N__51211;
    wire N__51210;
    wire N__51209;
    wire N__51208;
    wire N__51207;
    wire N__51206;
    wire N__51205;
    wire N__51204;
    wire N__51203;
    wire N__51202;
    wire N__51201;
    wire N__51200;
    wire N__51199;
    wire N__51198;
    wire N__51197;
    wire N__51196;
    wire N__51195;
    wire N__51194;
    wire N__51193;
    wire N__51192;
    wire N__51191;
    wire N__51190;
    wire N__51189;
    wire N__51188;
    wire N__51187;
    wire N__51186;
    wire N__51185;
    wire N__51184;
    wire N__51183;
    wire N__51182;
    wire N__51181;
    wire N__51180;
    wire N__51179;
    wire N__51178;
    wire N__51177;
    wire N__51174;
    wire N__51171;
    wire N__51170;
    wire N__51169;
    wire N__51168;
    wire N__51165;
    wire N__51162;
    wire N__51161;
    wire N__51154;
    wire N__51151;
    wire N__51148;
    wire N__51147;
    wire N__51142;
    wire N__51139;
    wire N__51138;
    wire N__51137;
    wire N__51136;
    wire N__51135;
    wire N__51132;
    wire N__51131;
    wire N__51130;
    wire N__51129;
    wire N__51128;
    wire N__51127;
    wire N__51126;
    wire N__51117;
    wire N__51112;
    wire N__51109;
    wire N__51106;
    wire N__51105;
    wire N__51104;
    wire N__51103;
    wire N__51102;
    wire N__51097;
    wire N__51094;
    wire N__51089;
    wire N__51084;
    wire N__51081;
    wire N__51074;
    wire N__51073;
    wire N__51066;
    wire N__51061;
    wire N__51054;
    wire N__51043;
    wire N__51040;
    wire N__51033;
    wire N__51030;
    wire N__51027;
    wire N__51024;
    wire N__51021;
    wire N__51018;
    wire N__51015;
    wire N__51012;
    wire N__51005;
    wire N__51002;
    wire N__51001;
    wire N__50996;
    wire N__50995;
    wire N__50992;
    wire N__50989;
    wire N__50982;
    wire N__50977;
    wire N__50974;
    wire N__50971;
    wire N__50966;
    wire N__50965;
    wire N__50956;
    wire N__50953;
    wire N__50952;
    wire N__50951;
    wire N__50950;
    wire N__50949;
    wire N__50948;
    wire N__50947;
    wire N__50946;
    wire N__50945;
    wire N__50944;
    wire N__50943;
    wire N__50942;
    wire N__50941;
    wire N__50940;
    wire N__50939;
    wire N__50938;
    wire N__50937;
    wire N__50936;
    wire N__50935;
    wire N__50934;
    wire N__50933;
    wire N__50932;
    wire N__50931;
    wire N__50930;
    wire N__50929;
    wire N__50928;
    wire N__50927;
    wire N__50926;
    wire N__50925;
    wire N__50924;
    wire N__50923;
    wire N__50922;
    wire N__50921;
    wire N__50908;
    wire N__50901;
    wire N__50898;
    wire N__50889;
    wire N__50882;
    wire N__50879;
    wire N__50874;
    wire N__50871;
    wire N__50866;
    wire N__50863;
    wire N__50854;
    wire N__50849;
    wire N__50844;
    wire N__50841;
    wire N__50834;
    wire N__50831;
    wire N__50828;
    wire N__50825;
    wire N__50822;
    wire N__50819;
    wire N__50812;
    wire N__50807;
    wire N__50804;
    wire N__50799;
    wire N__50790;
    wire N__50775;
    wire N__50764;
    wire N__50753;
    wire N__50744;
    wire N__50737;
    wire N__50728;
    wire N__50721;
    wire N__50712;
    wire N__50703;
    wire N__50694;
    wire N__50689;
    wire N__50678;
    wire N__50673;
    wire N__50644;
    wire N__50641;
    wire N__50638;
    wire N__50637;
    wire N__50636;
    wire N__50635;
    wire N__50634;
    wire N__50631;
    wire N__50628;
    wire N__50623;
    wire N__50620;
    wire N__50617;
    wire N__50614;
    wire N__50611;
    wire N__50602;
    wire N__50601;
    wire N__50600;
    wire N__50599;
    wire N__50598;
    wire N__50597;
    wire N__50596;
    wire N__50595;
    wire N__50594;
    wire N__50593;
    wire N__50592;
    wire N__50591;
    wire N__50590;
    wire N__50589;
    wire N__50588;
    wire N__50587;
    wire N__50586;
    wire N__50585;
    wire N__50584;
    wire N__50583;
    wire N__50582;
    wire N__50581;
    wire N__50580;
    wire N__50579;
    wire N__50578;
    wire N__50577;
    wire N__50576;
    wire N__50575;
    wire N__50574;
    wire N__50573;
    wire N__50572;
    wire N__50571;
    wire N__50570;
    wire N__50569;
    wire N__50568;
    wire N__50567;
    wire N__50566;
    wire N__50565;
    wire N__50564;
    wire N__50563;
    wire N__50562;
    wire N__50561;
    wire N__50560;
    wire N__50559;
    wire N__50558;
    wire N__50557;
    wire N__50556;
    wire N__50555;
    wire N__50554;
    wire N__50553;
    wire N__50552;
    wire N__50551;
    wire N__50550;
    wire N__50549;
    wire N__50548;
    wire N__50547;
    wire N__50546;
    wire N__50545;
    wire N__50544;
    wire N__50543;
    wire N__50542;
    wire N__50541;
    wire N__50540;
    wire N__50539;
    wire N__50538;
    wire N__50537;
    wire N__50536;
    wire N__50535;
    wire N__50534;
    wire N__50533;
    wire N__50532;
    wire N__50531;
    wire N__50530;
    wire N__50529;
    wire N__50528;
    wire N__50527;
    wire N__50526;
    wire N__50525;
    wire N__50524;
    wire N__50523;
    wire N__50522;
    wire N__50521;
    wire N__50520;
    wire N__50519;
    wire N__50518;
    wire N__50517;
    wire N__50516;
    wire N__50515;
    wire N__50514;
    wire N__50513;
    wire N__50512;
    wire N__50511;
    wire N__50510;
    wire N__50509;
    wire N__50508;
    wire N__50507;
    wire N__50506;
    wire N__50505;
    wire N__50504;
    wire N__50503;
    wire N__50502;
    wire N__50501;
    wire N__50500;
    wire N__50499;
    wire N__50498;
    wire N__50497;
    wire N__50496;
    wire N__50495;
    wire N__50494;
    wire N__50493;
    wire N__50492;
    wire N__50491;
    wire N__50490;
    wire N__50489;
    wire N__50488;
    wire N__50487;
    wire N__50486;
    wire N__50485;
    wire N__50484;
    wire N__50483;
    wire N__50482;
    wire N__50481;
    wire N__50480;
    wire N__50479;
    wire N__50478;
    wire N__50477;
    wire N__50476;
    wire N__50475;
    wire N__50474;
    wire N__50473;
    wire N__50472;
    wire N__50471;
    wire N__50470;
    wire N__50469;
    wire N__50468;
    wire N__50467;
    wire N__50466;
    wire N__50465;
    wire N__50464;
    wire N__50463;
    wire N__50462;
    wire N__50461;
    wire N__50460;
    wire N__50459;
    wire N__50458;
    wire N__50457;
    wire N__50456;
    wire N__50455;
    wire N__50454;
    wire N__50453;
    wire N__50452;
    wire N__50451;
    wire N__50450;
    wire N__50449;
    wire N__50448;
    wire N__50447;
    wire N__50446;
    wire N__50445;
    wire N__50444;
    wire N__50443;
    wire N__50442;
    wire N__50441;
    wire N__50440;
    wire N__50439;
    wire N__50438;
    wire N__50437;
    wire N__50436;
    wire N__50435;
    wire N__50434;
    wire N__50433;
    wire N__50432;
    wire N__50431;
    wire N__50430;
    wire N__50429;
    wire N__50428;
    wire N__50427;
    wire N__50426;
    wire N__50425;
    wire N__50424;
    wire N__50423;
    wire N__50422;
    wire N__50421;
    wire N__50420;
    wire N__50419;
    wire N__50418;
    wire N__50417;
    wire N__50416;
    wire N__50415;
    wire N__50414;
    wire N__50413;
    wire N__50412;
    wire N__50411;
    wire N__50410;
    wire N__50409;
    wire N__50408;
    wire N__50407;
    wire N__50406;
    wire N__50405;
    wire N__50404;
    wire N__50403;
    wire N__50402;
    wire N__50401;
    wire N__50400;
    wire N__50399;
    wire N__50398;
    wire N__50397;
    wire N__50396;
    wire N__50395;
    wire N__50394;
    wire N__50393;
    wire N__50392;
    wire N__50391;
    wire N__50390;
    wire N__50389;
    wire N__50388;
    wire N__50387;
    wire N__50386;
    wire N__50385;
    wire N__50384;
    wire N__50383;
    wire N__50382;
    wire N__50381;
    wire N__50380;
    wire N__50379;
    wire N__50378;
    wire N__50377;
    wire N__49924;
    wire N__49921;
    wire N__49918;
    wire N__49917;
    wire N__49916;
    wire N__49913;
    wire N__49910;
    wire N__49907;
    wire N__49906;
    wire N__49901;
    wire N__49898;
    wire N__49897;
    wire N__49894;
    wire N__49891;
    wire N__49888;
    wire N__49885;
    wire N__49882;
    wire N__49879;
    wire N__49878;
    wire N__49873;
    wire N__49868;
    wire N__49865;
    wire N__49862;
    wire N__49855;
    wire N__49854;
    wire N__49851;
    wire N__49848;
    wire N__49847;
    wire N__49844;
    wire N__49843;
    wire N__49840;
    wire N__49837;
    wire N__49834;
    wire N__49831;
    wire N__49828;
    wire N__49825;
    wire N__49822;
    wire N__49813;
    wire N__49810;
    wire N__49809;
    wire N__49806;
    wire N__49803;
    wire N__49802;
    wire N__49801;
    wire N__49796;
    wire N__49793;
    wire N__49790;
    wire N__49785;
    wire N__49784;
    wire N__49781;
    wire N__49780;
    wire N__49777;
    wire N__49774;
    wire N__49771;
    wire N__49768;
    wire N__49763;
    wire N__49756;
    wire N__49755;
    wire N__49752;
    wire N__49749;
    wire N__49744;
    wire N__49743;
    wire N__49742;
    wire N__49739;
    wire N__49736;
    wire N__49735;
    wire N__49732;
    wire N__49729;
    wire N__49726;
    wire N__49723;
    wire N__49720;
    wire N__49717;
    wire N__49714;
    wire N__49707;
    wire N__49702;
    wire N__49699;
    wire N__49698;
    wire N__49695;
    wire N__49692;
    wire N__49687;
    wire N__49686;
    wire N__49685;
    wire N__49684;
    wire N__49681;
    wire N__49676;
    wire N__49673;
    wire N__49670;
    wire N__49663;
    wire N__49660;
    wire N__49659;
    wire N__49658;
    wire N__49655;
    wire N__49652;
    wire N__49651;
    wire N__49648;
    wire N__49643;
    wire N__49638;
    wire N__49633;
    wire N__49630;
    wire N__49629;
    wire N__49626;
    wire N__49623;
    wire N__49620;
    wire N__49617;
    wire N__49614;
    wire N__49611;
    wire N__49608;
    wire N__49603;
    wire N__49600;
    wire N__49597;
    wire N__49596;
    wire N__49595;
    wire N__49592;
    wire N__49589;
    wire N__49586;
    wire N__49583;
    wire N__49576;
    wire N__49573;
    wire N__49570;
    wire N__49567;
    wire N__49564;
    wire N__49561;
    wire N__49558;
    wire N__49557;
    wire N__49554;
    wire N__49551;
    wire N__49548;
    wire N__49545;
    wire N__49540;
    wire N__49537;
    wire N__49536;
    wire N__49535;
    wire N__49532;
    wire N__49529;
    wire N__49526;
    wire N__49525;
    wire N__49518;
    wire N__49515;
    wire N__49512;
    wire N__49507;
    wire N__49504;
    wire N__49503;
    wire N__49500;
    wire N__49497;
    wire N__49494;
    wire N__49491;
    wire N__49488;
    wire N__49485;
    wire N__49480;
    wire N__49477;
    wire N__49476;
    wire N__49473;
    wire N__49470;
    wire N__49469;
    wire N__49466;
    wire N__49463;
    wire N__49460;
    wire N__49459;
    wire N__49456;
    wire N__49453;
    wire N__49450;
    wire N__49447;
    wire N__49442;
    wire N__49439;
    wire N__49432;
    wire N__49431;
    wire N__49428;
    wire N__49427;
    wire N__49424;
    wire N__49423;
    wire N__49420;
    wire N__49417;
    wire N__49416;
    wire N__49415;
    wire N__49412;
    wire N__49409;
    wire N__49406;
    wire N__49403;
    wire N__49398;
    wire N__49393;
    wire N__49384;
    wire N__49381;
    wire N__49380;
    wire N__49379;
    wire N__49378;
    wire N__49375;
    wire N__49372;
    wire N__49369;
    wire N__49366;
    wire N__49365;
    wire N__49362;
    wire N__49357;
    wire N__49352;
    wire N__49345;
    wire N__49344;
    wire N__49343;
    wire N__49340;
    wire N__49337;
    wire N__49334;
    wire N__49331;
    wire N__49328;
    wire N__49325;
    wire N__49324;
    wire N__49323;
    wire N__49320;
    wire N__49317;
    wire N__49314;
    wire N__49309;
    wire N__49300;
    wire N__49297;
    wire N__49294;
    wire N__49291;
    wire N__49290;
    wire N__49287;
    wire N__49284;
    wire N__49283;
    wire N__49280;
    wire N__49277;
    wire N__49274;
    wire N__49273;
    wire N__49272;
    wire N__49271;
    wire N__49266;
    wire N__49263;
    wire N__49260;
    wire N__49257;
    wire N__49254;
    wire N__49251;
    wire N__49246;
    wire N__49237;
    wire N__49234;
    wire N__49231;
    wire N__49228;
    wire N__49227;
    wire N__49224;
    wire N__49221;
    wire N__49216;
    wire N__49213;
    wire N__49210;
    wire N__49207;
    wire N__49204;
    wire N__49201;
    wire N__49198;
    wire N__49195;
    wire N__49194;
    wire N__49191;
    wire N__49188;
    wire N__49187;
    wire N__49184;
    wire N__49183;
    wire N__49182;
    wire N__49179;
    wire N__49176;
    wire N__49173;
    wire N__49168;
    wire N__49165;
    wire N__49156;
    wire N__49153;
    wire N__49150;
    wire N__49147;
    wire N__49144;
    wire N__49141;
    wire N__49138;
    wire N__49135;
    wire N__49132;
    wire N__49129;
    wire N__49126;
    wire N__49123;
    wire N__49120;
    wire N__49117;
    wire N__49114;
    wire N__49111;
    wire N__49110;
    wire N__49107;
    wire N__49106;
    wire N__49103;
    wire N__49102;
    wire N__49099;
    wire N__49096;
    wire N__49095;
    wire N__49092;
    wire N__49089;
    wire N__49086;
    wire N__49083;
    wire N__49080;
    wire N__49077;
    wire N__49074;
    wire N__49073;
    wire N__49068;
    wire N__49065;
    wire N__49062;
    wire N__49059;
    wire N__49056;
    wire N__49051;
    wire N__49042;
    wire N__49039;
    wire N__49038;
    wire N__49035;
    wire N__49032;
    wire N__49029;
    wire N__49024;
    wire N__49021;
    wire N__49018;
    wire N__49015;
    wire N__49012;
    wire N__49011;
    wire N__49008;
    wire N__49007;
    wire N__49004;
    wire N__49003;
    wire N__49000;
    wire N__48997;
    wire N__48994;
    wire N__48993;
    wire N__48990;
    wire N__48989;
    wire N__48986;
    wire N__48981;
    wire N__48978;
    wire N__48975;
    wire N__48972;
    wire N__48969;
    wire N__48966;
    wire N__48955;
    wire N__48952;
    wire N__48949;
    wire N__48946;
    wire N__48943;
    wire N__48940;
    wire N__48937;
    wire N__48936;
    wire N__48935;
    wire N__48934;
    wire N__48931;
    wire N__48928;
    wire N__48925;
    wire N__48922;
    wire N__48919;
    wire N__48916;
    wire N__48913;
    wire N__48912;
    wire N__48909;
    wire N__48906;
    wire N__48903;
    wire N__48900;
    wire N__48897;
    wire N__48894;
    wire N__48883;
    wire N__48882;
    wire N__48877;
    wire N__48876;
    wire N__48873;
    wire N__48872;
    wire N__48869;
    wire N__48866;
    wire N__48865;
    wire N__48862;
    wire N__48859;
    wire N__48856;
    wire N__48853;
    wire N__48844;
    wire N__48841;
    wire N__48840;
    wire N__48839;
    wire N__48836;
    wire N__48833;
    wire N__48830;
    wire N__48829;
    wire N__48828;
    wire N__48825;
    wire N__48822;
    wire N__48819;
    wire N__48816;
    wire N__48815;
    wire N__48812;
    wire N__48809;
    wire N__48806;
    wire N__48803;
    wire N__48800;
    wire N__48797;
    wire N__48794;
    wire N__48781;
    wire N__48780;
    wire N__48777;
    wire N__48774;
    wire N__48769;
    wire N__48768;
    wire N__48767;
    wire N__48766;
    wire N__48763;
    wire N__48760;
    wire N__48757;
    wire N__48754;
    wire N__48751;
    wire N__48748;
    wire N__48745;
    wire N__48744;
    wire N__48741;
    wire N__48738;
    wire N__48733;
    wire N__48732;
    wire N__48729;
    wire N__48724;
    wire N__48721;
    wire N__48718;
    wire N__48715;
    wire N__48706;
    wire N__48705;
    wire N__48702;
    wire N__48701;
    wire N__48698;
    wire N__48695;
    wire N__48694;
    wire N__48691;
    wire N__48688;
    wire N__48685;
    wire N__48682;
    wire N__48679;
    wire N__48676;
    wire N__48667;
    wire N__48666;
    wire N__48665;
    wire N__48662;
    wire N__48659;
    wire N__48656;
    wire N__48655;
    wire N__48654;
    wire N__48653;
    wire N__48652;
    wire N__48651;
    wire N__48650;
    wire N__48649;
    wire N__48642;
    wire N__48641;
    wire N__48640;
    wire N__48639;
    wire N__48638;
    wire N__48637;
    wire N__48636;
    wire N__48631;
    wire N__48630;
    wire N__48629;
    wire N__48626;
    wire N__48625;
    wire N__48624;
    wire N__48623;
    wire N__48618;
    wire N__48615;
    wire N__48614;
    wire N__48611;
    wire N__48608;
    wire N__48605;
    wire N__48604;
    wire N__48601;
    wire N__48596;
    wire N__48595;
    wire N__48594;
    wire N__48593;
    wire N__48590;
    wire N__48587;
    wire N__48586;
    wire N__48585;
    wire N__48584;
    wire N__48583;
    wire N__48582;
    wire N__48581;
    wire N__48580;
    wire N__48579;
    wire N__48578;
    wire N__48575;
    wire N__48572;
    wire N__48569;
    wire N__48568;
    wire N__48565;
    wire N__48564;
    wire N__48561;
    wire N__48558;
    wire N__48555;
    wire N__48552;
    wire N__48549;
    wire N__48546;
    wire N__48543;
    wire N__48542;
    wire N__48541;
    wire N__48536;
    wire N__48535;
    wire N__48532;
    wire N__48527;
    wire N__48524;
    wire N__48517;
    wire N__48514;
    wire N__48513;
    wire N__48512;
    wire N__48509;
    wire N__48506;
    wire N__48503;
    wire N__48500;
    wire N__48497;
    wire N__48494;
    wire N__48493;
    wire N__48492;
    wire N__48491;
    wire N__48490;
    wire N__48489;
    wire N__48486;
    wire N__48481;
    wire N__48478;
    wire N__48475;
    wire N__48472;
    wire N__48469;
    wire N__48466;
    wire N__48465;
    wire N__48462;
    wire N__48461;
    wire N__48460;
    wire N__48459;
    wire N__48458;
    wire N__48457;
    wire N__48456;
    wire N__48453;
    wire N__48450;
    wire N__48447;
    wire N__48438;
    wire N__48433;
    wire N__48430;
    wire N__48427;
    wire N__48418;
    wire N__48415;
    wire N__48412;
    wire N__48409;
    wire N__48402;
    wire N__48397;
    wire N__48394;
    wire N__48393;
    wire N__48392;
    wire N__48391;
    wire N__48388;
    wire N__48381;
    wire N__48378;
    wire N__48375;
    wire N__48372;
    wire N__48365;
    wire N__48360;
    wire N__48355;
    wire N__48354;
    wire N__48353;
    wire N__48350;
    wire N__48341;
    wire N__48338;
    wire N__48331;
    wire N__48328;
    wire N__48323;
    wire N__48318;
    wire N__48315;
    wire N__48304;
    wire N__48299;
    wire N__48296;
    wire N__48279;
    wire N__48276;
    wire N__48273;
    wire N__48270;
    wire N__48265;
    wire N__48260;
    wire N__48251;
    wire N__48244;
    wire N__48229;
    wire N__48228;
    wire N__48227;
    wire N__48226;
    wire N__48225;
    wire N__48224;
    wire N__48223;
    wire N__48222;
    wire N__48221;
    wire N__48216;
    wire N__48215;
    wire N__48214;
    wire N__48213;
    wire N__48212;
    wire N__48211;
    wire N__48210;
    wire N__48209;
    wire N__48208;
    wire N__48207;
    wire N__48202;
    wire N__48195;
    wire N__48194;
    wire N__48191;
    wire N__48190;
    wire N__48189;
    wire N__48188;
    wire N__48187;
    wire N__48186;
    wire N__48183;
    wire N__48180;
    wire N__48177;
    wire N__48172;
    wire N__48171;
    wire N__48168;
    wire N__48167;
    wire N__48166;
    wire N__48165;
    wire N__48164;
    wire N__48161;
    wire N__48154;
    wire N__48151;
    wire N__48146;
    wire N__48143;
    wire N__48142;
    wire N__48141;
    wire N__48140;
    wire N__48137;
    wire N__48134;
    wire N__48131;
    wire N__48128;
    wire N__48125;
    wire N__48122;
    wire N__48121;
    wire N__48120;
    wire N__48111;
    wire N__48108;
    wire N__48107;
    wire N__48106;
    wire N__48105;
    wire N__48104;
    wire N__48101;
    wire N__48098;
    wire N__48097;
    wire N__48096;
    wire N__48093;
    wire N__48092;
    wire N__48089;
    wire N__48086;
    wire N__48081;
    wire N__48074;
    wire N__48067;
    wire N__48066;
    wire N__48065;
    wire N__48060;
    wire N__48053;
    wire N__48052;
    wire N__48051;
    wire N__48048;
    wire N__48045;
    wire N__48044;
    wire N__48043;
    wire N__48042;
    wire N__48039;
    wire N__48034;
    wire N__48031;
    wire N__48030;
    wire N__48027;
    wire N__48024;
    wire N__48021;
    wire N__48016;
    wire N__48013;
    wire N__48010;
    wire N__48009;
    wire N__48006;
    wire N__48003;
    wire N__47998;
    wire N__47991;
    wire N__47988;
    wire N__47985;
    wire N__47980;
    wire N__47977;
    wire N__47974;
    wire N__47969;
    wire N__47964;
    wire N__47963;
    wire N__47962;
    wire N__47961;
    wire N__47960;
    wire N__47957;
    wire N__47954;
    wire N__47949;
    wire N__47946;
    wire N__47943;
    wire N__47938;
    wire N__47933;
    wire N__47930;
    wire N__47927;
    wire N__47924;
    wire N__47917;
    wire N__47910;
    wire N__47901;
    wire N__47898;
    wire N__47895;
    wire N__47890;
    wire N__47881;
    wire N__47874;
    wire N__47865;
    wire N__47860;
    wire N__47855;
    wire N__47848;
    wire N__47839;
    wire N__47836;
    wire N__47833;
    wire N__47830;
    wire N__47827;
    wire N__47824;
    wire N__47821;
    wire N__47818;
    wire N__47817;
    wire N__47816;
    wire N__47815;
    wire N__47814;
    wire N__47811;
    wire N__47808;
    wire N__47805;
    wire N__47804;
    wire N__47801;
    wire N__47798;
    wire N__47791;
    wire N__47788;
    wire N__47787;
    wire N__47784;
    wire N__47781;
    wire N__47776;
    wire N__47773;
    wire N__47770;
    wire N__47767;
    wire N__47762;
    wire N__47761;
    wire N__47758;
    wire N__47755;
    wire N__47752;
    wire N__47749;
    wire N__47740;
    wire N__47737;
    wire N__47734;
    wire N__47731;
    wire N__47728;
    wire N__47725;
    wire N__47722;
    wire N__47719;
    wire N__47716;
    wire N__47715;
    wire N__47714;
    wire N__47713;
    wire N__47712;
    wire N__47711;
    wire N__47710;
    wire N__47709;
    wire N__47708;
    wire N__47707;
    wire N__47706;
    wire N__47705;
    wire N__47702;
    wire N__47699;
    wire N__47696;
    wire N__47693;
    wire N__47690;
    wire N__47687;
    wire N__47684;
    wire N__47681;
    wire N__47678;
    wire N__47675;
    wire N__47674;
    wire N__47671;
    wire N__47668;
    wire N__47661;
    wire N__47660;
    wire N__47659;
    wire N__47658;
    wire N__47651;
    wire N__47646;
    wire N__47645;
    wire N__47644;
    wire N__47643;
    wire N__47642;
    wire N__47639;
    wire N__47636;
    wire N__47633;
    wire N__47632;
    wire N__47631;
    wire N__47624;
    wire N__47621;
    wire N__47618;
    wire N__47615;
    wire N__47612;
    wire N__47609;
    wire N__47606;
    wire N__47601;
    wire N__47598;
    wire N__47595;
    wire N__47590;
    wire N__47587;
    wire N__47584;
    wire N__47579;
    wire N__47578;
    wire N__47569;
    wire N__47560;
    wire N__47557;
    wire N__47550;
    wire N__47547;
    wire N__47536;
    wire N__47533;
    wire N__47530;
    wire N__47527;
    wire N__47524;
    wire N__47521;
    wire N__47518;
    wire N__47515;
    wire N__47512;
    wire N__47509;
    wire N__47506;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47488;
    wire N__47485;
    wire N__47484;
    wire N__47481;
    wire N__47478;
    wire N__47475;
    wire N__47472;
    wire N__47467;
    wire N__47464;
    wire N__47461;
    wire N__47458;
    wire N__47455;
    wire N__47452;
    wire N__47451;
    wire N__47448;
    wire N__47445;
    wire N__47440;
    wire N__47437;
    wire N__47434;
    wire N__47431;
    wire N__47428;
    wire N__47425;
    wire N__47422;
    wire N__47419;
    wire N__47416;
    wire N__47415;
    wire N__47412;
    wire N__47411;
    wire N__47410;
    wire N__47409;
    wire N__47406;
    wire N__47403;
    wire N__47398;
    wire N__47395;
    wire N__47392;
    wire N__47389;
    wire N__47386;
    wire N__47377;
    wire N__47376;
    wire N__47373;
    wire N__47372;
    wire N__47371;
    wire N__47368;
    wire N__47365;
    wire N__47362;
    wire N__47361;
    wire N__47360;
    wire N__47357;
    wire N__47354;
    wire N__47351;
    wire N__47348;
    wire N__47345;
    wire N__47342;
    wire N__47339;
    wire N__47332;
    wire N__47329;
    wire N__47320;
    wire N__47317;
    wire N__47314;
    wire N__47313;
    wire N__47312;
    wire N__47309;
    wire N__47306;
    wire N__47303;
    wire N__47302;
    wire N__47301;
    wire N__47296;
    wire N__47293;
    wire N__47290;
    wire N__47287;
    wire N__47282;
    wire N__47279;
    wire N__47276;
    wire N__47271;
    wire N__47270;
    wire N__47267;
    wire N__47264;
    wire N__47261;
    wire N__47258;
    wire N__47255;
    wire N__47248;
    wire N__47247;
    wire N__47244;
    wire N__47241;
    wire N__47238;
    wire N__47237;
    wire N__47232;
    wire N__47231;
    wire N__47228;
    wire N__47225;
    wire N__47224;
    wire N__47221;
    wire N__47216;
    wire N__47213;
    wire N__47210;
    wire N__47203;
    wire N__47200;
    wire N__47199;
    wire N__47198;
    wire N__47195;
    wire N__47192;
    wire N__47189;
    wire N__47188;
    wire N__47185;
    wire N__47182;
    wire N__47181;
    wire N__47178;
    wire N__47175;
    wire N__47172;
    wire N__47169;
    wire N__47166;
    wire N__47163;
    wire N__47152;
    wire N__47149;
    wire N__47146;
    wire N__47143;
    wire N__47140;
    wire N__47139;
    wire N__47138;
    wire N__47135;
    wire N__47132;
    wire N__47129;
    wire N__47126;
    wire N__47123;
    wire N__47120;
    wire N__47117;
    wire N__47112;
    wire N__47109;
    wire N__47106;
    wire N__47101;
    wire N__47098;
    wire N__47097;
    wire N__47096;
    wire N__47093;
    wire N__47090;
    wire N__47087;
    wire N__47084;
    wire N__47081;
    wire N__47078;
    wire N__47075;
    wire N__47072;
    wire N__47069;
    wire N__47064;
    wire N__47061;
    wire N__47056;
    wire N__47053;
    wire N__47050;
    wire N__47049;
    wire N__47046;
    wire N__47045;
    wire N__47042;
    wire N__47039;
    wire N__47034;
    wire N__47029;
    wire N__47026;
    wire N__47023;
    wire N__47022;
    wire N__47019;
    wire N__47016;
    wire N__47011;
    wire N__47008;
    wire N__47005;
    wire N__47004;
    wire N__47001;
    wire N__46998;
    wire N__46993;
    wire N__46990;
    wire N__46987;
    wire N__46984;
    wire N__46981;
    wire N__46978;
    wire N__46975;
    wire N__46972;
    wire N__46969;
    wire N__46968;
    wire N__46967;
    wire N__46966;
    wire N__46963;
    wire N__46960;
    wire N__46955;
    wire N__46952;
    wire N__46949;
    wire N__46946;
    wire N__46943;
    wire N__46940;
    wire N__46937;
    wire N__46934;
    wire N__46927;
    wire N__46926;
    wire N__46921;
    wire N__46918;
    wire N__46915;
    wire N__46912;
    wire N__46911;
    wire N__46908;
    wire N__46905;
    wire N__46902;
    wire N__46899;
    wire N__46898;
    wire N__46895;
    wire N__46892;
    wire N__46889;
    wire N__46882;
    wire N__46879;
    wire N__46878;
    wire N__46875;
    wire N__46872;
    wire N__46867;
    wire N__46864;
    wire N__46863;
    wire N__46860;
    wire N__46857;
    wire N__46856;
    wire N__46855;
    wire N__46854;
    wire N__46853;
    wire N__46848;
    wire N__46845;
    wire N__46842;
    wire N__46839;
    wire N__46836;
    wire N__46831;
    wire N__46822;
    wire N__46821;
    wire N__46820;
    wire N__46817;
    wire N__46812;
    wire N__46809;
    wire N__46804;
    wire N__46803;
    wire N__46800;
    wire N__46799;
    wire N__46798;
    wire N__46795;
    wire N__46792;
    wire N__46791;
    wire N__46788;
    wire N__46785;
    wire N__46780;
    wire N__46777;
    wire N__46772;
    wire N__46769;
    wire N__46766;
    wire N__46763;
    wire N__46756;
    wire N__46755;
    wire N__46752;
    wire N__46749;
    wire N__46746;
    wire N__46743;
    wire N__46740;
    wire N__46739;
    wire N__46734;
    wire N__46731;
    wire N__46726;
    wire N__46723;
    wire N__46720;
    wire N__46719;
    wire N__46716;
    wire N__46713;
    wire N__46710;
    wire N__46707;
    wire N__46702;
    wire N__46701;
    wire N__46698;
    wire N__46697;
    wire N__46694;
    wire N__46691;
    wire N__46690;
    wire N__46689;
    wire N__46686;
    wire N__46683;
    wire N__46680;
    wire N__46677;
    wire N__46674;
    wire N__46671;
    wire N__46664;
    wire N__46661;
    wire N__46654;
    wire N__46651;
    wire N__46648;
    wire N__46647;
    wire N__46646;
    wire N__46643;
    wire N__46640;
    wire N__46637;
    wire N__46630;
    wire N__46627;
    wire N__46624;
    wire N__46623;
    wire N__46622;
    wire N__46621;
    wire N__46620;
    wire N__46617;
    wire N__46616;
    wire N__46613;
    wire N__46610;
    wire N__46607;
    wire N__46606;
    wire N__46603;
    wire N__46600;
    wire N__46597;
    wire N__46590;
    wire N__46589;
    wire N__46586;
    wire N__46583;
    wire N__46580;
    wire N__46577;
    wire N__46574;
    wire N__46571;
    wire N__46568;
    wire N__46567;
    wire N__46564;
    wire N__46555;
    wire N__46552;
    wire N__46549;
    wire N__46546;
    wire N__46543;
    wire N__46540;
    wire N__46537;
    wire N__46534;
    wire N__46531;
    wire N__46526;
    wire N__46519;
    wire N__46518;
    wire N__46515;
    wire N__46512;
    wire N__46509;
    wire N__46506;
    wire N__46501;
    wire N__46498;
    wire N__46495;
    wire N__46492;
    wire N__46491;
    wire N__46490;
    wire N__46489;
    wire N__46488;
    wire N__46487;
    wire N__46486;
    wire N__46485;
    wire N__46482;
    wire N__46481;
    wire N__46480;
    wire N__46479;
    wire N__46476;
    wire N__46475;
    wire N__46472;
    wire N__46467;
    wire N__46466;
    wire N__46459;
    wire N__46456;
    wire N__46453;
    wire N__46450;
    wire N__46449;
    wire N__46448;
    wire N__46447;
    wire N__46444;
    wire N__46441;
    wire N__46438;
    wire N__46437;
    wire N__46436;
    wire N__46435;
    wire N__46434;
    wire N__46433;
    wire N__46432;
    wire N__46427;
    wire N__46424;
    wire N__46423;
    wire N__46422;
    wire N__46421;
    wire N__46420;
    wire N__46419;
    wire N__46418;
    wire N__46417;
    wire N__46416;
    wire N__46415;
    wire N__46408;
    wire N__46405;
    wire N__46404;
    wire N__46403;
    wire N__46402;
    wire N__46401;
    wire N__46400;
    wire N__46399;
    wire N__46396;
    wire N__46395;
    wire N__46390;
    wire N__46383;
    wire N__46380;
    wire N__46369;
    wire N__46366;
    wire N__46363;
    wire N__46362;
    wire N__46359;
    wire N__46356;
    wire N__46353;
    wire N__46344;
    wire N__46339;
    wire N__46336;
    wire N__46333;
    wire N__46322;
    wire N__46321;
    wire N__46318;
    wire N__46315;
    wire N__46312;
    wire N__46307;
    wire N__46306;
    wire N__46305;
    wire N__46304;
    wire N__46303;
    wire N__46302;
    wire N__46301;
    wire N__46300;
    wire N__46299;
    wire N__46298;
    wire N__46293;
    wire N__46288;
    wire N__46285;
    wire N__46268;
    wire N__46263;
    wire N__46256;
    wire N__46253;
    wire N__46242;
    wire N__46235;
    wire N__46232;
    wire N__46227;
    wire N__46224;
    wire N__46221;
    wire N__46218;
    wire N__46201;
    wire N__46200;
    wire N__46199;
    wire N__46196;
    wire N__46193;
    wire N__46192;
    wire N__46189;
    wire N__46186;
    wire N__46183;
    wire N__46180;
    wire N__46177;
    wire N__46174;
    wire N__46171;
    wire N__46166;
    wire N__46163;
    wire N__46160;
    wire N__46155;
    wire N__46150;
    wire N__46149;
    wire N__46146;
    wire N__46143;
    wire N__46140;
    wire N__46139;
    wire N__46138;
    wire N__46137;
    wire N__46134;
    wire N__46133;
    wire N__46132;
    wire N__46131;
    wire N__46130;
    wire N__46129;
    wire N__46128;
    wire N__46125;
    wire N__46122;
    wire N__46119;
    wire N__46116;
    wire N__46113;
    wire N__46110;
    wire N__46107;
    wire N__46106;
    wire N__46103;
    wire N__46100;
    wire N__46097;
    wire N__46094;
    wire N__46089;
    wire N__46086;
    wire N__46083;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46071;
    wire N__46066;
    wire N__46063;
    wire N__46058;
    wire N__46051;
    wire N__46048;
    wire N__46041;
    wire N__46036;
    wire N__46033;
    wire N__46024;
    wire N__46021;
    wire N__46018;
    wire N__46017;
    wire N__46014;
    wire N__46011;
    wire N__46008;
    wire N__46005;
    wire N__46000;
    wire N__45999;
    wire N__45998;
    wire N__45997;
    wire N__45996;
    wire N__45995;
    wire N__45994;
    wire N__45993;
    wire N__45992;
    wire N__45991;
    wire N__45990;
    wire N__45989;
    wire N__45988;
    wire N__45987;
    wire N__45986;
    wire N__45983;
    wire N__45982;
    wire N__45979;
    wire N__45978;
    wire N__45977;
    wire N__45976;
    wire N__45971;
    wire N__45968;
    wire N__45957;
    wire N__45956;
    wire N__45955;
    wire N__45954;
    wire N__45953;
    wire N__45952;
    wire N__45951;
    wire N__45948;
    wire N__45947;
    wire N__45944;
    wire N__45943;
    wire N__45940;
    wire N__45937;
    wire N__45936;
    wire N__45935;
    wire N__45932;
    wire N__45931;
    wire N__45930;
    wire N__45929;
    wire N__45928;
    wire N__45925;
    wire N__45924;
    wire N__45921;
    wire N__45920;
    wire N__45915;
    wire N__45912;
    wire N__45911;
    wire N__45908;
    wire N__45907;
    wire N__45906;
    wire N__45905;
    wire N__45898;
    wire N__45889;
    wire N__45886;
    wire N__45883;
    wire N__45880;
    wire N__45879;
    wire N__45876;
    wire N__45875;
    wire N__45874;
    wire N__45869;
    wire N__45864;
    wire N__45861;
    wire N__45858;
    wire N__45855;
    wire N__45852;
    wire N__45849;
    wire N__45848;
    wire N__45845;
    wire N__45844;
    wire N__45841;
    wire N__45838;
    wire N__45835;
    wire N__45830;
    wire N__45825;
    wire N__45820;
    wire N__45817;
    wire N__45812;
    wire N__45807;
    wire N__45804;
    wire N__45803;
    wire N__45802;
    wire N__45801;
    wire N__45798;
    wire N__45795;
    wire N__45792;
    wire N__45789;
    wire N__45786;
    wire N__45785;
    wire N__45784;
    wire N__45783;
    wire N__45782;
    wire N__45781;
    wire N__45778;
    wire N__45771;
    wire N__45762;
    wire N__45761;
    wire N__45760;
    wire N__45757;
    wire N__45754;
    wire N__45751;
    wire N__45748;
    wire N__45745;
    wire N__45742;
    wire N__45739;
    wire N__45734;
    wire N__45725;
    wire N__45718;
    wire N__45713;
    wire N__45706;
    wire N__45695;
    wire N__45688;
    wire N__45683;
    wire N__45680;
    wire N__45667;
    wire N__45662;
    wire N__45651;
    wire N__45640;
    wire N__45637;
    wire N__45634;
    wire N__45631;
    wire N__45628;
    wire N__45625;
    wire N__45624;
    wire N__45621;
    wire N__45618;
    wire N__45617;
    wire N__45616;
    wire N__45613;
    wire N__45606;
    wire N__45601;
    wire N__45598;
    wire N__45597;
    wire N__45596;
    wire N__45593;
    wire N__45590;
    wire N__45587;
    wire N__45582;
    wire N__45577;
    wire N__45574;
    wire N__45571;
    wire N__45568;
    wire N__45565;
    wire N__45562;
    wire N__45559;
    wire N__45556;
    wire N__45553;
    wire N__45550;
    wire N__45549;
    wire N__45548;
    wire N__45547;
    wire N__45546;
    wire N__45545;
    wire N__45544;
    wire N__45541;
    wire N__45538;
    wire N__45537;
    wire N__45536;
    wire N__45533;
    wire N__45526;
    wire N__45523;
    wire N__45520;
    wire N__45517;
    wire N__45516;
    wire N__45515;
    wire N__45514;
    wire N__45511;
    wire N__45510;
    wire N__45507;
    wire N__45504;
    wire N__45499;
    wire N__45496;
    wire N__45493;
    wire N__45492;
    wire N__45491;
    wire N__45488;
    wire N__45487;
    wire N__45486;
    wire N__45483;
    wire N__45480;
    wire N__45477;
    wire N__45474;
    wire N__45471;
    wire N__45462;
    wire N__45457;
    wire N__45456;
    wire N__45455;
    wire N__45454;
    wire N__45451;
    wire N__45446;
    wire N__45443;
    wire N__45436;
    wire N__45435;
    wire N__45428;
    wire N__45425;
    wire N__45422;
    wire N__45419;
    wire N__45416;
    wire N__45411;
    wire N__45408;
    wire N__45405;
    wire N__45402;
    wire N__45399;
    wire N__45382;
    wire N__45379;
    wire N__45378;
    wire N__45375;
    wire N__45372;
    wire N__45367;
    wire N__45364;
    wire N__45363;
    wire N__45362;
    wire N__45361;
    wire N__45358;
    wire N__45355;
    wire N__45352;
    wire N__45349;
    wire N__45348;
    wire N__45343;
    wire N__45340;
    wire N__45337;
    wire N__45336;
    wire N__45333;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45310;
    wire N__45301;
    wire N__45300;
    wire N__45297;
    wire N__45294;
    wire N__45293;
    wire N__45292;
    wire N__45289;
    wire N__45286;
    wire N__45283;
    wire N__45280;
    wire N__45279;
    wire N__45272;
    wire N__45269;
    wire N__45266;
    wire N__45261;
    wire N__45256;
    wire N__45253;
    wire N__45252;
    wire N__45249;
    wire N__45248;
    wire N__45245;
    wire N__45242;
    wire N__45239;
    wire N__45238;
    wire N__45235;
    wire N__45230;
    wire N__45227;
    wire N__45224;
    wire N__45221;
    wire N__45214;
    wire N__45213;
    wire N__45210;
    wire N__45207;
    wire N__45206;
    wire N__45205;
    wire N__45202;
    wire N__45201;
    wire N__45198;
    wire N__45195;
    wire N__45192;
    wire N__45191;
    wire N__45188;
    wire N__45185;
    wire N__45182;
    wire N__45177;
    wire N__45174;
    wire N__45169;
    wire N__45166;
    wire N__45161;
    wire N__45158;
    wire N__45151;
    wire N__45148;
    wire N__45145;
    wire N__45144;
    wire N__45141;
    wire N__45138;
    wire N__45133;
    wire N__45130;
    wire N__45127;
    wire N__45124;
    wire N__45121;
    wire N__45118;
    wire N__45115;
    wire N__45114;
    wire N__45111;
    wire N__45108;
    wire N__45107;
    wire N__45106;
    wire N__45103;
    wire N__45100;
    wire N__45099;
    wire N__45094;
    wire N__45089;
    wire N__45086;
    wire N__45079;
    wire N__45076;
    wire N__45075;
    wire N__45074;
    wire N__45071;
    wire N__45070;
    wire N__45069;
    wire N__45064;
    wire N__45061;
    wire N__45058;
    wire N__45057;
    wire N__45054;
    wire N__45051;
    wire N__45046;
    wire N__45043;
    wire N__45034;
    wire N__45031;
    wire N__45028;
    wire N__45025;
    wire N__45022;
    wire N__45021;
    wire N__45020;
    wire N__45017;
    wire N__45012;
    wire N__45009;
    wire N__45004;
    wire N__45001;
    wire N__45000;
    wire N__44997;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44985;
    wire N__44982;
    wire N__44977;
    wire N__44974;
    wire N__44973;
    wire N__44970;
    wire N__44967;
    wire N__44964;
    wire N__44961;
    wire N__44958;
    wire N__44955;
    wire N__44950;
    wire N__44947;
    wire N__44946;
    wire N__44945;
    wire N__44944;
    wire N__44943;
    wire N__44940;
    wire N__44937;
    wire N__44934;
    wire N__44931;
    wire N__44928;
    wire N__44925;
    wire N__44922;
    wire N__44919;
    wire N__44918;
    wire N__44915;
    wire N__44912;
    wire N__44907;
    wire N__44904;
    wire N__44901;
    wire N__44896;
    wire N__44887;
    wire N__44886;
    wire N__44883;
    wire N__44882;
    wire N__44879;
    wire N__44878;
    wire N__44877;
    wire N__44874;
    wire N__44871;
    wire N__44868;
    wire N__44863;
    wire N__44854;
    wire N__44853;
    wire N__44852;
    wire N__44849;
    wire N__44846;
    wire N__44843;
    wire N__44842;
    wire N__44841;
    wire N__44838;
    wire N__44835;
    wire N__44832;
    wire N__44829;
    wire N__44826;
    wire N__44823;
    wire N__44820;
    wire N__44817;
    wire N__44806;
    wire N__44803;
    wire N__44800;
    wire N__44797;
    wire N__44794;
    wire N__44791;
    wire N__44788;
    wire N__44785;
    wire N__44784;
    wire N__44783;
    wire N__44782;
    wire N__44779;
    wire N__44776;
    wire N__44773;
    wire N__44770;
    wire N__44765;
    wire N__44762;
    wire N__44761;
    wire N__44758;
    wire N__44755;
    wire N__44752;
    wire N__44749;
    wire N__44746;
    wire N__44737;
    wire N__44736;
    wire N__44735;
    wire N__44734;
    wire N__44731;
    wire N__44728;
    wire N__44723;
    wire N__44720;
    wire N__44717;
    wire N__44716;
    wire N__44713;
    wire N__44708;
    wire N__44705;
    wire N__44700;
    wire N__44695;
    wire N__44694;
    wire N__44691;
    wire N__44688;
    wire N__44687;
    wire N__44686;
    wire N__44683;
    wire N__44680;
    wire N__44677;
    wire N__44674;
    wire N__44667;
    wire N__44666;
    wire N__44663;
    wire N__44660;
    wire N__44657;
    wire N__44654;
    wire N__44647;
    wire N__44646;
    wire N__44643;
    wire N__44642;
    wire N__44639;
    wire N__44636;
    wire N__44633;
    wire N__44632;
    wire N__44629;
    wire N__44626;
    wire N__44621;
    wire N__44614;
    wire N__44611;
    wire N__44610;
    wire N__44607;
    wire N__44606;
    wire N__44605;
    wire N__44602;
    wire N__44599;
    wire N__44596;
    wire N__44593;
    wire N__44584;
    wire N__44581;
    wire N__44578;
    wire N__44575;
    wire N__44572;
    wire N__44569;
    wire N__44568;
    wire N__44567;
    wire N__44566;
    wire N__44563;
    wire N__44558;
    wire N__44557;
    wire N__44554;
    wire N__44551;
    wire N__44548;
    wire N__44547;
    wire N__44544;
    wire N__44541;
    wire N__44538;
    wire N__44535;
    wire N__44532;
    wire N__44527;
    wire N__44518;
    wire N__44515;
    wire N__44512;
    wire N__44509;
    wire N__44506;
    wire N__44503;
    wire N__44500;
    wire N__44497;
    wire N__44494;
    wire N__44491;
    wire N__44488;
    wire N__44487;
    wire N__44484;
    wire N__44481;
    wire N__44480;
    wire N__44477;
    wire N__44474;
    wire N__44471;
    wire N__44470;
    wire N__44463;
    wire N__44462;
    wire N__44459;
    wire N__44456;
    wire N__44453;
    wire N__44450;
    wire N__44443;
    wire N__44442;
    wire N__44441;
    wire N__44438;
    wire N__44435;
    wire N__44434;
    wire N__44431;
    wire N__44428;
    wire N__44425;
    wire N__44422;
    wire N__44421;
    wire N__44418;
    wire N__44411;
    wire N__44408;
    wire N__44405;
    wire N__44402;
    wire N__44395;
    wire N__44394;
    wire N__44393;
    wire N__44390;
    wire N__44385;
    wire N__44382;
    wire N__44379;
    wire N__44378;
    wire N__44375;
    wire N__44372;
    wire N__44369;
    wire N__44366;
    wire N__44363;
    wire N__44356;
    wire N__44355;
    wire N__44354;
    wire N__44351;
    wire N__44348;
    wire N__44347;
    wire N__44346;
    wire N__44345;
    wire N__44342;
    wire N__44339;
    wire N__44336;
    wire N__44333;
    wire N__44328;
    wire N__44323;
    wire N__44320;
    wire N__44315;
    wire N__44308;
    wire N__44307;
    wire N__44304;
    wire N__44301;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44289;
    wire N__44284;
    wire N__44283;
    wire N__44282;
    wire N__44279;
    wire N__44276;
    wire N__44273;
    wire N__44272;
    wire N__44269;
    wire N__44266;
    wire N__44263;
    wire N__44260;
    wire N__44257;
    wire N__44254;
    wire N__44251;
    wire N__44242;
    wire N__44241;
    wire N__44238;
    wire N__44235;
    wire N__44232;
    wire N__44231;
    wire N__44230;
    wire N__44225;
    wire N__44222;
    wire N__44221;
    wire N__44218;
    wire N__44215;
    wire N__44212;
    wire N__44209;
    wire N__44200;
    wire N__44197;
    wire N__44196;
    wire N__44195;
    wire N__44192;
    wire N__44189;
    wire N__44186;
    wire N__44183;
    wire N__44180;
    wire N__44173;
    wire N__44172;
    wire N__44169;
    wire N__44166;
    wire N__44165;
    wire N__44164;
    wire N__44161;
    wire N__44160;
    wire N__44157;
    wire N__44154;
    wire N__44151;
    wire N__44148;
    wire N__44145;
    wire N__44140;
    wire N__44139;
    wire N__44136;
    wire N__44133;
    wire N__44130;
    wire N__44127;
    wire N__44124;
    wire N__44121;
    wire N__44110;
    wire N__44107;
    wire N__44106;
    wire N__44103;
    wire N__44100;
    wire N__44097;
    wire N__44092;
    wire N__44091;
    wire N__44090;
    wire N__44087;
    wire N__44082;
    wire N__44081;
    wire N__44078;
    wire N__44075;
    wire N__44072;
    wire N__44069;
    wire N__44068;
    wire N__44065;
    wire N__44062;
    wire N__44059;
    wire N__44056;
    wire N__44051;
    wire N__44044;
    wire N__44041;
    wire N__44040;
    wire N__44039;
    wire N__44038;
    wire N__44035;
    wire N__44032;
    wire N__44029;
    wire N__44026;
    wire N__44019;
    wire N__44014;
    wire N__44013;
    wire N__44012;
    wire N__44009;
    wire N__44006;
    wire N__44003;
    wire N__44002;
    wire N__43997;
    wire N__43994;
    wire N__43991;
    wire N__43990;
    wire N__43987;
    wire N__43984;
    wire N__43981;
    wire N__43978;
    wire N__43973;
    wire N__43970;
    wire N__43963;
    wire N__43960;
    wire N__43959;
    wire N__43958;
    wire N__43955;
    wire N__43952;
    wire N__43949;
    wire N__43948;
    wire N__43947;
    wire N__43944;
    wire N__43941;
    wire N__43938;
    wire N__43935;
    wire N__43932;
    wire N__43929;
    wire N__43924;
    wire N__43915;
    wire N__43912;
    wire N__43909;
    wire N__43908;
    wire N__43907;
    wire N__43906;
    wire N__43903;
    wire N__43902;
    wire N__43899;
    wire N__43896;
    wire N__43891;
    wire N__43888;
    wire N__43885;
    wire N__43884;
    wire N__43881;
    wire N__43878;
    wire N__43873;
    wire N__43870;
    wire N__43867;
    wire N__43864;
    wire N__43861;
    wire N__43852;
    wire N__43849;
    wire N__43848;
    wire N__43847;
    wire N__43844;
    wire N__43841;
    wire N__43838;
    wire N__43833;
    wire N__43832;
    wire N__43831;
    wire N__43828;
    wire N__43825;
    wire N__43822;
    wire N__43819;
    wire N__43816;
    wire N__43811;
    wire N__43804;
    wire N__43801;
    wire N__43798;
    wire N__43795;
    wire N__43792;
    wire N__43789;
    wire N__43786;
    wire N__43783;
    wire N__43780;
    wire N__43777;
    wire N__43774;
    wire N__43771;
    wire N__43768;
    wire N__43767;
    wire N__43766;
    wire N__43763;
    wire N__43760;
    wire N__43757;
    wire N__43756;
    wire N__43753;
    wire N__43750;
    wire N__43747;
    wire N__43744;
    wire N__43739;
    wire N__43732;
    wire N__43729;
    wire N__43728;
    wire N__43725;
    wire N__43724;
    wire N__43721;
    wire N__43718;
    wire N__43715;
    wire N__43712;
    wire N__43709;
    wire N__43704;
    wire N__43699;
    wire N__43696;
    wire N__43693;
    wire N__43690;
    wire N__43687;
    wire N__43686;
    wire N__43683;
    wire N__43682;
    wire N__43679;
    wire N__43678;
    wire N__43675;
    wire N__43672;
    wire N__43669;
    wire N__43666;
    wire N__43663;
    wire N__43658;
    wire N__43651;
    wire N__43648;
    wire N__43647;
    wire N__43646;
    wire N__43643;
    wire N__43640;
    wire N__43637;
    wire N__43636;
    wire N__43633;
    wire N__43630;
    wire N__43627;
    wire N__43626;
    wire N__43623;
    wire N__43620;
    wire N__43617;
    wire N__43614;
    wire N__43611;
    wire N__43600;
    wire N__43597;
    wire N__43594;
    wire N__43591;
    wire N__43588;
    wire N__43585;
    wire N__43584;
    wire N__43581;
    wire N__43578;
    wire N__43575;
    wire N__43574;
    wire N__43573;
    wire N__43572;
    wire N__43569;
    wire N__43566;
    wire N__43563;
    wire N__43560;
    wire N__43557;
    wire N__43554;
    wire N__43549;
    wire N__43546;
    wire N__43537;
    wire N__43534;
    wire N__43531;
    wire N__43528;
    wire N__43525;
    wire N__43524;
    wire N__43523;
    wire N__43520;
    wire N__43519;
    wire N__43516;
    wire N__43513;
    wire N__43510;
    wire N__43507;
    wire N__43504;
    wire N__43501;
    wire N__43498;
    wire N__43489;
    wire N__43486;
    wire N__43483;
    wire N__43480;
    wire N__43477;
    wire N__43474;
    wire N__43473;
    wire N__43472;
    wire N__43469;
    wire N__43466;
    wire N__43465;
    wire N__43464;
    wire N__43463;
    wire N__43460;
    wire N__43457;
    wire N__43454;
    wire N__43451;
    wire N__43448;
    wire N__43445;
    wire N__43438;
    wire N__43433;
    wire N__43430;
    wire N__43427;
    wire N__43424;
    wire N__43417;
    wire N__43414;
    wire N__43411;
    wire N__43410;
    wire N__43407;
    wire N__43404;
    wire N__43401;
    wire N__43398;
    wire N__43395;
    wire N__43392;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43380;
    wire N__43377;
    wire N__43374;
    wire N__43373;
    wire N__43372;
    wire N__43369;
    wire N__43366;
    wire N__43363;
    wire N__43360;
    wire N__43357;
    wire N__43354;
    wire N__43351;
    wire N__43346;
    wire N__43341;
    wire N__43336;
    wire N__43335;
    wire N__43332;
    wire N__43329;
    wire N__43324;
    wire N__43321;
    wire N__43318;
    wire N__43315;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43305;
    wire N__43304;
    wire N__43301;
    wire N__43300;
    wire N__43297;
    wire N__43294;
    wire N__43291;
    wire N__43286;
    wire N__43279;
    wire N__43278;
    wire N__43277;
    wire N__43274;
    wire N__43271;
    wire N__43268;
    wire N__43267;
    wire N__43266;
    wire N__43263;
    wire N__43258;
    wire N__43255;
    wire N__43252;
    wire N__43247;
    wire N__43244;
    wire N__43237;
    wire N__43234;
    wire N__43231;
    wire N__43228;
    wire N__43227;
    wire N__43224;
    wire N__43221;
    wire N__43216;
    wire N__43215;
    wire N__43212;
    wire N__43209;
    wire N__43204;
    wire N__43201;
    wire N__43198;
    wire N__43195;
    wire N__43192;
    wire N__43189;
    wire N__43186;
    wire N__43183;
    wire N__43182;
    wire N__43179;
    wire N__43176;
    wire N__43171;
    wire N__43168;
    wire N__43165;
    wire N__43162;
    wire N__43159;
    wire N__43156;
    wire N__43153;
    wire N__43152;
    wire N__43151;
    wire N__43150;
    wire N__43149;
    wire N__43148;
    wire N__43147;
    wire N__43146;
    wire N__43143;
    wire N__43140;
    wire N__43139;
    wire N__43136;
    wire N__43133;
    wire N__43130;
    wire N__43127;
    wire N__43124;
    wire N__43121;
    wire N__43120;
    wire N__43119;
    wire N__43116;
    wire N__43113;
    wire N__43112;
    wire N__43109;
    wire N__43106;
    wire N__43103;
    wire N__43096;
    wire N__43093;
    wire N__43090;
    wire N__43087;
    wire N__43082;
    wire N__43079;
    wire N__43078;
    wire N__43075;
    wire N__43072;
    wire N__43069;
    wire N__43064;
    wire N__43055;
    wire N__43052;
    wire N__43039;
    wire N__43036;
    wire N__43033;
    wire N__43030;
    wire N__43027;
    wire N__43024;
    wire N__43021;
    wire N__43020;
    wire N__43017;
    wire N__43014;
    wire N__43013;
    wire N__43012;
    wire N__43011;
    wire N__43008;
    wire N__43005;
    wire N__43002;
    wire N__42999;
    wire N__42996;
    wire N__42989;
    wire N__42982;
    wire N__42981;
    wire N__42978;
    wire N__42975;
    wire N__42972;
    wire N__42969;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42958;
    wire N__42957;
    wire N__42954;
    wire N__42949;
    wire N__42944;
    wire N__42937;
    wire N__42936;
    wire N__42933;
    wire N__42930;
    wire N__42927;
    wire N__42922;
    wire N__42921;
    wire N__42918;
    wire N__42915;
    wire N__42910;
    wire N__42909;
    wire N__42906;
    wire N__42903;
    wire N__42898;
    wire N__42895;
    wire N__42892;
    wire N__42889;
    wire N__42886;
    wire N__42883;
    wire N__42882;
    wire N__42879;
    wire N__42876;
    wire N__42873;
    wire N__42870;
    wire N__42865;
    wire N__42864;
    wire N__42863;
    wire N__42862;
    wire N__42861;
    wire N__42860;
    wire N__42855;
    wire N__42852;
    wire N__42851;
    wire N__42848;
    wire N__42847;
    wire N__42844;
    wire N__42843;
    wire N__42842;
    wire N__42839;
    wire N__42838;
    wire N__42835;
    wire N__42832;
    wire N__42829;
    wire N__42826;
    wire N__42823;
    wire N__42822;
    wire N__42817;
    wire N__42812;
    wire N__42809;
    wire N__42804;
    wire N__42799;
    wire N__42798;
    wire N__42795;
    wire N__42792;
    wire N__42781;
    wire N__42778;
    wire N__42775;
    wire N__42770;
    wire N__42763;
    wire N__42762;
    wire N__42761;
    wire N__42760;
    wire N__42759;
    wire N__42758;
    wire N__42755;
    wire N__42754;
    wire N__42753;
    wire N__42752;
    wire N__42751;
    wire N__42750;
    wire N__42749;
    wire N__42746;
    wire N__42745;
    wire N__42742;
    wire N__42739;
    wire N__42736;
    wire N__42733;
    wire N__42728;
    wire N__42727;
    wire N__42726;
    wire N__42725;
    wire N__42722;
    wire N__42719;
    wire N__42716;
    wire N__42713;
    wire N__42712;
    wire N__42711;
    wire N__42710;
    wire N__42709;
    wire N__42708;
    wire N__42705;
    wire N__42702;
    wire N__42701;
    wire N__42698;
    wire N__42695;
    wire N__42692;
    wire N__42687;
    wire N__42684;
    wire N__42681;
    wire N__42680;
    wire N__42675;
    wire N__42670;
    wire N__42661;
    wire N__42660;
    wire N__42657;
    wire N__42654;
    wire N__42653;
    wire N__42652;
    wire N__42649;
    wire N__42648;
    wire N__42647;
    wire N__42646;
    wire N__42645;
    wire N__42644;
    wire N__42641;
    wire N__42638;
    wire N__42635;
    wire N__42624;
    wire N__42623;
    wire N__42622;
    wire N__42619;
    wire N__42616;
    wire N__42611;
    wire N__42608;
    wire N__42607;
    wire N__42604;
    wire N__42603;
    wire N__42598;
    wire N__42593;
    wire N__42592;
    wire N__42589;
    wire N__42584;
    wire N__42581;
    wire N__42580;
    wire N__42577;
    wire N__42576;
    wire N__42575;
    wire N__42574;
    wire N__42571;
    wire N__42568;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42546;
    wire N__42543;
    wire N__42538;
    wire N__42533;
    wire N__42530;
    wire N__42525;
    wire N__42522;
    wire N__42515;
    wire N__42510;
    wire N__42503;
    wire N__42498;
    wire N__42495;
    wire N__42484;
    wire N__42469;
    wire N__42468;
    wire N__42467;
    wire N__42466;
    wire N__42465;
    wire N__42464;
    wire N__42461;
    wire N__42458;
    wire N__42455;
    wire N__42452;
    wire N__42449;
    wire N__42446;
    wire N__42443;
    wire N__42440;
    wire N__42439;
    wire N__42436;
    wire N__42431;
    wire N__42428;
    wire N__42425;
    wire N__42422;
    wire N__42419;
    wire N__42414;
    wire N__42403;
    wire N__42402;
    wire N__42401;
    wire N__42400;
    wire N__42397;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42383;
    wire N__42380;
    wire N__42375;
    wire N__42372;
    wire N__42371;
    wire N__42368;
    wire N__42365;
    wire N__42362;
    wire N__42357;
    wire N__42354;
    wire N__42349;
    wire N__42340;
    wire N__42337;
    wire N__42334;
    wire N__42331;
    wire N__42328;
    wire N__42327;
    wire N__42326;
    wire N__42323;
    wire N__42320;
    wire N__42317;
    wire N__42316;
    wire N__42315;
    wire N__42310;
    wire N__42307;
    wire N__42302;
    wire N__42299;
    wire N__42296;
    wire N__42289;
    wire N__42288;
    wire N__42285;
    wire N__42284;
    wire N__42281;
    wire N__42278;
    wire N__42275;
    wire N__42270;
    wire N__42267;
    wire N__42264;
    wire N__42259;
    wire N__42256;
    wire N__42253;
    wire N__42250;
    wire N__42249;
    wire N__42246;
    wire N__42243;
    wire N__42238;
    wire N__42235;
    wire N__42232;
    wire N__42229;
    wire N__42228;
    wire N__42225;
    wire N__42222;
    wire N__42217;
    wire N__42214;
    wire N__42211;
    wire N__42208;
    wire N__42205;
    wire N__42204;
    wire N__42203;
    wire N__42202;
    wire N__42199;
    wire N__42194;
    wire N__42191;
    wire N__42188;
    wire N__42185;
    wire N__42180;
    wire N__42177;
    wire N__42172;
    wire N__42171;
    wire N__42166;
    wire N__42163;
    wire N__42160;
    wire N__42157;
    wire N__42156;
    wire N__42155;
    wire N__42152;
    wire N__42149;
    wire N__42146;
    wire N__42141;
    wire N__42138;
    wire N__42135;
    wire N__42132;
    wire N__42131;
    wire N__42126;
    wire N__42123;
    wire N__42118;
    wire N__42115;
    wire N__42112;
    wire N__42109;
    wire N__42106;
    wire N__42103;
    wire N__42100;
    wire N__42097;
    wire N__42094;
    wire N__42091;
    wire N__42088;
    wire N__42085;
    wire N__42082;
    wire N__42079;
    wire N__42076;
    wire N__42073;
    wire N__42072;
    wire N__42069;
    wire N__42068;
    wire N__42067;
    wire N__42066;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42051;
    wire N__42048;
    wire N__42043;
    wire N__42034;
    wire N__42033;
    wire N__42028;
    wire N__42025;
    wire N__42024;
    wire N__42023;
    wire N__42020;
    wire N__42015;
    wire N__42010;
    wire N__42007;
    wire N__42004;
    wire N__42001;
    wire N__41998;
    wire N__41995;
    wire N__41994;
    wire N__41991;
    wire N__41988;
    wire N__41985;
    wire N__41982;
    wire N__41979;
    wire N__41974;
    wire N__41971;
    wire N__41968;
    wire N__41965;
    wire N__41962;
    wire N__41959;
    wire N__41958;
    wire N__41957;
    wire N__41956;
    wire N__41953;
    wire N__41950;
    wire N__41945;
    wire N__41938;
    wire N__41935;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41923;
    wire N__41920;
    wire N__41917;
    wire N__41914;
    wire N__41911;
    wire N__41908;
    wire N__41905;
    wire N__41902;
    wire N__41899;
    wire N__41896;
    wire N__41893;
    wire N__41890;
    wire N__41889;
    wire N__41886;
    wire N__41883;
    wire N__41878;
    wire N__41875;
    wire N__41872;
    wire N__41869;
    wire N__41868;
    wire N__41867;
    wire N__41866;
    wire N__41863;
    wire N__41860;
    wire N__41859;
    wire N__41856;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41844;
    wire N__41833;
    wire N__41832;
    wire N__41831;
    wire N__41828;
    wire N__41825;
    wire N__41822;
    wire N__41819;
    wire N__41816;
    wire N__41815;
    wire N__41812;
    wire N__41809;
    wire N__41806;
    wire N__41803;
    wire N__41800;
    wire N__41795;
    wire N__41788;
    wire N__41785;
    wire N__41782;
    wire N__41779;
    wire N__41776;
    wire N__41773;
    wire N__41770;
    wire N__41767;
    wire N__41764;
    wire N__41761;
    wire N__41758;
    wire N__41755;
    wire N__41754;
    wire N__41753;
    wire N__41752;
    wire N__41749;
    wire N__41746;
    wire N__41743;
    wire N__41740;
    wire N__41737;
    wire N__41734;
    wire N__41733;
    wire N__41730;
    wire N__41727;
    wire N__41724;
    wire N__41721;
    wire N__41718;
    wire N__41713;
    wire N__41704;
    wire N__41703;
    wire N__41700;
    wire N__41697;
    wire N__41696;
    wire N__41691;
    wire N__41690;
    wire N__41689;
    wire N__41686;
    wire N__41683;
    wire N__41680;
    wire N__41677;
    wire N__41668;
    wire N__41665;
    wire N__41662;
    wire N__41659;
    wire N__41656;
    wire N__41653;
    wire N__41650;
    wire N__41647;
    wire N__41646;
    wire N__41641;
    wire N__41638;
    wire N__41635;
    wire N__41632;
    wire N__41629;
    wire N__41626;
    wire N__41623;
    wire N__41620;
    wire N__41617;
    wire N__41614;
    wire N__41611;
    wire N__41608;
    wire N__41605;
    wire N__41602;
    wire N__41599;
    wire N__41596;
    wire N__41595;
    wire N__41594;
    wire N__41591;
    wire N__41588;
    wire N__41585;
    wire N__41582;
    wire N__41579;
    wire N__41576;
    wire N__41571;
    wire N__41570;
    wire N__41569;
    wire N__41566;
    wire N__41563;
    wire N__41558;
    wire N__41551;
    wire N__41548;
    wire N__41545;
    wire N__41542;
    wire N__41539;
    wire N__41536;
    wire N__41535;
    wire N__41534;
    wire N__41531;
    wire N__41526;
    wire N__41521;
    wire N__41518;
    wire N__41515;
    wire N__41514;
    wire N__41513;
    wire N__41510;
    wire N__41509;
    wire N__41506;
    wire N__41503;
    wire N__41500;
    wire N__41497;
    wire N__41488;
    wire N__41487;
    wire N__41484;
    wire N__41481;
    wire N__41476;
    wire N__41473;
    wire N__41470;
    wire N__41469;
    wire N__41466;
    wire N__41465;
    wire N__41464;
    wire N__41461;
    wire N__41458;
    wire N__41455;
    wire N__41454;
    wire N__41451;
    wire N__41448;
    wire N__41445;
    wire N__41444;
    wire N__41441;
    wire N__41438;
    wire N__41433;
    wire N__41430;
    wire N__41427;
    wire N__41424;
    wire N__41413;
    wire N__41410;
    wire N__41407;
    wire N__41406;
    wire N__41403;
    wire N__41400;
    wire N__41399;
    wire N__41398;
    wire N__41395;
    wire N__41392;
    wire N__41387;
    wire N__41380;
    wire N__41379;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41367;
    wire N__41364;
    wire N__41359;
    wire N__41356;
    wire N__41353;
    wire N__41350;
    wire N__41347;
    wire N__41346;
    wire N__41345;
    wire N__41344;
    wire N__41343;
    wire N__41340;
    wire N__41337;
    wire N__41334;
    wire N__41331;
    wire N__41328;
    wire N__41325;
    wire N__41322;
    wire N__41319;
    wire N__41318;
    wire N__41313;
    wire N__41308;
    wire N__41305;
    wire N__41302;
    wire N__41297;
    wire N__41294;
    wire N__41287;
    wire N__41284;
    wire N__41281;
    wire N__41278;
    wire N__41275;
    wire N__41272;
    wire N__41269;
    wire N__41268;
    wire N__41265;
    wire N__41264;
    wire N__41263;
    wire N__41260;
    wire N__41255;
    wire N__41252;
    wire N__41249;
    wire N__41242;
    wire N__41239;
    wire N__41238;
    wire N__41235;
    wire N__41232;
    wire N__41229;
    wire N__41226;
    wire N__41221;
    wire N__41218;
    wire N__41217;
    wire N__41214;
    wire N__41211;
    wire N__41208;
    wire N__41205;
    wire N__41204;
    wire N__41203;
    wire N__41198;
    wire N__41195;
    wire N__41192;
    wire N__41189;
    wire N__41186;
    wire N__41185;
    wire N__41182;
    wire N__41179;
    wire N__41176;
    wire N__41173;
    wire N__41170;
    wire N__41161;
    wire N__41160;
    wire N__41159;
    wire N__41158;
    wire N__41155;
    wire N__41150;
    wire N__41147;
    wire N__41140;
    wire N__41137;
    wire N__41136;
    wire N__41135;
    wire N__41132;
    wire N__41131;
    wire N__41128;
    wire N__41125;
    wire N__41122;
    wire N__41119;
    wire N__41110;
    wire N__41109;
    wire N__41106;
    wire N__41103;
    wire N__41100;
    wire N__41097;
    wire N__41094;
    wire N__41091;
    wire N__41086;
    wire N__41083;
    wire N__41080;
    wire N__41077;
    wire N__41074;
    wire N__41071;
    wire N__41068;
    wire N__41067;
    wire N__41064;
    wire N__41061;
    wire N__41058;
    wire N__41055;
    wire N__41050;
    wire N__41049;
    wire N__41046;
    wire N__41043;
    wire N__41042;
    wire N__41041;
    wire N__41040;
    wire N__41037;
    wire N__41034;
    wire N__41031;
    wire N__41026;
    wire N__41017;
    wire N__41014;
    wire N__41011;
    wire N__41008;
    wire N__41005;
    wire N__41002;
    wire N__40999;
    wire N__40996;
    wire N__40993;
    wire N__40990;
    wire N__40987;
    wire N__40984;
    wire N__40983;
    wire N__40980;
    wire N__40979;
    wire N__40978;
    wire N__40977;
    wire N__40974;
    wire N__40971;
    wire N__40968;
    wire N__40965;
    wire N__40962;
    wire N__40957;
    wire N__40954;
    wire N__40949;
    wire N__40942;
    wire N__40939;
    wire N__40936;
    wire N__40933;
    wire N__40930;
    wire N__40927;
    wire N__40924;
    wire N__40921;
    wire N__40918;
    wire N__40915;
    wire N__40912;
    wire N__40909;
    wire N__40906;
    wire N__40905;
    wire N__40904;
    wire N__40901;
    wire N__40900;
    wire N__40895;
    wire N__40892;
    wire N__40889;
    wire N__40886;
    wire N__40879;
    wire N__40876;
    wire N__40875;
    wire N__40872;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40862;
    wire N__40861;
    wire N__40860;
    wire N__40857;
    wire N__40852;
    wire N__40849;
    wire N__40846;
    wire N__40843;
    wire N__40840;
    wire N__40835;
    wire N__40828;
    wire N__40825;
    wire N__40822;
    wire N__40819;
    wire N__40816;
    wire N__40813;
    wire N__40810;
    wire N__40807;
    wire N__40804;
    wire N__40803;
    wire N__40800;
    wire N__40799;
    wire N__40796;
    wire N__40793;
    wire N__40790;
    wire N__40783;
    wire N__40782;
    wire N__40781;
    wire N__40778;
    wire N__40775;
    wire N__40774;
    wire N__40771;
    wire N__40768;
    wire N__40765;
    wire N__40762;
    wire N__40753;
    wire N__40750;
    wire N__40747;
    wire N__40744;
    wire N__40741;
    wire N__40738;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40726;
    wire N__40725;
    wire N__40724;
    wire N__40721;
    wire N__40718;
    wire N__40717;
    wire N__40714;
    wire N__40711;
    wire N__40708;
    wire N__40705;
    wire N__40696;
    wire N__40693;
    wire N__40692;
    wire N__40689;
    wire N__40686;
    wire N__40683;
    wire N__40680;
    wire N__40677;
    wire N__40674;
    wire N__40669;
    wire N__40668;
    wire N__40665;
    wire N__40662;
    wire N__40659;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40641;
    wire N__40638;
    wire N__40635;
    wire N__40634;
    wire N__40631;
    wire N__40628;
    wire N__40625;
    wire N__40620;
    wire N__40619;
    wire N__40618;
    wire N__40615;
    wire N__40612;
    wire N__40609;
    wire N__40606;
    wire N__40603;
    wire N__40594;
    wire N__40591;
    wire N__40588;
    wire N__40585;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40573;
    wire N__40570;
    wire N__40569;
    wire N__40566;
    wire N__40563;
    wire N__40560;
    wire N__40557;
    wire N__40552;
    wire N__40551;
    wire N__40550;
    wire N__40547;
    wire N__40544;
    wire N__40541;
    wire N__40536;
    wire N__40533;
    wire N__40530;
    wire N__40525;
    wire N__40524;
    wire N__40521;
    wire N__40518;
    wire N__40515;
    wire N__40512;
    wire N__40509;
    wire N__40508;
    wire N__40505;
    wire N__40504;
    wire N__40501;
    wire N__40498;
    wire N__40495;
    wire N__40492;
    wire N__40487;
    wire N__40480;
    wire N__40479;
    wire N__40478;
    wire N__40475;
    wire N__40474;
    wire N__40471;
    wire N__40468;
    wire N__40465;
    wire N__40462;
    wire N__40459;
    wire N__40456;
    wire N__40455;
    wire N__40454;
    wire N__40449;
    wire N__40444;
    wire N__40439;
    wire N__40436;
    wire N__40429;
    wire N__40426;
    wire N__40425;
    wire N__40420;
    wire N__40417;
    wire N__40414;
    wire N__40413;
    wire N__40412;
    wire N__40409;
    wire N__40408;
    wire N__40405;
    wire N__40402;
    wire N__40399;
    wire N__40396;
    wire N__40393;
    wire N__40386;
    wire N__40385;
    wire N__40384;
    wire N__40381;
    wire N__40378;
    wire N__40373;
    wire N__40366;
    wire N__40363;
    wire N__40360;
    wire N__40357;
    wire N__40354;
    wire N__40351;
    wire N__40348;
    wire N__40345;
    wire N__40342;
    wire N__40341;
    wire N__40340;
    wire N__40337;
    wire N__40336;
    wire N__40335;
    wire N__40332;
    wire N__40329;
    wire N__40326;
    wire N__40323;
    wire N__40322;
    wire N__40319;
    wire N__40316;
    wire N__40313;
    wire N__40308;
    wire N__40305;
    wire N__40294;
    wire N__40291;
    wire N__40290;
    wire N__40287;
    wire N__40284;
    wire N__40281;
    wire N__40278;
    wire N__40273;
    wire N__40270;
    wire N__40269;
    wire N__40266;
    wire N__40263;
    wire N__40260;
    wire N__40259;
    wire N__40254;
    wire N__40251;
    wire N__40248;
    wire N__40243;
    wire N__40242;
    wire N__40241;
    wire N__40238;
    wire N__40235;
    wire N__40232;
    wire N__40229;
    wire N__40228;
    wire N__40223;
    wire N__40220;
    wire N__40219;
    wire N__40216;
    wire N__40211;
    wire N__40208;
    wire N__40205;
    wire N__40202;
    wire N__40195;
    wire N__40192;
    wire N__40189;
    wire N__40188;
    wire N__40187;
    wire N__40184;
    wire N__40181;
    wire N__40178;
    wire N__40175;
    wire N__40170;
    wire N__40167;
    wire N__40162;
    wire N__40159;
    wire N__40156;
    wire N__40153;
    wire N__40152;
    wire N__40149;
    wire N__40148;
    wire N__40147;
    wire N__40146;
    wire N__40143;
    wire N__40140;
    wire N__40137;
    wire N__40132;
    wire N__40129;
    wire N__40126;
    wire N__40121;
    wire N__40118;
    wire N__40115;
    wire N__40112;
    wire N__40105;
    wire N__40104;
    wire N__40101;
    wire N__40098;
    wire N__40095;
    wire N__40092;
    wire N__40087;
    wire N__40084;
    wire N__40081;
    wire N__40080;
    wire N__40079;
    wire N__40078;
    wire N__40077;
    wire N__40074;
    wire N__40067;
    wire N__40064;
    wire N__40057;
    wire N__40056;
    wire N__40053;
    wire N__40050;
    wire N__40045;
    wire N__40044;
    wire N__40041;
    wire N__40038;
    wire N__40035;
    wire N__40032;
    wire N__40027;
    wire N__40026;
    wire N__40025;
    wire N__40024;
    wire N__40023;
    wire N__40018;
    wire N__40013;
    wire N__40010;
    wire N__40005;
    wire N__40000;
    wire N__39997;
    wire N__39994;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39984;
    wire N__39981;
    wire N__39976;
    wire N__39973;
    wire N__39970;
    wire N__39967;
    wire N__39964;
    wire N__39961;
    wire N__39958;
    wire N__39957;
    wire N__39954;
    wire N__39951;
    wire N__39948;
    wire N__39945;
    wire N__39942;
    wire N__39939;
    wire N__39934;
    wire N__39933;
    wire N__39932;
    wire N__39929;
    wire N__39924;
    wire N__39919;
    wire N__39916;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39903;
    wire N__39900;
    wire N__39899;
    wire N__39898;
    wire N__39895;
    wire N__39892;
    wire N__39887;
    wire N__39884;
    wire N__39877;
    wire N__39876;
    wire N__39875;
    wire N__39872;
    wire N__39871;
    wire N__39868;
    wire N__39865;
    wire N__39862;
    wire N__39859;
    wire N__39858;
    wire N__39851;
    wire N__39848;
    wire N__39845;
    wire N__39838;
    wire N__39837;
    wire N__39834;
    wire N__39833;
    wire N__39832;
    wire N__39827;
    wire N__39822;
    wire N__39817;
    wire N__39814;
    wire N__39813;
    wire N__39812;
    wire N__39809;
    wire N__39806;
    wire N__39803;
    wire N__39800;
    wire N__39795;
    wire N__39792;
    wire N__39787;
    wire N__39786;
    wire N__39783;
    wire N__39782;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39768;
    wire N__39765;
    wire N__39760;
    wire N__39757;
    wire N__39754;
    wire N__39751;
    wire N__39748;
    wire N__39745;
    wire N__39742;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39729;
    wire N__39724;
    wire N__39721;
    wire N__39720;
    wire N__39717;
    wire N__39714;
    wire N__39709;
    wire N__39706;
    wire N__39705;
    wire N__39704;
    wire N__39701;
    wire N__39698;
    wire N__39695;
    wire N__39692;
    wire N__39689;
    wire N__39686;
    wire N__39683;
    wire N__39680;
    wire N__39675;
    wire N__39670;
    wire N__39669;
    wire N__39668;
    wire N__39661;
    wire N__39660;
    wire N__39657;
    wire N__39654;
    wire N__39651;
    wire N__39646;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39636;
    wire N__39635;
    wire N__39634;
    wire N__39631;
    wire N__39628;
    wire N__39623;
    wire N__39622;
    wire N__39619;
    wire N__39616;
    wire N__39613;
    wire N__39610;
    wire N__39605;
    wire N__39598;
    wire N__39597;
    wire N__39594;
    wire N__39593;
    wire N__39590;
    wire N__39589;
    wire N__39586;
    wire N__39583;
    wire N__39580;
    wire N__39577;
    wire N__39576;
    wire N__39573;
    wire N__39568;
    wire N__39565;
    wire N__39562;
    wire N__39559;
    wire N__39554;
    wire N__39547;
    wire N__39546;
    wire N__39545;
    wire N__39542;
    wire N__39539;
    wire N__39534;
    wire N__39533;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39523;
    wire N__39522;
    wire N__39519;
    wire N__39514;
    wire N__39511;
    wire N__39508;
    wire N__39505;
    wire N__39496;
    wire N__39495;
    wire N__39494;
    wire N__39491;
    wire N__39488;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39478;
    wire N__39477;
    wire N__39474;
    wire N__39469;
    wire N__39464;
    wire N__39459;
    wire N__39454;
    wire N__39451;
    wire N__39448;
    wire N__39445;
    wire N__39442;
    wire N__39439;
    wire N__39436;
    wire N__39435;
    wire N__39434;
    wire N__39431;
    wire N__39428;
    wire N__39425;
    wire N__39422;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39408;
    wire N__39403;
    wire N__39400;
    wire N__39397;
    wire N__39396;
    wire N__39393;
    wire N__39390;
    wire N__39385;
    wire N__39382;
    wire N__39379;
    wire N__39376;
    wire N__39375;
    wire N__39374;
    wire N__39369;
    wire N__39368;
    wire N__39365;
    wire N__39362;
    wire N__39359;
    wire N__39358;
    wire N__39355;
    wire N__39352;
    wire N__39349;
    wire N__39346;
    wire N__39343;
    wire N__39334;
    wire N__39333;
    wire N__39330;
    wire N__39327;
    wire N__39326;
    wire N__39325;
    wire N__39322;
    wire N__39319;
    wire N__39314;
    wire N__39311;
    wire N__39304;
    wire N__39301;
    wire N__39298;
    wire N__39295;
    wire N__39292;
    wire N__39289;
    wire N__39286;
    wire N__39283;
    wire N__39280;
    wire N__39277;
    wire N__39276;
    wire N__39275;
    wire N__39274;
    wire N__39271;
    wire N__39268;
    wire N__39265;
    wire N__39262;
    wire N__39259;
    wire N__39256;
    wire N__39253;
    wire N__39244;
    wire N__39241;
    wire N__39238;
    wire N__39235;
    wire N__39232;
    wire N__39229;
    wire N__39226;
    wire N__39223;
    wire N__39220;
    wire N__39217;
    wire N__39214;
    wire N__39211;
    wire N__39210;
    wire N__39207;
    wire N__39204;
    wire N__39203;
    wire N__39202;
    wire N__39199;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39183;
    wire N__39180;
    wire N__39175;
    wire N__39172;
    wire N__39163;
    wire N__39160;
    wire N__39159;
    wire N__39156;
    wire N__39153;
    wire N__39152;
    wire N__39151;
    wire N__39148;
    wire N__39145;
    wire N__39140;
    wire N__39133;
    wire N__39132;
    wire N__39129;
    wire N__39128;
    wire N__39127;
    wire N__39126;
    wire N__39123;
    wire N__39120;
    wire N__39117;
    wire N__39114;
    wire N__39111;
    wire N__39108;
    wire N__39103;
    wire N__39094;
    wire N__39091;
    wire N__39090;
    wire N__39087;
    wire N__39084;
    wire N__39083;
    wire N__39082;
    wire N__39077;
    wire N__39074;
    wire N__39073;
    wire N__39070;
    wire N__39067;
    wire N__39064;
    wire N__39061;
    wire N__39058;
    wire N__39049;
    wire N__39048;
    wire N__39045;
    wire N__39042;
    wire N__39039;
    wire N__39038;
    wire N__39035;
    wire N__39032;
    wire N__39029;
    wire N__39022;
    wire N__39021;
    wire N__39018;
    wire N__39015;
    wire N__39014;
    wire N__39013;
    wire N__39010;
    wire N__39007;
    wire N__39004;
    wire N__39001;
    wire N__38998;
    wire N__38993;
    wire N__38986;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38976;
    wire N__38973;
    wire N__38970;
    wire N__38965;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38950;
    wire N__38947;
    wire N__38944;
    wire N__38941;
    wire N__38938;
    wire N__38935;
    wire N__38932;
    wire N__38929;
    wire N__38926;
    wire N__38923;
    wire N__38920;
    wire N__38917;
    wire N__38914;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38902;
    wire N__38899;
    wire N__38896;
    wire N__38893;
    wire N__38892;
    wire N__38891;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38878;
    wire N__38873;
    wire N__38866;
    wire N__38863;
    wire N__38862;
    wire N__38859;
    wire N__38856;
    wire N__38851;
    wire N__38848;
    wire N__38845;
    wire N__38842;
    wire N__38839;
    wire N__38836;
    wire N__38833;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38821;
    wire N__38818;
    wire N__38815;
    wire N__38812;
    wire N__38809;
    wire N__38806;
    wire N__38803;
    wire N__38800;
    wire N__38797;
    wire N__38794;
    wire N__38791;
    wire N__38788;
    wire N__38785;
    wire N__38782;
    wire N__38779;
    wire N__38776;
    wire N__38775;
    wire N__38774;
    wire N__38773;
    wire N__38770;
    wire N__38767;
    wire N__38762;
    wire N__38759;
    wire N__38752;
    wire N__38751;
    wire N__38748;
    wire N__38745;
    wire N__38742;
    wire N__38739;
    wire N__38734;
    wire N__38731;
    wire N__38728;
    wire N__38725;
    wire N__38724;
    wire N__38721;
    wire N__38718;
    wire N__38717;
    wire N__38714;
    wire N__38711;
    wire N__38708;
    wire N__38707;
    wire N__38704;
    wire N__38701;
    wire N__38696;
    wire N__38693;
    wire N__38690;
    wire N__38683;
    wire N__38680;
    wire N__38679;
    wire N__38676;
    wire N__38673;
    wire N__38668;
    wire N__38665;
    wire N__38664;
    wire N__38661;
    wire N__38658;
    wire N__38655;
    wire N__38650;
    wire N__38647;
    wire N__38644;
    wire N__38641;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38626;
    wire N__38625;
    wire N__38622;
    wire N__38619;
    wire N__38616;
    wire N__38611;
    wire N__38608;
    wire N__38607;
    wire N__38604;
    wire N__38601;
    wire N__38600;
    wire N__38597;
    wire N__38594;
    wire N__38591;
    wire N__38586;
    wire N__38581;
    wire N__38580;
    wire N__38577;
    wire N__38574;
    wire N__38571;
    wire N__38570;
    wire N__38569;
    wire N__38564;
    wire N__38561;
    wire N__38558;
    wire N__38555;
    wire N__38552;
    wire N__38545;
    wire N__38542;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38524;
    wire N__38523;
    wire N__38522;
    wire N__38519;
    wire N__38518;
    wire N__38515;
    wire N__38514;
    wire N__38511;
    wire N__38508;
    wire N__38505;
    wire N__38502;
    wire N__38499;
    wire N__38494;
    wire N__38485;
    wire N__38482;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38470;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38462;
    wire N__38459;
    wire N__38456;
    wire N__38455;
    wire N__38452;
    wire N__38447;
    wire N__38444;
    wire N__38441;
    wire N__38440;
    wire N__38439;
    wire N__38436;
    wire N__38431;
    wire N__38426;
    wire N__38419;
    wire N__38416;
    wire N__38415;
    wire N__38412;
    wire N__38409;
    wire N__38404;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38389;
    wire N__38386;
    wire N__38383;
    wire N__38380;
    wire N__38379;
    wire N__38376;
    wire N__38373;
    wire N__38370;
    wire N__38365;
    wire N__38362;
    wire N__38361;
    wire N__38358;
    wire N__38355;
    wire N__38352;
    wire N__38347;
    wire N__38344;
    wire N__38341;
    wire N__38338;
    wire N__38335;
    wire N__38332;
    wire N__38331;
    wire N__38328;
    wire N__38325;
    wire N__38322;
    wire N__38317;
    wire N__38314;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38302;
    wire N__38299;
    wire N__38298;
    wire N__38295;
    wire N__38292;
    wire N__38289;
    wire N__38284;
    wire N__38281;
    wire N__38278;
    wire N__38275;
    wire N__38272;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38262;
    wire N__38257;
    wire N__38254;
    wire N__38253;
    wire N__38250;
    wire N__38247;
    wire N__38242;
    wire N__38241;
    wire N__38238;
    wire N__38235;
    wire N__38232;
    wire N__38229;
    wire N__38224;
    wire N__38223;
    wire N__38220;
    wire N__38217;
    wire N__38214;
    wire N__38209;
    wire N__38206;
    wire N__38205;
    wire N__38202;
    wire N__38199;
    wire N__38194;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38170;
    wire N__38167;
    wire N__38164;
    wire N__38163;
    wire N__38160;
    wire N__38157;
    wire N__38154;
    wire N__38151;
    wire N__38146;
    wire N__38143;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38131;
    wire N__38128;
    wire N__38125;
    wire N__38122;
    wire N__38119;
    wire N__38116;
    wire N__38115;
    wire N__38110;
    wire N__38107;
    wire N__38106;
    wire N__38103;
    wire N__38102;
    wire N__38101;
    wire N__38098;
    wire N__38097;
    wire N__38096;
    wire N__38093;
    wire N__38088;
    wire N__38085;
    wire N__38082;
    wire N__38079;
    wire N__38072;
    wire N__38065;
    wire N__38064;
    wire N__38061;
    wire N__38058;
    wire N__38053;
    wire N__38050;
    wire N__38047;
    wire N__38044;
    wire N__38041;
    wire N__38038;
    wire N__38035;
    wire N__38034;
    wire N__38033;
    wire N__38030;
    wire N__38029;
    wire N__38026;
    wire N__38025;
    wire N__38022;
    wire N__38019;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__37996;
    wire N__37993;
    wire N__37990;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37960;
    wire N__37957;
    wire N__37954;
    wire N__37953;
    wire N__37950;
    wire N__37947;
    wire N__37946;
    wire N__37945;
    wire N__37940;
    wire N__37937;
    wire N__37936;
    wire N__37933;
    wire N__37930;
    wire N__37927;
    wire N__37924;
    wire N__37921;
    wire N__37912;
    wire N__37911;
    wire N__37910;
    wire N__37905;
    wire N__37902;
    wire N__37901;
    wire N__37898;
    wire N__37897;
    wire N__37896;
    wire N__37893;
    wire N__37890;
    wire N__37887;
    wire N__37884;
    wire N__37881;
    wire N__37876;
    wire N__37867;
    wire N__37864;
    wire N__37863;
    wire N__37860;
    wire N__37857;
    wire N__37854;
    wire N__37849;
    wire N__37848;
    wire N__37847;
    wire N__37844;
    wire N__37839;
    wire N__37838;
    wire N__37837;
    wire N__37834;
    wire N__37831;
    wire N__37828;
    wire N__37825;
    wire N__37822;
    wire N__37819;
    wire N__37816;
    wire N__37807;
    wire N__37804;
    wire N__37801;
    wire N__37798;
    wire N__37795;
    wire N__37792;
    wire N__37789;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37774;
    wire N__37771;
    wire N__37768;
    wire N__37767;
    wire N__37766;
    wire N__37763;
    wire N__37760;
    wire N__37757;
    wire N__37756;
    wire N__37753;
    wire N__37748;
    wire N__37745;
    wire N__37738;
    wire N__37737;
    wire N__37736;
    wire N__37733;
    wire N__37732;
    wire N__37731;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37716;
    wire N__37713;
    wire N__37708;
    wire N__37703;
    wire N__37698;
    wire N__37693;
    wire N__37692;
    wire N__37689;
    wire N__37686;
    wire N__37683;
    wire N__37680;
    wire N__37675;
    wire N__37672;
    wire N__37669;
    wire N__37668;
    wire N__37665;
    wire N__37664;
    wire N__37661;
    wire N__37658;
    wire N__37653;
    wire N__37652;
    wire N__37651;
    wire N__37648;
    wire N__37645;
    wire N__37642;
    wire N__37639;
    wire N__37636;
    wire N__37631;
    wire N__37624;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37606;
    wire N__37603;
    wire N__37600;
    wire N__37597;
    wire N__37594;
    wire N__37591;
    wire N__37588;
    wire N__37587;
    wire N__37584;
    wire N__37581;
    wire N__37580;
    wire N__37579;
    wire N__37574;
    wire N__37571;
    wire N__37568;
    wire N__37565;
    wire N__37562;
    wire N__37555;
    wire N__37554;
    wire N__37553;
    wire N__37552;
    wire N__37549;
    wire N__37548;
    wire N__37545;
    wire N__37542;
    wire N__37541;
    wire N__37540;
    wire N__37539;
    wire N__37538;
    wire N__37535;
    wire N__37532;
    wire N__37529;
    wire N__37524;
    wire N__37519;
    wire N__37516;
    wire N__37513;
    wire N__37508;
    wire N__37505;
    wire N__37498;
    wire N__37495;
    wire N__37492;
    wire N__37483;
    wire N__37480;
    wire N__37479;
    wire N__37478;
    wire N__37477;
    wire N__37476;
    wire N__37473;
    wire N__37472;
    wire N__37467;
    wire N__37462;
    wire N__37459;
    wire N__37456;
    wire N__37455;
    wire N__37454;
    wire N__37453;
    wire N__37444;
    wire N__37439;
    wire N__37436;
    wire N__37435;
    wire N__37434;
    wire N__37433;
    wire N__37432;
    wire N__37431;
    wire N__37430;
    wire N__37427;
    wire N__37422;
    wire N__37417;
    wire N__37414;
    wire N__37409;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37387;
    wire N__37384;
    wire N__37383;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37370;
    wire N__37367;
    wire N__37364;
    wire N__37361;
    wire N__37354;
    wire N__37353;
    wire N__37350;
    wire N__37349;
    wire N__37348;
    wire N__37345;
    wire N__37344;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37329;
    wire N__37326;
    wire N__37323;
    wire N__37312;
    wire N__37309;
    wire N__37306;
    wire N__37305;
    wire N__37304;
    wire N__37303;
    wire N__37302;
    wire N__37299;
    wire N__37296;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37281;
    wire N__37276;
    wire N__37267;
    wire N__37264;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37254;
    wire N__37251;
    wire N__37248;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37236;
    wire N__37233;
    wire N__37230;
    wire N__37227;
    wire N__37222;
    wire N__37219;
    wire N__37216;
    wire N__37213;
    wire N__37210;
    wire N__37207;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37195;
    wire N__37192;
    wire N__37191;
    wire N__37188;
    wire N__37185;
    wire N__37180;
    wire N__37177;
    wire N__37174;
    wire N__37171;
    wire N__37168;
    wire N__37165;
    wire N__37162;
    wire N__37159;
    wire N__37156;
    wire N__37153;
    wire N__37150;
    wire N__37149;
    wire N__37148;
    wire N__37147;
    wire N__37144;
    wire N__37141;
    wire N__37138;
    wire N__37135;
    wire N__37126;
    wire N__37123;
    wire N__37120;
    wire N__37117;
    wire N__37116;
    wire N__37113;
    wire N__37110;
    wire N__37109;
    wire N__37106;
    wire N__37105;
    wire N__37102;
    wire N__37099;
    wire N__37096;
    wire N__37093;
    wire N__37090;
    wire N__37081;
    wire N__37078;
    wire N__37077;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37065;
    wire N__37060;
    wire N__37057;
    wire N__37054;
    wire N__37053;
    wire N__37050;
    wire N__37047;
    wire N__37044;
    wire N__37043;
    wire N__37042;
    wire N__37041;
    wire N__37036;
    wire N__37033;
    wire N__37028;
    wire N__37021;
    wire N__37018;
    wire N__37015;
    wire N__37012;
    wire N__37009;
    wire N__37006;
    wire N__37003;
    wire N__37000;
    wire N__36997;
    wire N__36994;
    wire N__36991;
    wire N__36988;
    wire N__36987;
    wire N__36984;
    wire N__36981;
    wire N__36978;
    wire N__36975;
    wire N__36972;
    wire N__36967;
    wire N__36964;
    wire N__36961;
    wire N__36958;
    wire N__36955;
    wire N__36952;
    wire N__36949;
    wire N__36946;
    wire N__36943;
    wire N__36940;
    wire N__36937;
    wire N__36934;
    wire N__36931;
    wire N__36928;
    wire N__36925;
    wire N__36922;
    wire N__36919;
    wire N__36916;
    wire N__36913;
    wire N__36910;
    wire N__36907;
    wire N__36904;
    wire N__36901;
    wire N__36898;
    wire N__36895;
    wire N__36892;
    wire N__36889;
    wire N__36888;
    wire N__36885;
    wire N__36882;
    wire N__36877;
    wire N__36874;
    wire N__36871;
    wire N__36870;
    wire N__36867;
    wire N__36864;
    wire N__36861;
    wire N__36856;
    wire N__36853;
    wire N__36850;
    wire N__36849;
    wire N__36846;
    wire N__36843;
    wire N__36838;
    wire N__36835;
    wire N__36832;
    wire N__36829;
    wire N__36828;
    wire N__36827;
    wire N__36824;
    wire N__36821;
    wire N__36820;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36803;
    wire N__36796;
    wire N__36793;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36781;
    wire N__36778;
    wire N__36775;
    wire N__36772;
    wire N__36769;
    wire N__36766;
    wire N__36763;
    wire N__36760;
    wire N__36757;
    wire N__36756;
    wire N__36753;
    wire N__36750;
    wire N__36747;
    wire N__36744;
    wire N__36741;
    wire N__36736;
    wire N__36735;
    wire N__36732;
    wire N__36731;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36718;
    wire N__36715;
    wire N__36712;
    wire N__36709;
    wire N__36708;
    wire N__36705;
    wire N__36702;
    wire N__36699;
    wire N__36696;
    wire N__36693;
    wire N__36690;
    wire N__36679;
    wire N__36676;
    wire N__36673;
    wire N__36670;
    wire N__36669;
    wire N__36666;
    wire N__36663;
    wire N__36660;
    wire N__36655;
    wire N__36652;
    wire N__36649;
    wire N__36646;
    wire N__36645;
    wire N__36642;
    wire N__36639;
    wire N__36636;
    wire N__36631;
    wire N__36628;
    wire N__36625;
    wire N__36622;
    wire N__36621;
    wire N__36620;
    wire N__36619;
    wire N__36616;
    wire N__36613;
    wire N__36610;
    wire N__36609;
    wire N__36606;
    wire N__36603;
    wire N__36600;
    wire N__36597;
    wire N__36596;
    wire N__36593;
    wire N__36590;
    wire N__36587;
    wire N__36582;
    wire N__36579;
    wire N__36576;
    wire N__36565;
    wire N__36562;
    wire N__36559;
    wire N__36556;
    wire N__36555;
    wire N__36552;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36538;
    wire N__36535;
    wire N__36532;
    wire N__36529;
    wire N__36528;
    wire N__36525;
    wire N__36522;
    wire N__36517;
    wire N__36514;
    wire N__36511;
    wire N__36508;
    wire N__36507;
    wire N__36504;
    wire N__36501;
    wire N__36496;
    wire N__36493;
    wire N__36492;
    wire N__36489;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36475;
    wire N__36472;
    wire N__36469;
    wire N__36466;
    wire N__36465;
    wire N__36462;
    wire N__36459;
    wire N__36454;
    wire N__36451;
    wire N__36448;
    wire N__36445;
    wire N__36442;
    wire N__36441;
    wire N__36440;
    wire N__36439;
    wire N__36436;
    wire N__36433;
    wire N__36428;
    wire N__36425;
    wire N__36424;
    wire N__36419;
    wire N__36418;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36406;
    wire N__36401;
    wire N__36394;
    wire N__36391;
    wire N__36390;
    wire N__36387;
    wire N__36384;
    wire N__36381;
    wire N__36376;
    wire N__36373;
    wire N__36372;
    wire N__36369;
    wire N__36366;
    wire N__36363;
    wire N__36358;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36346;
    wire N__36343;
    wire N__36340;
    wire N__36339;
    wire N__36336;
    wire N__36333;
    wire N__36330;
    wire N__36327;
    wire N__36322;
    wire N__36319;
    wire N__36316;
    wire N__36313;
    wire N__36312;
    wire N__36309;
    wire N__36306;
    wire N__36303;
    wire N__36300;
    wire N__36295;
    wire N__36292;
    wire N__36289;
    wire N__36286;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36274;
    wire N__36271;
    wire N__36268;
    wire N__36267;
    wire N__36264;
    wire N__36261;
    wire N__36258;
    wire N__36255;
    wire N__36250;
    wire N__36249;
    wire N__36246;
    wire N__36245;
    wire N__36242;
    wire N__36239;
    wire N__36236;
    wire N__36233;
    wire N__36232;
    wire N__36231;
    wire N__36228;
    wire N__36225;
    wire N__36224;
    wire N__36221;
    wire N__36218;
    wire N__36215;
    wire N__36212;
    wire N__36209;
    wire N__36206;
    wire N__36201;
    wire N__36190;
    wire N__36187;
    wire N__36184;
    wire N__36181;
    wire N__36178;
    wire N__36175;
    wire N__36172;
    wire N__36169;
    wire N__36166;
    wire N__36163;
    wire N__36160;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36148;
    wire N__36145;
    wire N__36142;
    wire N__36139;
    wire N__36136;
    wire N__36133;
    wire N__36130;
    wire N__36127;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36112;
    wire N__36109;
    wire N__36108;
    wire N__36105;
    wire N__36102;
    wire N__36097;
    wire N__36094;
    wire N__36091;
    wire N__36088;
    wire N__36085;
    wire N__36082;
    wire N__36079;
    wire N__36076;
    wire N__36075;
    wire N__36074;
    wire N__36073;
    wire N__36070;
    wire N__36069;
    wire N__36066;
    wire N__36061;
    wire N__36058;
    wire N__36055;
    wire N__36052;
    wire N__36043;
    wire N__36042;
    wire N__36041;
    wire N__36038;
    wire N__36033;
    wire N__36028;
    wire N__36025;
    wire N__36022;
    wire N__36019;
    wire N__36016;
    wire N__36013;
    wire N__36010;
    wire N__36007;
    wire N__36004;
    wire N__36001;
    wire N__35998;
    wire N__35995;
    wire N__35992;
    wire N__35989;
    wire N__35986;
    wire N__35983;
    wire N__35980;
    wire N__35977;
    wire N__35974;
    wire N__35971;
    wire N__35968;
    wire N__35965;
    wire N__35962;
    wire N__35959;
    wire N__35956;
    wire N__35953;
    wire N__35950;
    wire N__35947;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35937;
    wire N__35934;
    wire N__35931;
    wire N__35928;
    wire N__35925;
    wire N__35922;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35908;
    wire N__35905;
    wire N__35902;
    wire N__35899;
    wire N__35896;
    wire N__35893;
    wire N__35892;
    wire N__35887;
    wire N__35884;
    wire N__35881;
    wire N__35878;
    wire N__35875;
    wire N__35874;
    wire N__35873;
    wire N__35870;
    wire N__35869;
    wire N__35866;
    wire N__35863;
    wire N__35860;
    wire N__35857;
    wire N__35854;
    wire N__35853;
    wire N__35846;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35830;
    wire N__35827;
    wire N__35824;
    wire N__35821;
    wire N__35818;
    wire N__35815;
    wire N__35814;
    wire N__35811;
    wire N__35810;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35800;
    wire N__35797;
    wire N__35794;
    wire N__35791;
    wire N__35788;
    wire N__35779;
    wire N__35776;
    wire N__35773;
    wire N__35772;
    wire N__35769;
    wire N__35768;
    wire N__35767;
    wire N__35764;
    wire N__35763;
    wire N__35762;
    wire N__35761;
    wire N__35760;
    wire N__35753;
    wire N__35746;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35734;
    wire N__35731;
    wire N__35728;
    wire N__35725;
    wire N__35722;
    wire N__35717;
    wire N__35714;
    wire N__35711;
    wire N__35708;
    wire N__35701;
    wire N__35700;
    wire N__35697;
    wire N__35694;
    wire N__35691;
    wire N__35686;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35674;
    wire N__35671;
    wire N__35668;
    wire N__35665;
    wire N__35662;
    wire N__35659;
    wire N__35656;
    wire N__35653;
    wire N__35650;
    wire N__35647;
    wire N__35644;
    wire N__35641;
    wire N__35638;
    wire N__35635;
    wire N__35632;
    wire N__35629;
    wire N__35626;
    wire N__35623;
    wire N__35620;
    wire N__35617;
    wire N__35616;
    wire N__35615;
    wire N__35612;
    wire N__35609;
    wire N__35606;
    wire N__35605;
    wire N__35604;
    wire N__35603;
    wire N__35602;
    wire N__35599;
    wire N__35596;
    wire N__35593;
    wire N__35590;
    wire N__35587;
    wire N__35584;
    wire N__35581;
    wire N__35576;
    wire N__35571;
    wire N__35568;
    wire N__35565;
    wire N__35564;
    wire N__35561;
    wire N__35556;
    wire N__35551;
    wire N__35548;
    wire N__35545;
    wire N__35542;
    wire N__35539;
    wire N__35534;
    wire N__35527;
    wire N__35524;
    wire N__35523;
    wire N__35522;
    wire N__35521;
    wire N__35520;
    wire N__35519;
    wire N__35518;
    wire N__35515;
    wire N__35512;
    wire N__35511;
    wire N__35508;
    wire N__35505;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35490;
    wire N__35487;
    wire N__35484;
    wire N__35479;
    wire N__35472;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35460;
    wire N__35457;
    wire N__35454;
    wire N__35443;
    wire N__35440;
    wire N__35437;
    wire N__35434;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35424;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35391;
    wire N__35390;
    wire N__35387;
    wire N__35386;
    wire N__35385;
    wire N__35382;
    wire N__35381;
    wire N__35380;
    wire N__35377;
    wire N__35374;
    wire N__35369;
    wire N__35360;
    wire N__35357;
    wire N__35350;
    wire N__35349;
    wire N__35348;
    wire N__35347;
    wire N__35344;
    wire N__35343;
    wire N__35342;
    wire N__35335;
    wire N__35332;
    wire N__35329;
    wire N__35326;
    wire N__35321;
    wire N__35314;
    wire N__35311;
    wire N__35308;
    wire N__35305;
    wire N__35304;
    wire N__35301;
    wire N__35298;
    wire N__35293;
    wire N__35290;
    wire N__35287;
    wire N__35286;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35272;
    wire N__35271;
    wire N__35268;
    wire N__35265;
    wire N__35260;
    wire N__35257;
    wire N__35254;
    wire N__35251;
    wire N__35248;
    wire N__35247;
    wire N__35242;
    wire N__35239;
    wire N__35238;
    wire N__35237;
    wire N__35236;
    wire N__35233;
    wire N__35232;
    wire N__35227;
    wire N__35224;
    wire N__35219;
    wire N__35216;
    wire N__35215;
    wire N__35212;
    wire N__35209;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35185;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35170;
    wire N__35167;
    wire N__35166;
    wire N__35165;
    wire N__35160;
    wire N__35159;
    wire N__35156;
    wire N__35153;
    wire N__35150;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35134;
    wire N__35131;
    wire N__35128;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35086;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35071;
    wire N__35068;
    wire N__35065;
    wire N__35064;
    wire N__35063;
    wire N__35062;
    wire N__35059;
    wire N__35056;
    wire N__35053;
    wire N__35050;
    wire N__35047;
    wire N__35038;
    wire N__35037;
    wire N__35036;
    wire N__35035;
    wire N__35034;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35022;
    wire N__35019;
    wire N__35018;
    wire N__35017;
    wire N__35014;
    wire N__35005;
    wire N__35004;
    wire N__35001;
    wire N__34998;
    wire N__34993;
    wire N__34990;
    wire N__34981;
    wire N__34978;
    wire N__34977;
    wire N__34976;
    wire N__34973;
    wire N__34970;
    wire N__34967;
    wire N__34964;
    wire N__34961;
    wire N__34958;
    wire N__34957;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34930;
    wire N__34927;
    wire N__34924;
    wire N__34921;
    wire N__34918;
    wire N__34915;
    wire N__34914;
    wire N__34913;
    wire N__34912;
    wire N__34909;
    wire N__34906;
    wire N__34903;
    wire N__34900;
    wire N__34891;
    wire N__34888;
    wire N__34885;
    wire N__34882;
    wire N__34879;
    wire N__34876;
    wire N__34873;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34855;
    wire N__34852;
    wire N__34849;
    wire N__34846;
    wire N__34843;
    wire N__34840;
    wire N__34837;
    wire N__34834;
    wire N__34831;
    wire N__34828;
    wire N__34825;
    wire N__34822;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34810;
    wire N__34807;
    wire N__34806;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34792;
    wire N__34789;
    wire N__34786;
    wire N__34785;
    wire N__34782;
    wire N__34779;
    wire N__34776;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34756;
    wire N__34753;
    wire N__34752;
    wire N__34749;
    wire N__34746;
    wire N__34743;
    wire N__34738;
    wire N__34735;
    wire N__34732;
    wire N__34729;
    wire N__34728;
    wire N__34725;
    wire N__34722;
    wire N__34719;
    wire N__34714;
    wire N__34711;
    wire N__34708;
    wire N__34705;
    wire N__34704;
    wire N__34701;
    wire N__34698;
    wire N__34695;
    wire N__34690;
    wire N__34687;
    wire N__34684;
    wire N__34683;
    wire N__34680;
    wire N__34677;
    wire N__34672;
    wire N__34669;
    wire N__34666;
    wire N__34663;
    wire N__34662;
    wire N__34661;
    wire N__34660;
    wire N__34659;
    wire N__34656;
    wire N__34655;
    wire N__34654;
    wire N__34653;
    wire N__34652;
    wire N__34651;
    wire N__34650;
    wire N__34649;
    wire N__34648;
    wire N__34647;
    wire N__34646;
    wire N__34645;
    wire N__34644;
    wire N__34643;
    wire N__34642;
    wire N__34641;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34629;
    wire N__34626;
    wire N__34623;
    wire N__34620;
    wire N__34617;
    wire N__34614;
    wire N__34613;
    wire N__34610;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34598;
    wire N__34595;
    wire N__34592;
    wire N__34589;
    wire N__34586;
    wire N__34583;
    wire N__34580;
    wire N__34577;
    wire N__34574;
    wire N__34565;
    wire N__34564;
    wire N__34563;
    wire N__34562;
    wire N__34561;
    wire N__34560;
    wire N__34559;
    wire N__34558;
    wire N__34555;
    wire N__34550;
    wire N__34547;
    wire N__34544;
    wire N__34537;
    wire N__34530;
    wire N__34527;
    wire N__34524;
    wire N__34521;
    wire N__34516;
    wire N__34511;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34499;
    wire N__34496;
    wire N__34493;
    wire N__34490;
    wire N__34485;
    wire N__34476;
    wire N__34467;
    wire N__34464;
    wire N__34441;
    wire N__34438;
    wire N__34435;
    wire N__34432;
    wire N__34431;
    wire N__34430;
    wire N__34427;
    wire N__34424;
    wire N__34421;
    wire N__34418;
    wire N__34411;
    wire N__34408;
    wire N__34405;
    wire N__34402;
    wire N__34399;
    wire N__34396;
    wire N__34393;
    wire N__34392;
    wire N__34389;
    wire N__34386;
    wire N__34383;
    wire N__34378;
    wire N__34375;
    wire N__34372;
    wire N__34369;
    wire N__34366;
    wire N__34363;
    wire N__34360;
    wire N__34357;
    wire N__34356;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34348;
    wire N__34345;
    wire N__34342;
    wire N__34339;
    wire N__34336;
    wire N__34333;
    wire N__34330;
    wire N__34321;
    wire N__34318;
    wire N__34317;
    wire N__34314;
    wire N__34311;
    wire N__34310;
    wire N__34309;
    wire N__34304;
    wire N__34299;
    wire N__34294;
    wire N__34291;
    wire N__34288;
    wire N__34285;
    wire N__34282;
    wire N__34281;
    wire N__34280;
    wire N__34277;
    wire N__34276;
    wire N__34275;
    wire N__34272;
    wire N__34269;
    wire N__34266;
    wire N__34263;
    wire N__34262;
    wire N__34259;
    wire N__34256;
    wire N__34249;
    wire N__34248;
    wire N__34247;
    wire N__34246;
    wire N__34243;
    wire N__34238;
    wire N__34235;
    wire N__34228;
    wire N__34219;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34204;
    wire N__34201;
    wire N__34198;
    wire N__34197;
    wire N__34196;
    wire N__34195;
    wire N__34194;
    wire N__34189;
    wire N__34186;
    wire N__34181;
    wire N__34176;
    wire N__34171;
    wire N__34168;
    wire N__34165;
    wire N__34162;
    wire N__34159;
    wire N__34156;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34140;
    wire N__34137;
    wire N__34134;
    wire N__34133;
    wire N__34130;
    wire N__34127;
    wire N__34124;
    wire N__34121;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34096;
    wire N__34093;
    wire N__34090;
    wire N__34087;
    wire N__34084;
    wire N__34081;
    wire N__34078;
    wire N__34075;
    wire N__34074;
    wire N__34071;
    wire N__34068;
    wire N__34065;
    wire N__34060;
    wire N__34057;
    wire N__34054;
    wire N__34053;
    wire N__34050;
    wire N__34047;
    wire N__34044;
    wire N__34039;
    wire N__34036;
    wire N__34035;
    wire N__34032;
    wire N__34029;
    wire N__34024;
    wire N__34021;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34009;
    wire N__34006;
    wire N__34003;
    wire N__34000;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33987;
    wire N__33984;
    wire N__33981;
    wire N__33976;
    wire N__33973;
    wire N__33972;
    wire N__33969;
    wire N__33966;
    wire N__33963;
    wire N__33958;
    wire N__33955;
    wire N__33952;
    wire N__33949;
    wire N__33946;
    wire N__33943;
    wire N__33940;
    wire N__33937;
    wire N__33934;
    wire N__33931;
    wire N__33928;
    wire N__33925;
    wire N__33922;
    wire N__33919;
    wire N__33916;
    wire N__33913;
    wire N__33910;
    wire N__33907;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33885;
    wire N__33882;
    wire N__33881;
    wire N__33880;
    wire N__33877;
    wire N__33876;
    wire N__33875;
    wire N__33874;
    wire N__33871;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33859;
    wire N__33858;
    wire N__33855;
    wire N__33852;
    wire N__33849;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33834;
    wire N__33829;
    wire N__33822;
    wire N__33819;
    wire N__33816;
    wire N__33813;
    wire N__33810;
    wire N__33807;
    wire N__33798;
    wire N__33795;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33780;
    wire N__33777;
    wire N__33774;
    wire N__33771;
    wire N__33766;
    wire N__33765;
    wire N__33764;
    wire N__33763;
    wire N__33760;
    wire N__33759;
    wire N__33758;
    wire N__33755;
    wire N__33754;
    wire N__33753;
    wire N__33748;
    wire N__33747;
    wire N__33746;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33731;
    wire N__33728;
    wire N__33725;
    wire N__33722;
    wire N__33719;
    wire N__33716;
    wire N__33713;
    wire N__33710;
    wire N__33707;
    wire N__33704;
    wire N__33699;
    wire N__33696;
    wire N__33689;
    wire N__33684;
    wire N__33681;
    wire N__33676;
    wire N__33671;
    wire N__33666;
    wire N__33661;
    wire N__33658;
    wire N__33655;
    wire N__33652;
    wire N__33649;
    wire N__33646;
    wire N__33643;
    wire N__33640;
    wire N__33639;
    wire N__33634;
    wire N__33631;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33619;
    wire N__33616;
    wire N__33613;
    wire N__33610;
    wire N__33607;
    wire N__33604;
    wire N__33601;
    wire N__33598;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33564;
    wire N__33561;
    wire N__33558;
    wire N__33557;
    wire N__33556;
    wire N__33553;
    wire N__33548;
    wire N__33545;
    wire N__33538;
    wire N__33535;
    wire N__33534;
    wire N__33533;
    wire N__33532;
    wire N__33531;
    wire N__33530;
    wire N__33527;
    wire N__33524;
    wire N__33523;
    wire N__33522;
    wire N__33521;
    wire N__33518;
    wire N__33517;
    wire N__33516;
    wire N__33515;
    wire N__33512;
    wire N__33509;
    wire N__33506;
    wire N__33501;
    wire N__33494;
    wire N__33493;
    wire N__33490;
    wire N__33487;
    wire N__33482;
    wire N__33479;
    wire N__33478;
    wire N__33477;
    wire N__33476;
    wire N__33467;
    wire N__33464;
    wire N__33455;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33433;
    wire N__33430;
    wire N__33429;
    wire N__33426;
    wire N__33425;
    wire N__33422;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33412;
    wire N__33409;
    wire N__33406;
    wire N__33403;
    wire N__33402;
    wire N__33401;
    wire N__33398;
    wire N__33397;
    wire N__33392;
    wire N__33389;
    wire N__33386;
    wire N__33383;
    wire N__33380;
    wire N__33377;
    wire N__33372;
    wire N__33365;
    wire N__33358;
    wire N__33357;
    wire N__33356;
    wire N__33353;
    wire N__33352;
    wire N__33349;
    wire N__33346;
    wire N__33343;
    wire N__33340;
    wire N__33335;
    wire N__33328;
    wire N__33325;
    wire N__33322;
    wire N__33321;
    wire N__33320;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33295;
    wire N__33292;
    wire N__33289;
    wire N__33286;
    wire N__33283;
    wire N__33280;
    wire N__33279;
    wire N__33278;
    wire N__33277;
    wire N__33276;
    wire N__33273;
    wire N__33270;
    wire N__33269;
    wire N__33268;
    wire N__33267;
    wire N__33266;
    wire N__33265;
    wire N__33262;
    wire N__33261;
    wire N__33260;
    wire N__33259;
    wire N__33258;
    wire N__33257;
    wire N__33256;
    wire N__33255;
    wire N__33254;
    wire N__33251;
    wire N__33248;
    wire N__33247;
    wire N__33242;
    wire N__33239;
    wire N__33236;
    wire N__33233;
    wire N__33230;
    wire N__33227;
    wire N__33226;
    wire N__33225;
    wire N__33222;
    wire N__33219;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33209;
    wire N__33208;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33195;
    wire N__33190;
    wire N__33187;
    wire N__33186;
    wire N__33185;
    wire N__33184;
    wire N__33183;
    wire N__33182;
    wire N__33181;
    wire N__33168;
    wire N__33165;
    wire N__33162;
    wire N__33161;
    wire N__33150;
    wire N__33147;
    wire N__33144;
    wire N__33135;
    wire N__33132;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33102;
    wire N__33099;
    wire N__33098;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33079;
    wire N__33076;
    wire N__33073;
    wire N__33068;
    wire N__33065;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33053;
    wire N__33048;
    wire N__33045;
    wire N__33040;
    wire N__33037;
    wire N__33030;
    wire N__33027;
    wire N__33022;
    wire N__33007;
    wire N__33006;
    wire N__33005;
    wire N__33004;
    wire N__33003;
    wire N__33002;
    wire N__33001;
    wire N__33000;
    wire N__32999;
    wire N__32998;
    wire N__32997;
    wire N__32996;
    wire N__32993;
    wire N__32990;
    wire N__32989;
    wire N__32988;
    wire N__32985;
    wire N__32982;
    wire N__32979;
    wire N__32976;
    wire N__32973;
    wire N__32970;
    wire N__32967;
    wire N__32964;
    wire N__32961;
    wire N__32960;
    wire N__32959;
    wire N__32956;
    wire N__32951;
    wire N__32948;
    wire N__32947;
    wire N__32946;
    wire N__32943;
    wire N__32938;
    wire N__32935;
    wire N__32922;
    wire N__32919;
    wire N__32918;
    wire N__32915;
    wire N__32914;
    wire N__32913;
    wire N__32912;
    wire N__32911;
    wire N__32910;
    wire N__32903;
    wire N__32900;
    wire N__32897;
    wire N__32896;
    wire N__32895;
    wire N__32894;
    wire N__32893;
    wire N__32892;
    wire N__32889;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32859;
    wire N__32852;
    wire N__32849;
    wire N__32848;
    wire N__32847;
    wire N__32842;
    wire N__32839;
    wire N__32836;
    wire N__32835;
    wire N__32834;
    wire N__32827;
    wire N__32826;
    wire N__32823;
    wire N__32816;
    wire N__32807;
    wire N__32804;
    wire N__32803;
    wire N__32802;
    wire N__32799;
    wire N__32796;
    wire N__32791;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32783;
    wire N__32780;
    wire N__32777;
    wire N__32768;
    wire N__32765;
    wire N__32762;
    wire N__32755;
    wire N__32752;
    wire N__32747;
    wire N__32744;
    wire N__32725;
    wire N__32722;
    wire N__32719;
    wire N__32716;
    wire N__32713;
    wire N__32710;
    wire N__32709;
    wire N__32706;
    wire N__32705;
    wire N__32704;
    wire N__32701;
    wire N__32698;
    wire N__32695;
    wire N__32692;
    wire N__32691;
    wire N__32690;
    wire N__32687;
    wire N__32682;
    wire N__32679;
    wire N__32676;
    wire N__32673;
    wire N__32670;
    wire N__32669;
    wire N__32666;
    wire N__32659;
    wire N__32656;
    wire N__32653;
    wire N__32650;
    wire N__32645;
    wire N__32642;
    wire N__32639;
    wire N__32636;
    wire N__32633;
    wire N__32626;
    wire N__32623;
    wire N__32620;
    wire N__32617;
    wire N__32614;
    wire N__32611;
    wire N__32610;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32600;
    wire N__32597;
    wire N__32590;
    wire N__32589;
    wire N__32588;
    wire N__32585;
    wire N__32584;
    wire N__32583;
    wire N__32578;
    wire N__32575;
    wire N__32572;
    wire N__32571;
    wire N__32568;
    wire N__32567;
    wire N__32566;
    wire N__32563;
    wire N__32560;
    wire N__32549;
    wire N__32542;
    wire N__32539;
    wire N__32536;
    wire N__32533;
    wire N__32530;
    wire N__32529;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32515;
    wire N__32512;
    wire N__32509;
    wire N__32506;
    wire N__32503;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32491;
    wire N__32488;
    wire N__32485;
    wire N__32482;
    wire N__32479;
    wire N__32478;
    wire N__32475;
    wire N__32472;
    wire N__32467;
    wire N__32464;
    wire N__32461;
    wire N__32458;
    wire N__32455;
    wire N__32454;
    wire N__32451;
    wire N__32448;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32438;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32424;
    wire N__32419;
    wire N__32416;
    wire N__32413;
    wire N__32410;
    wire N__32407;
    wire N__32404;
    wire N__32403;
    wire N__32398;
    wire N__32397;
    wire N__32396;
    wire N__32393;
    wire N__32390;
    wire N__32389;
    wire N__32386;
    wire N__32383;
    wire N__32380;
    wire N__32377;
    wire N__32368;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32344;
    wire N__32341;
    wire N__32338;
    wire N__32335;
    wire N__32332;
    wire N__32329;
    wire N__32326;
    wire N__32325;
    wire N__32324;
    wire N__32319;
    wire N__32318;
    wire N__32317;
    wire N__32314;
    wire N__32311;
    wire N__32310;
    wire N__32307;
    wire N__32306;
    wire N__32303;
    wire N__32300;
    wire N__32299;
    wire N__32296;
    wire N__32293;
    wire N__32292;
    wire N__32289;
    wire N__32286;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32272;
    wire N__32269;
    wire N__32268;
    wire N__32265;
    wire N__32262;
    wire N__32261;
    wire N__32260;
    wire N__32253;
    wire N__32248;
    wire N__32245;
    wire N__32240;
    wire N__32235;
    wire N__32232;
    wire N__32229;
    wire N__32218;
    wire N__32215;
    wire N__32212;
    wire N__32209;
    wire N__32206;
    wire N__32203;
    wire N__32200;
    wire N__32197;
    wire N__32194;
    wire N__32193;
    wire N__32192;
    wire N__32191;
    wire N__32190;
    wire N__32187;
    wire N__32182;
    wire N__32177;
    wire N__32170;
    wire N__32169;
    wire N__32166;
    wire N__32163;
    wire N__32158;
    wire N__32155;
    wire N__32152;
    wire N__32149;
    wire N__32146;
    wire N__32143;
    wire N__32140;
    wire N__32137;
    wire N__32134;
    wire N__32131;
    wire N__32128;
    wire N__32125;
    wire N__32122;
    wire N__32121;
    wire N__32118;
    wire N__32115;
    wire N__32112;
    wire N__32107;
    wire N__32104;
    wire N__32101;
    wire N__32098;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32086;
    wire N__32083;
    wire N__32082;
    wire N__32079;
    wire N__32076;
    wire N__32073;
    wire N__32068;
    wire N__32067;
    wire N__32062;
    wire N__32059;
    wire N__32056;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32041;
    wire N__32038;
    wire N__32035;
    wire N__32032;
    wire N__32029;
    wire N__32026;
    wire N__32023;
    wire N__32020;
    wire N__32017;
    wire N__32014;
    wire N__32011;
    wire N__32008;
    wire N__32007;
    wire N__32002;
    wire N__32001;
    wire N__32000;
    wire N__31999;
    wire N__31998;
    wire N__31997;
    wire N__31996;
    wire N__31995;
    wire N__31994;
    wire N__31993;
    wire N__31992;
    wire N__31991;
    wire N__31990;
    wire N__31989;
    wire N__31988;
    wire N__31985;
    wire N__31976;
    wire N__31967;
    wire N__31964;
    wire N__31961;
    wire N__31956;
    wire N__31951;
    wire N__31936;
    wire N__31935;
    wire N__31934;
    wire N__31933;
    wire N__31926;
    wire N__31925;
    wire N__31924;
    wire N__31923;
    wire N__31922;
    wire N__31921;
    wire N__31920;
    wire N__31919;
    wire N__31918;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31908;
    wire N__31905;
    wire N__31896;
    wire N__31893;
    wire N__31888;
    wire N__31885;
    wire N__31880;
    wire N__31879;
    wire N__31878;
    wire N__31877;
    wire N__31874;
    wire N__31867;
    wire N__31864;
    wire N__31861;
    wire N__31856;
    wire N__31853;
    wire N__31848;
    wire N__31839;
    wire N__31834;
    wire N__31831;
    wire N__31830;
    wire N__31827;
    wire N__31826;
    wire N__31823;
    wire N__31820;
    wire N__31819;
    wire N__31816;
    wire N__31813;
    wire N__31812;
    wire N__31809;
    wire N__31804;
    wire N__31801;
    wire N__31798;
    wire N__31797;
    wire N__31796;
    wire N__31795;
    wire N__31794;
    wire N__31789;
    wire N__31784;
    wire N__31781;
    wire N__31778;
    wire N__31775;
    wire N__31772;
    wire N__31759;
    wire N__31758;
    wire N__31755;
    wire N__31752;
    wire N__31749;
    wire N__31744;
    wire N__31741;
    wire N__31738;
    wire N__31737;
    wire N__31736;
    wire N__31735;
    wire N__31732;
    wire N__31729;
    wire N__31728;
    wire N__31725;
    wire N__31722;
    wire N__31721;
    wire N__31718;
    wire N__31715;
    wire N__31712;
    wire N__31707;
    wire N__31706;
    wire N__31703;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31687;
    wire N__31684;
    wire N__31681;
    wire N__31672;
    wire N__31671;
    wire N__31670;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31660;
    wire N__31657;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31645;
    wire N__31644;
    wire N__31643;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31633;
    wire N__31630;
    wire N__31623;
    wire N__31612;
    wire N__31609;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31592;
    wire N__31589;
    wire N__31584;
    wire N__31579;
    wire N__31576;
    wire N__31573;
    wire N__31572;
    wire N__31567;
    wire N__31564;
    wire N__31561;
    wire N__31558;
    wire N__31555;
    wire N__31552;
    wire N__31551;
    wire N__31550;
    wire N__31547;
    wire N__31546;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31536;
    wire N__31533;
    wire N__31532;
    wire N__31529;
    wire N__31526;
    wire N__31525;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31514;
    wire N__31513;
    wire N__31510;
    wire N__31505;
    wire N__31500;
    wire N__31499;
    wire N__31498;
    wire N__31497;
    wire N__31496;
    wire N__31489;
    wire N__31488;
    wire N__31487;
    wire N__31486;
    wire N__31485;
    wire N__31482;
    wire N__31481;
    wire N__31478;
    wire N__31475;
    wire N__31470;
    wire N__31467;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31449;
    wire N__31442;
    wire N__31435;
    wire N__31420;
    wire N__31417;
    wire N__31414;
    wire N__31411;
    wire N__31408;
    wire N__31407;
    wire N__31404;
    wire N__31403;
    wire N__31400;
    wire N__31397;
    wire N__31394;
    wire N__31389;
    wire N__31384;
    wire N__31383;
    wire N__31380;
    wire N__31379;
    wire N__31378;
    wire N__31377;
    wire N__31374;
    wire N__31371;
    wire N__31368;
    wire N__31365;
    wire N__31362;
    wire N__31361;
    wire N__31356;
    wire N__31353;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31343;
    wire N__31338;
    wire N__31333;
    wire N__31330;
    wire N__31327;
    wire N__31322;
    wire N__31315;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31294;
    wire N__31293;
    wire N__31288;
    wire N__31285;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31273;
    wire N__31270;
    wire N__31267;
    wire N__31264;
    wire N__31261;
    wire N__31258;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31240;
    wire N__31237;
    wire N__31234;
    wire N__31231;
    wire N__31230;
    wire N__31229;
    wire N__31228;
    wire N__31225;
    wire N__31222;
    wire N__31221;
    wire N__31218;
    wire N__31217;
    wire N__31216;
    wire N__31213;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31202;
    wire N__31199;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31181;
    wire N__31178;
    wire N__31175;
    wire N__31172;
    wire N__31169;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31150;
    wire N__31141;
    wire N__31138;
    wire N__31137;
    wire N__31136;
    wire N__31135;
    wire N__31134;
    wire N__31133;
    wire N__31130;
    wire N__31127;
    wire N__31124;
    wire N__31121;
    wire N__31116;
    wire N__31115;
    wire N__31114;
    wire N__31113;
    wire N__31112;
    wire N__31111;
    wire N__31110;
    wire N__31109;
    wire N__31108;
    wire N__31107;
    wire N__31104;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31086;
    wire N__31079;
    wire N__31072;
    wire N__31057;
    wire N__31054;
    wire N__31053;
    wire N__31050;
    wire N__31047;
    wire N__31044;
    wire N__31039;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31029;
    wire N__31028;
    wire N__31027;
    wire N__31026;
    wire N__31023;
    wire N__31022;
    wire N__31021;
    wire N__31018;
    wire N__31015;
    wire N__31014;
    wire N__31013;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__31001;
    wire N__30998;
    wire N__30997;
    wire N__30996;
    wire N__30995;
    wire N__30994;
    wire N__30989;
    wire N__30986;
    wire N__30983;
    wire N__30974;
    wire N__30969;
    wire N__30964;
    wire N__30961;
    wire N__30958;
    wire N__30943;
    wire N__30940;
    wire N__30937;
    wire N__30934;
    wire N__30931;
    wire N__30928;
    wire N__30925;
    wire N__30922;
    wire N__30919;
    wire N__30916;
    wire N__30913;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30898;
    wire N__30897;
    wire N__30894;
    wire N__30891;
    wire N__30888;
    wire N__30883;
    wire N__30880;
    wire N__30877;
    wire N__30876;
    wire N__30875;
    wire N__30874;
    wire N__30871;
    wire N__30868;
    wire N__30865;
    wire N__30864;
    wire N__30861;
    wire N__30854;
    wire N__30853;
    wire N__30852;
    wire N__30849;
    wire N__30848;
    wire N__30845;
    wire N__30842;
    wire N__30837;
    wire N__30834;
    wire N__30831;
    wire N__30830;
    wire N__30827;
    wire N__30824;
    wire N__30821;
    wire N__30816;
    wire N__30813;
    wire N__30802;
    wire N__30799;
    wire N__30796;
    wire N__30793;
    wire N__30790;
    wire N__30787;
    wire N__30784;
    wire N__30781;
    wire N__30780;
    wire N__30779;
    wire N__30776;
    wire N__30771;
    wire N__30770;
    wire N__30769;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30761;
    wire N__30760;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30749;
    wire N__30744;
    wire N__30739;
    wire N__30736;
    wire N__30735;
    wire N__30730;
    wire N__30727;
    wire N__30724;
    wire N__30721;
    wire N__30716;
    wire N__30713;
    wire N__30710;
    wire N__30697;
    wire N__30696;
    wire N__30695;
    wire N__30694;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30683;
    wire N__30680;
    wire N__30679;
    wire N__30676;
    wire N__30669;
    wire N__30666;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30656;
    wire N__30653;
    wire N__30650;
    wire N__30649;
    wire N__30646;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30628;
    wire N__30619;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30604;
    wire N__30603;
    wire N__30598;
    wire N__30597;
    wire N__30594;
    wire N__30591;
    wire N__30588;
    wire N__30583;
    wire N__30580;
    wire N__30579;
    wire N__30576;
    wire N__30575;
    wire N__30572;
    wire N__30569;
    wire N__30566;
    wire N__30563;
    wire N__30556;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30543;
    wire N__30538;
    wire N__30535;
    wire N__30532;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30524;
    wire N__30523;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30513;
    wire N__30512;
    wire N__30509;
    wire N__30506;
    wire N__30505;
    wire N__30500;
    wire N__30497;
    wire N__30494;
    wire N__30489;
    wire N__30488;
    wire N__30487;
    wire N__30484;
    wire N__30479;
    wire N__30476;
    wire N__30473;
    wire N__30470;
    wire N__30467;
    wire N__30464;
    wire N__30461;
    wire N__30454;
    wire N__30451;
    wire N__30442;
    wire N__30441;
    wire N__30438;
    wire N__30437;
    wire N__30436;
    wire N__30435;
    wire N__30434;
    wire N__30431;
    wire N__30428;
    wire N__30423;
    wire N__30422;
    wire N__30421;
    wire N__30418;
    wire N__30415;
    wire N__30412;
    wire N__30407;
    wire N__30402;
    wire N__30397;
    wire N__30390;
    wire N__30387;
    wire N__30384;
    wire N__30379;
    wire N__30378;
    wire N__30377;
    wire N__30372;
    wire N__30371;
    wire N__30368;
    wire N__30365;
    wire N__30362;
    wire N__30359;
    wire N__30356;
    wire N__30349;
    wire N__30346;
    wire N__30343;
    wire N__30340;
    wire N__30339;
    wire N__30336;
    wire N__30335;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30323;
    wire N__30316;
    wire N__30315;
    wire N__30312;
    wire N__30309;
    wire N__30306;
    wire N__30305;
    wire N__30304;
    wire N__30301;
    wire N__30300;
    wire N__30299;
    wire N__30296;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30282;
    wire N__30271;
    wire N__30268;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30255;
    wire N__30252;
    wire N__30249;
    wire N__30244;
    wire N__30241;
    wire N__30238;
    wire N__30237;
    wire N__30234;
    wire N__30231;
    wire N__30228;
    wire N__30223;
    wire N__30220;
    wire N__30219;
    wire N__30216;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30204;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30192;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30182;
    wire N__30177;
    wire N__30172;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30142;
    wire N__30139;
    wire N__30136;
    wire N__30133;
    wire N__30130;
    wire N__30129;
    wire N__30126;
    wire N__30123;
    wire N__30118;
    wire N__30117;
    wire N__30114;
    wire N__30111;
    wire N__30110;
    wire N__30109;
    wire N__30104;
    wire N__30101;
    wire N__30098;
    wire N__30095;
    wire N__30088;
    wire N__30085;
    wire N__30084;
    wire N__30081;
    wire N__30078;
    wire N__30073;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30057;
    wire N__30056;
    wire N__30055;
    wire N__30052;
    wire N__30049;
    wire N__30044;
    wire N__30041;
    wire N__30034;
    wire N__30031;
    wire N__30028;
    wire N__30027;
    wire N__30026;
    wire N__30025;
    wire N__30022;
    wire N__30019;
    wire N__30018;
    wire N__30015;
    wire N__30012;
    wire N__30009;
    wire N__30006;
    wire N__30003;
    wire N__30000;
    wire N__29995;
    wire N__29992;
    wire N__29983;
    wire N__29982;
    wire N__29981;
    wire N__29978;
    wire N__29975;
    wire N__29974;
    wire N__29973;
    wire N__29972;
    wire N__29969;
    wire N__29968;
    wire N__29967;
    wire N__29966;
    wire N__29955;
    wire N__29954;
    wire N__29949;
    wire N__29946;
    wire N__29945;
    wire N__29942;
    wire N__29941;
    wire N__29938;
    wire N__29935;
    wire N__29930;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29920;
    wire N__29919;
    wire N__29918;
    wire N__29917;
    wire N__29912;
    wire N__29907;
    wire N__29904;
    wire N__29901;
    wire N__29898;
    wire N__29895;
    wire N__29894;
    wire N__29893;
    wire N__29890;
    wire N__29889;
    wire N__29886;
    wire N__29885;
    wire N__29884;
    wire N__29881;
    wire N__29878;
    wire N__29873;
    wire N__29868;
    wire N__29865;
    wire N__29862;
    wire N__29851;
    wire N__29836;
    wire N__29833;
    wire N__29830;
    wire N__29827;
    wire N__29824;
    wire N__29823;
    wire N__29820;
    wire N__29817;
    wire N__29816;
    wire N__29813;
    wire N__29810;
    wire N__29809;
    wire N__29806;
    wire N__29803;
    wire N__29800;
    wire N__29797;
    wire N__29788;
    wire N__29785;
    wire N__29782;
    wire N__29779;
    wire N__29776;
    wire N__29775;
    wire N__29772;
    wire N__29769;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29752;
    wire N__29749;
    wire N__29746;
    wire N__29745;
    wire N__29744;
    wire N__29743;
    wire N__29736;
    wire N__29735;
    wire N__29734;
    wire N__29733;
    wire N__29732;
    wire N__29729;
    wire N__29728;
    wire N__29727;
    wire N__29726;
    wire N__29723;
    wire N__29716;
    wire N__29713;
    wire N__29712;
    wire N__29711;
    wire N__29710;
    wire N__29709;
    wire N__29708;
    wire N__29707;
    wire N__29706;
    wire N__29705;
    wire N__29702;
    wire N__29695;
    wire N__29690;
    wire N__29685;
    wire N__29684;
    wire N__29681;
    wire N__29680;
    wire N__29679;
    wire N__29672;
    wire N__29669;
    wire N__29666;
    wire N__29665;
    wire N__29662;
    wire N__29661;
    wire N__29660;
    wire N__29659;
    wire N__29658;
    wire N__29657;
    wire N__29656;
    wire N__29653;
    wire N__29650;
    wire N__29649;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29633;
    wire N__29630;
    wire N__29619;
    wire N__29608;
    wire N__29603;
    wire N__29598;
    wire N__29581;
    wire N__29578;
    wire N__29575;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29560;
    wire N__29557;
    wire N__29554;
    wire N__29551;
    wire N__29548;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29536;
    wire N__29533;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29520;
    wire N__29517;
    wire N__29514;
    wire N__29509;
    wire N__29506;
    wire N__29505;
    wire N__29504;
    wire N__29503;
    wire N__29500;
    wire N__29493;
    wire N__29490;
    wire N__29485;
    wire N__29482;
    wire N__29479;
    wire N__29476;
    wire N__29475;
    wire N__29474;
    wire N__29473;
    wire N__29472;
    wire N__29469;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29455;
    wire N__29452;
    wire N__29449;
    wire N__29444;
    wire N__29439;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29427;
    wire N__29422;
    wire N__29419;
    wire N__29416;
    wire N__29413;
    wire N__29410;
    wire N__29407;
    wire N__29404;
    wire N__29401;
    wire N__29398;
    wire N__29395;
    wire N__29392;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29380;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29361;
    wire N__29358;
    wire N__29355;
    wire N__29352;
    wire N__29347;
    wire N__29344;
    wire N__29343;
    wire N__29342;
    wire N__29341;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29327;
    wire N__29326;
    wire N__29325;
    wire N__29322;
    wire N__29321;
    wire N__29320;
    wire N__29315;
    wire N__29310;
    wire N__29307;
    wire N__29302;
    wire N__29299;
    wire N__29296;
    wire N__29293;
    wire N__29288;
    wire N__29275;
    wire N__29272;
    wire N__29269;
    wire N__29266;
    wire N__29263;
    wire N__29260;
    wire N__29257;
    wire N__29256;
    wire N__29255;
    wire N__29252;
    wire N__29249;
    wire N__29244;
    wire N__29239;
    wire N__29236;
    wire N__29233;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29221;
    wire N__29218;
    wire N__29215;
    wire N__29212;
    wire N__29209;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29197;
    wire N__29194;
    wire N__29193;
    wire N__29188;
    wire N__29185;
    wire N__29184;
    wire N__29183;
    wire N__29182;
    wire N__29177;
    wire N__29172;
    wire N__29169;
    wire N__29166;
    wire N__29163;
    wire N__29160;
    wire N__29155;
    wire N__29152;
    wire N__29149;
    wire N__29146;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29134;
    wire N__29133;
    wire N__29132;
    wire N__29129;
    wire N__29126;
    wire N__29123;
    wire N__29116;
    wire N__29115;
    wire N__29114;
    wire N__29111;
    wire N__29106;
    wire N__29101;
    wire N__29098;
    wire N__29095;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29085;
    wire N__29082;
    wire N__29079;
    wire N__29076;
    wire N__29073;
    wire N__29070;
    wire N__29067;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29055;
    wire N__29052;
    wire N__29051;
    wire N__29050;
    wire N__29049;
    wire N__29046;
    wire N__29045;
    wire N__29042;
    wire N__29037;
    wire N__29036;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29022;
    wire N__29019;
    wire N__29014;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28993;
    wire N__28992;
    wire N__28989;
    wire N__28986;
    wire N__28983;
    wire N__28978;
    wire N__28977;
    wire N__28974;
    wire N__28971;
    wire N__28968;
    wire N__28965;
    wire N__28960;
    wire N__28957;
    wire N__28954;
    wire N__28953;
    wire N__28950;
    wire N__28947;
    wire N__28944;
    wire N__28939;
    wire N__28938;
    wire N__28935;
    wire N__28932;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28918;
    wire N__28915;
    wire N__28912;
    wire N__28909;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28894;
    wire N__28891;
    wire N__28888;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28876;
    wire N__28873;
    wire N__28872;
    wire N__28869;
    wire N__28866;
    wire N__28863;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28851;
    wire N__28848;
    wire N__28845;
    wire N__28842;
    wire N__28837;
    wire N__28834;
    wire N__28833;
    wire N__28828;
    wire N__28827;
    wire N__28824;
    wire N__28821;
    wire N__28816;
    wire N__28815;
    wire N__28812;
    wire N__28809;
    wire N__28804;
    wire N__28803;
    wire N__28802;
    wire N__28801;
    wire N__28800;
    wire N__28799;
    wire N__28798;
    wire N__28797;
    wire N__28796;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28785;
    wire N__28782;
    wire N__28779;
    wire N__28770;
    wire N__28765;
    wire N__28764;
    wire N__28763;
    wire N__28762;
    wire N__28761;
    wire N__28760;
    wire N__28755;
    wire N__28752;
    wire N__28747;
    wire N__28742;
    wire N__28739;
    wire N__28736;
    wire N__28729;
    wire N__28726;
    wire N__28723;
    wire N__28718;
    wire N__28705;
    wire N__28704;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28690;
    wire N__28689;
    wire N__28686;
    wire N__28683;
    wire N__28678;
    wire N__28677;
    wire N__28674;
    wire N__28671;
    wire N__28666;
    wire N__28663;
    wire N__28660;
    wire N__28657;
    wire N__28654;
    wire N__28651;
    wire N__28650;
    wire N__28649;
    wire N__28646;
    wire N__28645;
    wire N__28644;
    wire N__28643;
    wire N__28638;
    wire N__28635;
    wire N__28632;
    wire N__28627;
    wire N__28624;
    wire N__28615;
    wire N__28612;
    wire N__28611;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28591;
    wire N__28586;
    wire N__28579;
    wire N__28576;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28568;
    wire N__28565;
    wire N__28562;
    wire N__28561;
    wire N__28558;
    wire N__28555;
    wire N__28552;
    wire N__28549;
    wire N__28540;
    wire N__28537;
    wire N__28534;
    wire N__28531;
    wire N__28528;
    wire N__28525;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28514;
    wire N__28513;
    wire N__28510;
    wire N__28507;
    wire N__28502;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28486;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28467;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28453;
    wire N__28450;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28438;
    wire N__28435;
    wire N__28432;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28398;
    wire N__28397;
    wire N__28394;
    wire N__28393;
    wire N__28392;
    wire N__28389;
    wire N__28386;
    wire N__28383;
    wire N__28380;
    wire N__28377;
    wire N__28374;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28342;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28323;
    wire N__28322;
    wire N__28321;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28309;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28291;
    wire N__28290;
    wire N__28287;
    wire N__28284;
    wire N__28283;
    wire N__28282;
    wire N__28279;
    wire N__28274;
    wire N__28271;
    wire N__28268;
    wire N__28261;
    wire N__28258;
    wire N__28255;
    wire N__28254;
    wire N__28251;
    wire N__28250;
    wire N__28249;
    wire N__28246;
    wire N__28243;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28195;
    wire N__28192;
    wire N__28189;
    wire N__28186;
    wire N__28185;
    wire N__28184;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28169;
    wire N__28164;
    wire N__28161;
    wire N__28156;
    wire N__28153;
    wire N__28150;
    wire N__28147;
    wire N__28144;
    wire N__28141;
    wire N__28140;
    wire N__28139;
    wire N__28136;
    wire N__28133;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28120;
    wire N__28117;
    wire N__28114;
    wire N__28111;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28084;
    wire N__28083;
    wire N__28082;
    wire N__28081;
    wire N__28078;
    wire N__28075;
    wire N__28072;
    wire N__28069;
    wire N__28066;
    wire N__28063;
    wire N__28060;
    wire N__28057;
    wire N__28054;
    wire N__28049;
    wire N__28046;
    wire N__28043;
    wire N__28036;
    wire N__28033;
    wire N__28030;
    wire N__28029;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28017;
    wire N__28012;
    wire N__28009;
    wire N__28006;
    wire N__28003;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27991;
    wire N__27990;
    wire N__27987;
    wire N__27984;
    wire N__27983;
    wire N__27982;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27972;
    wire N__27969;
    wire N__27966;
    wire N__27963;
    wire N__27958;
    wire N__27955;
    wire N__27948;
    wire N__27943;
    wire N__27940;
    wire N__27939;
    wire N__27938;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27910;
    wire N__27907;
    wire N__27906;
    wire N__27903;
    wire N__27900;
    wire N__27897;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27880;
    wire N__27879;
    wire N__27878;
    wire N__27875;
    wire N__27872;
    wire N__27869;
    wire N__27866;
    wire N__27865;
    wire N__27864;
    wire N__27861;
    wire N__27856;
    wire N__27851;
    wire N__27848;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27828;
    wire N__27825;
    wire N__27824;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27808;
    wire N__27805;
    wire N__27804;
    wire N__27803;
    wire N__27802;
    wire N__27801;
    wire N__27800;
    wire N__27791;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27783;
    wire N__27782;
    wire N__27779;
    wire N__27776;
    wire N__27771;
    wire N__27770;
    wire N__27769;
    wire N__27768;
    wire N__27765;
    wire N__27764;
    wire N__27763;
    wire N__27762;
    wire N__27761;
    wire N__27758;
    wire N__27753;
    wire N__27750;
    wire N__27747;
    wire N__27746;
    wire N__27745;
    wire N__27744;
    wire N__27743;
    wire N__27742;
    wire N__27741;
    wire N__27736;
    wire N__27731;
    wire N__27724;
    wire N__27721;
    wire N__27714;
    wire N__27713;
    wire N__27712;
    wire N__27711;
    wire N__27710;
    wire N__27709;
    wire N__27708;
    wire N__27707;
    wire N__27706;
    wire N__27705;
    wire N__27704;
    wire N__27695;
    wire N__27690;
    wire N__27687;
    wire N__27680;
    wire N__27677;
    wire N__27674;
    wire N__27673;
    wire N__27672;
    wire N__27671;
    wire N__27666;
    wire N__27657;
    wire N__27650;
    wire N__27647;
    wire N__27644;
    wire N__27641;
    wire N__27636;
    wire N__27627;
    wire N__27610;
    wire N__27609;
    wire N__27608;
    wire N__27605;
    wire N__27600;
    wire N__27597;
    wire N__27596;
    wire N__27593;
    wire N__27590;
    wire N__27587;
    wire N__27584;
    wire N__27577;
    wire N__27576;
    wire N__27575;
    wire N__27574;
    wire N__27573;
    wire N__27570;
    wire N__27569;
    wire N__27568;
    wire N__27565;
    wire N__27560;
    wire N__27559;
    wire N__27558;
    wire N__27557;
    wire N__27556;
    wire N__27553;
    wire N__27552;
    wire N__27551;
    wire N__27550;
    wire N__27549;
    wire N__27548;
    wire N__27545;
    wire N__27540;
    wire N__27535;
    wire N__27534;
    wire N__27533;
    wire N__27532;
    wire N__27529;
    wire N__27520;
    wire N__27515;
    wire N__27510;
    wire N__27507;
    wire N__27500;
    wire N__27495;
    wire N__27492;
    wire N__27475;
    wire N__27472;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27464;
    wire N__27461;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27449;
    wire N__27446;
    wire N__27443;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27427;
    wire N__27426;
    wire N__27425;
    wire N__27422;
    wire N__27417;
    wire N__27412;
    wire N__27409;
    wire N__27406;
    wire N__27403;
    wire N__27402;
    wire N__27399;
    wire N__27396;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27379;
    wire N__27378;
    wire N__27377;
    wire N__27376;
    wire N__27375;
    wire N__27366;
    wire N__27363;
    wire N__27358;
    wire N__27357;
    wire N__27354;
    wire N__27353;
    wire N__27352;
    wire N__27349;
    wire N__27348;
    wire N__27347;
    wire N__27344;
    wire N__27339;
    wire N__27338;
    wire N__27335;
    wire N__27330;
    wire N__27325;
    wire N__27322;
    wire N__27313;
    wire N__27312;
    wire N__27311;
    wire N__27310;
    wire N__27309;
    wire N__27308;
    wire N__27303;
    wire N__27300;
    wire N__27297;
    wire N__27294;
    wire N__27291;
    wire N__27280;
    wire N__27277;
    wire N__27274;
    wire N__27271;
    wire N__27268;
    wire N__27265;
    wire N__27262;
    wire N__27259;
    wire N__27256;
    wire N__27253;
    wire N__27250;
    wire N__27249;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27231;
    wire N__27230;
    wire N__27229;
    wire N__27226;
    wire N__27223;
    wire N__27218;
    wire N__27215;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27189;
    wire N__27188;
    wire N__27185;
    wire N__27182;
    wire N__27179;
    wire N__27172;
    wire N__27171;
    wire N__27170;
    wire N__27169;
    wire N__27168;
    wire N__27165;
    wire N__27160;
    wire N__27155;
    wire N__27148;
    wire N__27147;
    wire N__27146;
    wire N__27145;
    wire N__27144;
    wire N__27143;
    wire N__27142;
    wire N__27135;
    wire N__27132;
    wire N__27125;
    wire N__27118;
    wire N__27117;
    wire N__27114;
    wire N__27111;
    wire N__27106;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27082;
    wire N__27079;
    wire N__27076;
    wire N__27073;
    wire N__27070;
    wire N__27067;
    wire N__27064;
    wire N__27061;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27049;
    wire N__27048;
    wire N__27043;
    wire N__27040;
    wire N__27039;
    wire N__27036;
    wire N__27033;
    wire N__27028;
    wire N__27027;
    wire N__27026;
    wire N__27021;
    wire N__27018;
    wire N__27013;
    wire N__27012;
    wire N__27009;
    wire N__27006;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26989;
    wire N__26986;
    wire N__26983;
    wire N__26980;
    wire N__26977;
    wire N__26974;
    wire N__26973;
    wire N__26970;
    wire N__26967;
    wire N__26962;
    wire N__26959;
    wire N__26958;
    wire N__26957;
    wire N__26954;
    wire N__26951;
    wire N__26948;
    wire N__26941;
    wire N__26940;
    wire N__26937;
    wire N__26936;
    wire N__26933;
    wire N__26932;
    wire N__26929;
    wire N__26926;
    wire N__26923;
    wire N__26920;
    wire N__26919;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26911;
    wire N__26910;
    wire N__26907;
    wire N__26902;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26881;
    wire N__26878;
    wire N__26875;
    wire N__26860;
    wire N__26859;
    wire N__26858;
    wire N__26853;
    wire N__26852;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26840;
    wire N__26833;
    wire N__26832;
    wire N__26831;
    wire N__26828;
    wire N__26825;
    wire N__26824;
    wire N__26821;
    wire N__26820;
    wire N__26817;
    wire N__26814;
    wire N__26811;
    wire N__26808;
    wire N__26805;
    wire N__26794;
    wire N__26793;
    wire N__26790;
    wire N__26785;
    wire N__26782;
    wire N__26781;
    wire N__26780;
    wire N__26775;
    wire N__26774;
    wire N__26773;
    wire N__26770;
    wire N__26767;
    wire N__26762;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26734;
    wire N__26733;
    wire N__26732;
    wire N__26729;
    wire N__26726;
    wire N__26725;
    wire N__26722;
    wire N__26719;
    wire N__26716;
    wire N__26713;
    wire N__26704;
    wire N__26703;
    wire N__26700;
    wire N__26699;
    wire N__26698;
    wire N__26695;
    wire N__26692;
    wire N__26689;
    wire N__26686;
    wire N__26679;
    wire N__26674;
    wire N__26671;
    wire N__26670;
    wire N__26669;
    wire N__26668;
    wire N__26665;
    wire N__26662;
    wire N__26657;
    wire N__26650;
    wire N__26649;
    wire N__26646;
    wire N__26645;
    wire N__26642;
    wire N__26639;
    wire N__26636;
    wire N__26635;
    wire N__26632;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26614;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26581;
    wire N__26578;
    wire N__26577;
    wire N__26574;
    wire N__26571;
    wire N__26568;
    wire N__26563;
    wire N__26562;
    wire N__26559;
    wire N__26556;
    wire N__26553;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26539;
    wire N__26538;
    wire N__26537;
    wire N__26536;
    wire N__26533;
    wire N__26532;
    wire N__26529;
    wire N__26526;
    wire N__26525;
    wire N__26522;
    wire N__26521;
    wire N__26520;
    wire N__26517;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26491;
    wire N__26490;
    wire N__26485;
    wire N__26482;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26462;
    wire N__26459;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26437;
    wire N__26436;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26428;
    wire N__26425;
    wire N__26422;
    wire N__26419;
    wire N__26416;
    wire N__26413;
    wire N__26410;
    wire N__26401;
    wire N__26398;
    wire N__26395;
    wire N__26392;
    wire N__26391;
    wire N__26390;
    wire N__26383;
    wire N__26382;
    wire N__26379;
    wire N__26378;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26356;
    wire N__26353;
    wire N__26350;
    wire N__26349;
    wire N__26346;
    wire N__26343;
    wire N__26340;
    wire N__26335;
    wire N__26332;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26322;
    wire N__26319;
    wire N__26316;
    wire N__26313;
    wire N__26308;
    wire N__26305;
    wire N__26304;
    wire N__26301;
    wire N__26298;
    wire N__26295;
    wire N__26290;
    wire N__26287;
    wire N__26286;
    wire N__26283;
    wire N__26280;
    wire N__26277;
    wire N__26272;
    wire N__26271;
    wire N__26268;
    wire N__26265;
    wire N__26262;
    wire N__26257;
    wire N__26254;
    wire N__26253;
    wire N__26250;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26242;
    wire N__26241;
    wire N__26238;
    wire N__26235;
    wire N__26232;
    wire N__26229;
    wire N__26226;
    wire N__26215;
    wire N__26212;
    wire N__26209;
    wire N__26208;
    wire N__26207;
    wire N__26204;
    wire N__26203;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26176;
    wire N__26175;
    wire N__26174;
    wire N__26173;
    wire N__26170;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26152;
    wire N__26151;
    wire N__26150;
    wire N__26145;
    wire N__26144;
    wire N__26141;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26131;
    wire N__26126;
    wire N__26123;
    wire N__26120;
    wire N__26117;
    wire N__26110;
    wire N__26109;
    wire N__26106;
    wire N__26103;
    wire N__26100;
    wire N__26097;
    wire N__26092;
    wire N__26091;
    wire N__26088;
    wire N__26085;
    wire N__26082;
    wire N__26077;
    wire N__26074;
    wire N__26071;
    wire N__26070;
    wire N__26067;
    wire N__26064;
    wire N__26061;
    wire N__26056;
    wire N__26053;
    wire N__26050;
    wire N__26049;
    wire N__26046;
    wire N__26043;
    wire N__26040;
    wire N__26035;
    wire N__26034;
    wire N__26031;
    wire N__26028;
    wire N__26023;
    wire N__26020;
    wire N__26017;
    wire N__26016;
    wire N__26013;
    wire N__26010;
    wire N__26007;
    wire N__26002;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25983;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25962;
    wire N__25959;
    wire N__25956;
    wire N__25951;
    wire N__25950;
    wire N__25949;
    wire N__25948;
    wire N__25945;
    wire N__25942;
    wire N__25937;
    wire N__25930;
    wire N__25929;
    wire N__25926;
    wire N__25925;
    wire N__25922;
    wire N__25919;
    wire N__25914;
    wire N__25909;
    wire N__25908;
    wire N__25905;
    wire N__25902;
    wire N__25899;
    wire N__25894;
    wire N__25891;
    wire N__25888;
    wire N__25887;
    wire N__25886;
    wire N__25883;
    wire N__25880;
    wire N__25879;
    wire N__25876;
    wire N__25871;
    wire N__25866;
    wire N__25861;
    wire N__25860;
    wire N__25855;
    wire N__25852;
    wire N__25851;
    wire N__25850;
    wire N__25847;
    wire N__25842;
    wire N__25837;
    wire N__25834;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25824;
    wire N__25819;
    wire N__25818;
    wire N__25817;
    wire N__25814;
    wire N__25809;
    wire N__25806;
    wire N__25801;
    wire N__25798;
    wire N__25795;
    wire N__25794;
    wire N__25791;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25774;
    wire N__25771;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25761;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25749;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25735;
    wire N__25732;
    wire N__25731;
    wire N__25728;
    wire N__25725;
    wire N__25724;
    wire N__25719;
    wire N__25716;
    wire N__25715;
    wire N__25714;
    wire N__25713;
    wire N__25712;
    wire N__25711;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25680;
    wire N__25675;
    wire N__25674;
    wire N__25673;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25665;
    wire N__25664;
    wire N__25661;
    wire N__25658;
    wire N__25653;
    wire N__25650;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25639;
    wire N__25638;
    wire N__25635;
    wire N__25630;
    wire N__25627;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25603;
    wire N__25602;
    wire N__25599;
    wire N__25596;
    wire N__25595;
    wire N__25594;
    wire N__25593;
    wire N__25590;
    wire N__25589;
    wire N__25586;
    wire N__25585;
    wire N__25582;
    wire N__25579;
    wire N__25576;
    wire N__25573;
    wire N__25570;
    wire N__25567;
    wire N__25564;
    wire N__25563;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25519;
    wire N__25516;
    wire N__25515;
    wire N__25514;
    wire N__25513;
    wire N__25510;
    wire N__25503;
    wire N__25498;
    wire N__25495;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25474;
    wire N__25471;
    wire N__25470;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25455;
    wire N__25452;
    wire N__25451;
    wire N__25446;
    wire N__25443;
    wire N__25438;
    wire N__25435;
    wire N__25432;
    wire N__25429;
    wire N__25426;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25414;
    wire N__25413;
    wire N__25412;
    wire N__25409;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25394;
    wire N__25387;
    wire N__25384;
    wire N__25381;
    wire N__25378;
    wire N__25375;
    wire N__25374;
    wire N__25373;
    wire N__25370;
    wire N__25367;
    wire N__25366;
    wire N__25363;
    wire N__25360;
    wire N__25357;
    wire N__25354;
    wire N__25345;
    wire N__25342;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25330;
    wire N__25329;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25314;
    wire N__25309;
    wire N__25306;
    wire N__25303;
    wire N__25300;
    wire N__25297;
    wire N__25294;
    wire N__25293;
    wire N__25292;
    wire N__25289;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25270;
    wire N__25267;
    wire N__25264;
    wire N__25261;
    wire N__25260;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25240;
    wire N__25237;
    wire N__25234;
    wire N__25231;
    wire N__25228;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25216;
    wire N__25213;
    wire N__25210;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25179;
    wire N__25176;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25168;
    wire N__25165;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25144;
    wire N__25141;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25123;
    wire N__25122;
    wire N__25121;
    wire N__25120;
    wire N__25117;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25096;
    wire N__25087;
    wire N__25086;
    wire N__25085;
    wire N__25084;
    wire N__25081;
    wire N__25080;
    wire N__25077;
    wire N__25074;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25066;
    wire N__25063;
    wire N__25062;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25045;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25029;
    wire N__25018;
    wire N__25017;
    wire N__25016;
    wire N__25013;
    wire N__25010;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24997;
    wire N__24994;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24975;
    wire N__24972;
    wire N__24967;
    wire N__24964;
    wire N__24961;
    wire N__24960;
    wire N__24957;
    wire N__24956;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24943;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24913;
    wire N__24910;
    wire N__24909;
    wire N__24908;
    wire N__24907;
    wire N__24904;
    wire N__24901;
    wire N__24898;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24886;
    wire N__24883;
    wire N__24880;
    wire N__24877;
    wire N__24868;
    wire N__24865;
    wire N__24864;
    wire N__24861;
    wire N__24860;
    wire N__24857;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24847;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24823;
    wire N__24822;
    wire N__24819;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24808;
    wire N__24805;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24789;
    wire N__24784;
    wire N__24781;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24761;
    wire N__24758;
    wire N__24755;
    wire N__24752;
    wire N__24751;
    wire N__24748;
    wire N__24743;
    wire N__24740;
    wire N__24735;
    wire N__24732;
    wire N__24727;
    wire N__24726;
    wire N__24723;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24712;
    wire N__24709;
    wire N__24704;
    wire N__24701;
    wire N__24698;
    wire N__24693;
    wire N__24688;
    wire N__24685;
    wire N__24682;
    wire N__24681;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24667;
    wire N__24664;
    wire N__24661;
    wire N__24658;
    wire N__24655;
    wire N__24652;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24625;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24615;
    wire N__24612;
    wire N__24609;
    wire N__24604;
    wire N__24603;
    wire N__24602;
    wire N__24601;
    wire N__24596;
    wire N__24593;
    wire N__24590;
    wire N__24587;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24562;
    wire N__24559;
    wire N__24556;
    wire N__24553;
    wire N__24550;
    wire N__24547;
    wire N__24546;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24535;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24516;
    wire N__24511;
    wire N__24510;
    wire N__24509;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24492;
    wire N__24491;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24479;
    wire N__24476;
    wire N__24475;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24454;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24446;
    wire N__24441;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24433;
    wire N__24430;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24420;
    wire N__24415;
    wire N__24412;
    wire N__24403;
    wire N__24402;
    wire N__24399;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24373;
    wire N__24368;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24352;
    wire N__24349;
    wire N__24348;
    wire N__24347;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24337;
    wire N__24334;
    wire N__24331;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24313;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24301;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24286;
    wire N__24283;
    wire N__24282;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24259;
    wire N__24256;
    wire N__24253;
    wire N__24250;
    wire N__24247;
    wire N__24244;
    wire N__24241;
    wire N__24238;
    wire N__24237;
    wire N__24232;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24183;
    wire N__24182;
    wire N__24179;
    wire N__24174;
    wire N__24173;
    wire N__24172;
    wire N__24171;
    wire N__24170;
    wire N__24169;
    wire N__24166;
    wire N__24163;
    wire N__24160;
    wire N__24157;
    wire N__24156;
    wire N__24153;
    wire N__24150;
    wire N__24147;
    wire N__24144;
    wire N__24139;
    wire N__24136;
    wire N__24131;
    wire N__24128;
    wire N__24115;
    wire N__24114;
    wire N__24113;
    wire N__24110;
    wire N__24105;
    wire N__24104;
    wire N__24103;
    wire N__24100;
    wire N__24097;
    wire N__24094;
    wire N__24091;
    wire N__24088;
    wire N__24083;
    wire N__24076;
    wire N__24075;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24067;
    wire N__24066;
    wire N__24065;
    wire N__24064;
    wire N__24063;
    wire N__24056;
    wire N__24053;
    wire N__24050;
    wire N__24049;
    wire N__24046;
    wire N__24045;
    wire N__24044;
    wire N__24043;
    wire N__24040;
    wire N__24039;
    wire N__24038;
    wire N__24035;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24023;
    wire N__24020;
    wire N__24015;
    wire N__24012;
    wire N__24007;
    wire N__24004;
    wire N__24001;
    wire N__23996;
    wire N__23991;
    wire N__23982;
    wire N__23971;
    wire N__23970;
    wire N__23969;
    wire N__23968;
    wire N__23965;
    wire N__23964;
    wire N__23963;
    wire N__23962;
    wire N__23961;
    wire N__23960;
    wire N__23959;
    wire N__23958;
    wire N__23957;
    wire N__23956;
    wire N__23955;
    wire N__23954;
    wire N__23953;
    wire N__23950;
    wire N__23945;
    wire N__23942;
    wire N__23937;
    wire N__23934;
    wire N__23933;
    wire N__23930;
    wire N__23925;
    wire N__23922;
    wire N__23919;
    wire N__23914;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23896;
    wire N__23893;
    wire N__23892;
    wire N__23879;
    wire N__23878;
    wire N__23877;
    wire N__23872;
    wire N__23869;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23844;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23811;
    wire N__23808;
    wire N__23805;
    wire N__23802;
    wire N__23797;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23785;
    wire N__23782;
    wire N__23781;
    wire N__23780;
    wire N__23775;
    wire N__23772;
    wire N__23767;
    wire N__23764;
    wire N__23763;
    wire N__23758;
    wire N__23755;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23745;
    wire N__23742;
    wire N__23739;
    wire N__23734;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23722;
    wire N__23721;
    wire N__23718;
    wire N__23715;
    wire N__23714;
    wire N__23709;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23695;
    wire N__23692;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23680;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23668;
    wire N__23665;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23655;
    wire N__23652;
    wire N__23649;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23629;
    wire N__23626;
    wire N__23625;
    wire N__23622;
    wire N__23619;
    wire N__23616;
    wire N__23611;
    wire N__23608;
    wire N__23607;
    wire N__23606;
    wire N__23605;
    wire N__23604;
    wire N__23601;
    wire N__23596;
    wire N__23591;
    wire N__23588;
    wire N__23581;
    wire N__23580;
    wire N__23577;
    wire N__23574;
    wire N__23573;
    wire N__23572;
    wire N__23569;
    wire N__23566;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23548;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23535;
    wire N__23532;
    wire N__23531;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23519;
    wire N__23512;
    wire N__23511;
    wire N__23508;
    wire N__23507;
    wire N__23504;
    wire N__23499;
    wire N__23494;
    wire N__23491;
    wire N__23488;
    wire N__23485;
    wire N__23484;
    wire N__23483;
    wire N__23480;
    wire N__23479;
    wire N__23476;
    wire N__23473;
    wire N__23470;
    wire N__23467;
    wire N__23464;
    wire N__23461;
    wire N__23458;
    wire N__23449;
    wire N__23446;
    wire N__23443;
    wire N__23440;
    wire N__23437;
    wire N__23434;
    wire N__23431;
    wire N__23430;
    wire N__23429;
    wire N__23428;
    wire N__23427;
    wire N__23426;
    wire N__23423;
    wire N__23422;
    wire N__23421;
    wire N__23420;
    wire N__23419;
    wire N__23418;
    wire N__23417;
    wire N__23416;
    wire N__23415;
    wire N__23410;
    wire N__23403;
    wire N__23402;
    wire N__23399;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23379;
    wire N__23378;
    wire N__23377;
    wire N__23376;
    wire N__23375;
    wire N__23374;
    wire N__23373;
    wire N__23372;
    wire N__23371;
    wire N__23370;
    wire N__23369;
    wire N__23368;
    wire N__23367;
    wire N__23366;
    wire N__23365;
    wire N__23364;
    wire N__23359;
    wire N__23358;
    wire N__23357;
    wire N__23356;
    wire N__23355;
    wire N__23354;
    wire N__23353;
    wire N__23352;
    wire N__23351;
    wire N__23348;
    wire N__23339;
    wire N__23336;
    wire N__23327;
    wire N__23312;
    wire N__23303;
    wire N__23300;
    wire N__23291;
    wire N__23282;
    wire N__23277;
    wire N__23260;
    wire N__23259;
    wire N__23258;
    wire N__23257;
    wire N__23256;
    wire N__23255;
    wire N__23254;
    wire N__23253;
    wire N__23246;
    wire N__23241;
    wire N__23240;
    wire N__23239;
    wire N__23238;
    wire N__23237;
    wire N__23236;
    wire N__23235;
    wire N__23234;
    wire N__23233;
    wire N__23226;
    wire N__23225;
    wire N__23224;
    wire N__23223;
    wire N__23218;
    wire N__23215;
    wire N__23206;
    wire N__23205;
    wire N__23204;
    wire N__23203;
    wire N__23202;
    wire N__23201;
    wire N__23200;
    wire N__23199;
    wire N__23198;
    wire N__23197;
    wire N__23196;
    wire N__23195;
    wire N__23192;
    wire N__23191;
    wire N__23190;
    wire N__23189;
    wire N__23188;
    wire N__23187;
    wire N__23186;
    wire N__23185;
    wire N__23184;
    wire N__23183;
    wire N__23182;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23157;
    wire N__23148;
    wire N__23133;
    wire N__23124;
    wire N__23113;
    wire N__23108;
    wire N__23103;
    wire N__23098;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23064;
    wire N__23063;
    wire N__23062;
    wire N__23061;
    wire N__23060;
    wire N__23059;
    wire N__23058;
    wire N__23057;
    wire N__23056;
    wire N__23053;
    wire N__23050;
    wire N__23049;
    wire N__23048;
    wire N__23047;
    wire N__23046;
    wire N__23045;
    wire N__23044;
    wire N__23043;
    wire N__23042;
    wire N__23041;
    wire N__23040;
    wire N__23039;
    wire N__23038;
    wire N__23037;
    wire N__23036;
    wire N__23035;
    wire N__23022;
    wire N__23017;
    wire N__23016;
    wire N__23009;
    wire N__23008;
    wire N__23007;
    wire N__23006;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22996;
    wire N__22995;
    wire N__22994;
    wire N__22993;
    wire N__22992;
    wire N__22991;
    wire N__22990;
    wire N__22989;
    wire N__22988;
    wire N__22983;
    wire N__22980;
    wire N__22979;
    wire N__22978;
    wire N__22977;
    wire N__22976;
    wire N__22975;
    wire N__22972;
    wire N__22971;
    wire N__22966;
    wire N__22955;
    wire N__22954;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22928;
    wire N__22927;
    wire N__22926;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22905;
    wire N__22904;
    wire N__22903;
    wire N__22902;
    wire N__22901;
    wire N__22900;
    wire N__22899;
    wire N__22898;
    wire N__22897;
    wire N__22896;
    wire N__22895;
    wire N__22892;
    wire N__22891;
    wire N__22888;
    wire N__22887;
    wire N__22886;
    wire N__22881;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22856;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22844;
    wire N__22829;
    wire N__22814;
    wire N__22799;
    wire N__22788;
    wire N__22779;
    wire N__22772;
    wire N__22753;
    wire N__22752;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22726;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22708;
    wire N__22707;
    wire N__22706;
    wire N__22705;
    wire N__22704;
    wire N__22703;
    wire N__22702;
    wire N__22701;
    wire N__22700;
    wire N__22699;
    wire N__22698;
    wire N__22697;
    wire N__22696;
    wire N__22695;
    wire N__22694;
    wire N__22693;
    wire N__22692;
    wire N__22691;
    wire N__22690;
    wire N__22683;
    wire N__22676;
    wire N__22675;
    wire N__22674;
    wire N__22673;
    wire N__22672;
    wire N__22669;
    wire N__22668;
    wire N__22667;
    wire N__22666;
    wire N__22665;
    wire N__22662;
    wire N__22659;
    wire N__22652;
    wire N__22641;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22604;
    wire N__22599;
    wire N__22594;
    wire N__22587;
    wire N__22576;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22563;
    wire N__22560;
    wire N__22557;
    wire N__22554;
    wire N__22551;
    wire N__22548;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22500;
    wire N__22497;
    wire N__22496;
    wire N__22495;
    wire N__22494;
    wire N__22493;
    wire N__22492;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22442;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22425;
    wire N__22422;
    wire N__22419;
    wire N__22418;
    wire N__22413;
    wire N__22410;
    wire N__22409;
    wire N__22408;
    wire N__22405;
    wire N__22400;
    wire N__22397;
    wire N__22392;
    wire N__22387;
    wire N__22384;
    wire N__22383;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22371;
    wire N__22368;
    wire N__22365;
    wire N__22362;
    wire N__22359;
    wire N__22354;
    wire N__22353;
    wire N__22350;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22332;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22318;
    wire N__22315;
    wire N__22312;
    wire N__22309;
    wire N__22306;
    wire N__22303;
    wire N__22300;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22288;
    wire N__22287;
    wire N__22284;
    wire N__22281;
    wire N__22280;
    wire N__22279;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22261;
    wire N__22258;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22206;
    wire N__22205;
    wire N__22200;
    wire N__22197;
    wire N__22194;
    wire N__22191;
    wire N__22188;
    wire N__22183;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22164;
    wire N__22163;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22153;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22110;
    wire N__22107;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22099;
    wire N__22096;
    wire N__22091;
    wire N__22088;
    wire N__22081;
    wire N__22078;
    wire N__22077;
    wire N__22074;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22057;
    wire N__22054;
    wire N__22053;
    wire N__22050;
    wire N__22049;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22037;
    wire N__22030;
    wire N__22027;
    wire N__22024;
    wire N__22021;
    wire N__22020;
    wire N__22019;
    wire N__22016;
    wire N__22015;
    wire N__22010;
    wire N__22009;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__21999;
    wire N__21994;
    wire N__21985;
    wire N__21982;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21961;
    wire N__21958;
    wire N__21955;
    wire N__21952;
    wire N__21949;
    wire N__21948;
    wire N__21945;
    wire N__21942;
    wire N__21939;
    wire N__21936;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21907;
    wire N__21906;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21886;
    wire N__21885;
    wire N__21884;
    wire N__21881;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21856;
    wire N__21855;
    wire N__21852;
    wire N__21851;
    wire N__21848;
    wire N__21847;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21811;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21786;
    wire N__21785;
    wire N__21778;
    wire N__21775;
    wire N__21774;
    wire N__21771;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21754;
    wire N__21753;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21738;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21711;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21688;
    wire N__21687;
    wire N__21686;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21658;
    wire N__21657;
    wire N__21654;
    wire N__21653;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21642;
    wire N__21641;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21633;
    wire N__21628;
    wire N__21625;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21607;
    wire N__21602;
    wire N__21597;
    wire N__21594;
    wire N__21591;
    wire N__21588;
    wire N__21583;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21567;
    wire N__21564;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21547;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21519;
    wire N__21518;
    wire N__21515;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21488;
    wire N__21485;
    wire N__21480;
    wire N__21477;
    wire N__21472;
    wire N__21471;
    wire N__21470;
    wire N__21467;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21445;
    wire N__21442;
    wire N__21439;
    wire N__21436;
    wire N__21433;
    wire N__21426;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21387;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21367;
    wire N__21364;
    wire N__21363;
    wire N__21360;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21328;
    wire N__21327;
    wire N__21326;
    wire N__21323;
    wire N__21318;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21295;
    wire N__21292;
    wire N__21291;
    wire N__21290;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21259;
    wire N__21256;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21238;
    wire N__21235;
    wire N__21234;
    wire N__21233;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21220;
    wire N__21217;
    wire N__21212;
    wire N__21209;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21187;
    wire N__21184;
    wire N__21181;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21169;
    wire N__21168;
    wire N__21167;
    wire N__21164;
    wire N__21159;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21129;
    wire N__21128;
    wire N__21127;
    wire N__21124;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21106;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21096;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21076;
    wire N__21073;
    wire N__21070;
    wire N__21067;
    wire N__21066;
    wire N__21065;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21055;
    wire N__21052;
    wire N__21043;
    wire N__21040;
    wire N__21037;
    wire N__21034;
    wire N__21031;
    wire N__21028;
    wire N__21025;
    wire N__21022;
    wire N__21019;
    wire N__21018;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21001;
    wire N__20998;
    wire N__20995;
    wire N__20992;
    wire N__20989;
    wire N__20988;
    wire N__20987;
    wire N__20986;
    wire N__20985;
    wire N__20984;
    wire N__20983;
    wire N__20982;
    wire N__20981;
    wire N__20980;
    wire N__20979;
    wire N__20978;
    wire N__20977;
    wire N__20976;
    wire N__20971;
    wire N__20964;
    wire N__20957;
    wire N__20944;
    wire N__20935;
    wire N__20932;
    wire N__20929;
    wire N__20928;
    wire N__20925;
    wire N__20924;
    wire N__20923;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20911;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20893;
    wire N__20890;
    wire N__20887;
    wire N__20884;
    wire N__20881;
    wire N__20878;
    wire N__20877;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20860;
    wire N__20857;
    wire N__20854;
    wire N__20851;
    wire N__20850;
    wire N__20849;
    wire N__20848;
    wire N__20847;
    wire N__20846;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20830;
    wire N__20827;
    wire N__20818;
    wire N__20815;
    wire N__20812;
    wire N__20811;
    wire N__20810;
    wire N__20809;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20783;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20763;
    wire N__20762;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20750;
    wire N__20747;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20718;
    wire N__20715;
    wire N__20712;
    wire N__20709;
    wire N__20706;
    wire N__20701;
    wire N__20698;
    wire N__20697;
    wire N__20694;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20686;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20671;
    wire N__20662;
    wire N__20659;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20647;
    wire N__20646;
    wire N__20641;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20629;
    wire N__20626;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20614;
    wire N__20611;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20599;
    wire N__20596;
    wire N__20595;
    wire N__20594;
    wire N__20591;
    wire N__20586;
    wire N__20581;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20563;
    wire N__20562;
    wire N__20559;
    wire N__20556;
    wire N__20553;
    wire N__20550;
    wire N__20547;
    wire N__20544;
    wire N__20539;
    wire N__20536;
    wire N__20535;
    wire N__20532;
    wire N__20529;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20512;
    wire N__20509;
    wire N__20508;
    wire N__20507;
    wire N__20504;
    wire N__20499;
    wire N__20496;
    wire N__20493;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20434;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20368;
    wire N__20365;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20332;
    wire N__20329;
    wire N__20326;
    wire N__20323;
    wire N__20320;
    wire N__20317;
    wire N__20314;
    wire N__20311;
    wire N__20308;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20296;
    wire N__20293;
    wire N__20290;
    wire N__20287;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20275;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20260;
    wire N__20257;
    wire N__20254;
    wire N__20251;
    wire N__20248;
    wire N__20245;
    wire N__20242;
    wire N__20239;
    wire N__20236;
    wire N__20233;
    wire N__20230;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20215;
    wire N__20212;
    wire N__20209;
    wire N__20206;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20194;
    wire N__20191;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20176;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20147;
    wire N__20142;
    wire N__20141;
    wire N__20140;
    wire N__20139;
    wire N__20138;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20101;
    wire N__20100;
    wire N__20097;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20074;
    wire N__20073;
    wire N__20072;
    wire N__20069;
    wire N__20064;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20052;
    wire N__20049;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20032;
    wire N__20029;
    wire N__20026;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20004;
    wire N__20003;
    wire N__20002;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19990;
    wire N__19987;
    wire N__19984;
    wire N__19975;
    wire N__19972;
    wire N__19971;
    wire N__19970;
    wire N__19969;
    wire N__19966;
    wire N__19963;
    wire N__19962;
    wire N__19961;
    wire N__19958;
    wire N__19957;
    wire N__19954;
    wire N__19949;
    wire N__19946;
    wire N__19941;
    wire N__19936;
    wire N__19927;
    wire N__19926;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19918;
    wire N__19917;
    wire N__19914;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19896;
    wire N__19893;
    wire N__19890;
    wire N__19885;
    wire N__19882;
    wire N__19873;
    wire N__19872;
    wire N__19869;
    wire N__19866;
    wire N__19865;
    wire N__19864;
    wire N__19863;
    wire N__19860;
    wire N__19855;
    wire N__19852;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19834;
    wire N__19831;
    wire N__19828;
    wire N__19827;
    wire N__19826;
    wire N__19825;
    wire N__19824;
    wire N__19821;
    wire N__19816;
    wire N__19811;
    wire N__19804;
    wire N__19803;
    wire N__19802;
    wire N__19797;
    wire N__19794;
    wire N__19793;
    wire N__19792;
    wire N__19787;
    wire N__19782;
    wire N__19779;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19756;
    wire N__19753;
    wire N__19752;
    wire N__19749;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19732;
    wire N__19729;
    wire N__19726;
    wire N__19723;
    wire N__19722;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19680;
    wire N__19679;
    wire N__19678;
    wire N__19673;
    wire N__19672;
    wire N__19669;
    wire N__19666;
    wire N__19663;
    wire N__19660;
    wire N__19659;
    wire N__19656;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19612;
    wire N__19611;
    wire N__19610;
    wire N__19603;
    wire N__19600;
    wire N__19599;
    wire N__19598;
    wire N__19597;
    wire N__19592;
    wire N__19587;
    wire N__19582;
    wire N__19579;
    wire N__19576;
    wire N__19573;
    wire N__19570;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19548;
    wire N__19543;
    wire N__19542;
    wire N__19541;
    wire N__19540;
    wire N__19537;
    wire N__19532;
    wire N__19529;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19476;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19459;
    wire N__19456;
    wire N__19455;
    wire N__19454;
    wire N__19453;
    wire N__19452;
    wire N__19451;
    wire N__19450;
    wire N__19449;
    wire N__19448;
    wire N__19447;
    wire N__19446;
    wire N__19445;
    wire N__19444;
    wire N__19443;
    wire N__19442;
    wire N__19441;
    wire N__19440;
    wire N__19439;
    wire N__19438;
    wire N__19437;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19413;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19403;
    wire N__19402;
    wire N__19399;
    wire N__19398;
    wire N__19395;
    wire N__19394;
    wire N__19391;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19383;
    wire N__19380;
    wire N__19379;
    wire N__19376;
    wire N__19375;
    wire N__19372;
    wire N__19371;
    wire N__19368;
    wire N__19365;
    wire N__19362;
    wire N__19355;
    wire N__19344;
    wire N__19333;
    wire N__19316;
    wire N__19299;
    wire N__19292;
    wire N__19287;
    wire N__19280;
    wire N__19273;
    wire N__19272;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19252;
    wire N__19251;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19241;
    wire N__19238;
    wire N__19233;
    wire N__19228;
    wire N__19225;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19201;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19183;
    wire N__19180;
    wire N__19177;
    wire N__19174;
    wire N__19171;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19144;
    wire N__19141;
    wire N__19138;
    wire N__19135;
    wire N__19132;
    wire N__19129;
    wire N__19126;
    wire N__19123;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19069;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19057;
    wire N__19054;
    wire N__19051;
    wire N__19048;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19009;
    wire N__19006;
    wire N__19003;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18943;
    wire N__18940;
    wire N__18937;
    wire N__18934;
    wire N__18931;
    wire N__18928;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18916;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18898;
    wire N__18895;
    wire N__18892;
    wire N__18889;
    wire N__18886;
    wire N__18883;
    wire N__18880;
    wire N__18877;
    wire N__18874;
    wire N__18871;
    wire N__18868;
    wire N__18865;
    wire N__18862;
    wire N__18859;
    wire N__18856;
    wire N__18853;
    wire N__18850;
    wire N__18847;
    wire N__18844;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18832;
    wire N__18829;
    wire N__18826;
    wire N__18823;
    wire N__18820;
    wire N__18817;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18799;
    wire N__18796;
    wire N__18793;
    wire N__18790;
    wire N__18787;
    wire N__18784;
    wire N__18781;
    wire N__18778;
    wire N__18775;
    wire N__18772;
    wire N__18771;
    wire N__18770;
    wire N__18769;
    wire N__18766;
    wire N__18763;
    wire N__18758;
    wire N__18757;
    wire N__18756;
    wire N__18753;
    wire N__18748;
    wire N__18747;
    wire N__18744;
    wire N__18741;
    wire N__18736;
    wire N__18733;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18717;
    wire N__18714;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18694;
    wire N__18691;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18675;
    wire N__18672;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18655;
    wire N__18652;
    wire N__18649;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18630;
    wire N__18627;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18595;
    wire N__18592;
    wire N__18589;
    wire N__18588;
    wire N__18587;
    wire N__18584;
    wire N__18579;
    wire N__18574;
    wire N__18573;
    wire N__18572;
    wire N__18569;
    wire N__18564;
    wire N__18561;
    wire N__18558;
    wire N__18553;
    wire N__18552;
    wire N__18551;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18539;
    wire N__18534;
    wire N__18531;
    wire N__18528;
    wire N__18525;
    wire N__18520;
    wire N__18519;
    wire N__18516;
    wire N__18513;
    wire N__18508;
    wire N__18505;
    wire N__18502;
    wire N__18499;
    wire N__18498;
    wire N__18497;
    wire N__18494;
    wire N__18489;
    wire N__18486;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18472;
    wire N__18471;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18454;
    wire N__18451;
    wire N__18450;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18432;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18420;
    wire N__18417;
    wire N__18414;
    wire N__18413;
    wire N__18412;
    wire N__18409;
    wire N__18406;
    wire N__18403;
    wire N__18400;
    wire N__18397;
    wire N__18392;
    wire N__18389;
    wire N__18382;
    wire N__18379;
    wire N__18378;
    wire N__18375;
    wire N__18372;
    wire N__18367;
    wire N__18366;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18349;
    wire N__18348;
    wire N__18343;
    wire N__18340;
    wire N__18337;
    wire N__18334;
    wire N__18331;
    wire N__18328;
    wire N__18325;
    wire N__18322;
    wire N__18319;
    wire N__18316;
    wire N__18313;
    wire N__18310;
    wire N__18307;
    wire N__18304;
    wire N__18301;
    wire N__18298;
    wire N__18295;
    wire N__18292;
    wire N__18289;
    wire N__18286;
    wire N__18283;
    wire N__18280;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18259;
    wire N__18256;
    wire N__18253;
    wire N__18250;
    wire N__18247;
    wire N__18244;
    wire N__18241;
    wire N__18238;
    wire N__18235;
    wire N__18232;
    wire N__18229;
    wire N__18226;
    wire N__18223;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18213;
    wire N__18212;
    wire N__18211;
    wire N__18210;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18192;
    wire N__18181;
    wire N__18180;
    wire N__18179;
    wire N__18178;
    wire N__18177;
    wire N__18176;
    wire N__18175;
    wire N__18174;
    wire N__18167;
    wire N__18156;
    wire N__18151;
    wire N__18148;
    wire N__18145;
    wire N__18142;
    wire N__18141;
    wire N__18140;
    wire N__18137;
    wire N__18132;
    wire N__18127;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18112;
    wire N__18109;
    wire N__18106;
    wire N__18103;
    wire N__18100;
    wire N__18099;
    wire N__18098;
    wire N__18097;
    wire N__18096;
    wire N__18095;
    wire N__18088;
    wire N__18081;
    wire N__18076;
    wire N__18073;
    wire N__18070;
    wire N__18069;
    wire N__18066;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18056;
    wire N__18049;
    wire N__18046;
    wire N__18043;
    wire N__18040;
    wire N__18037;
    wire N__18034;
    wire N__18031;
    wire N__18028;
    wire N__18025;
    wire N__18022;
    wire N__18019;
    wire N__18016;
    wire N__18013;
    wire N__18010;
    wire N__18009;
    wire N__18008;
    wire N__18005;
    wire N__18000;
    wire N__17995;
    wire N__17994;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17982;
    wire N__17977;
    wire N__17976;
    wire N__17975;
    wire N__17972;
    wire N__17967;
    wire N__17962;
    wire N__17961;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17944;
    wire N__17941;
    wire N__17940;
    wire N__17939;
    wire N__17938;
    wire N__17935;
    wire N__17928;
    wire N__17923;
    wire N__17920;
    wire N__17917;
    wire N__17914;
    wire N__17911;
    wire N__17910;
    wire N__17909;
    wire N__17908;
    wire N__17907;
    wire N__17906;
    wire N__17899;
    wire N__17892;
    wire N__17887;
    wire N__17886;
    wire N__17885;
    wire N__17882;
    wire N__17877;
    wire N__17872;
    wire N__17871;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17854;
    wire N__17851;
    wire N__17850;
    wire N__17849;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17833;
    wire N__17830;
    wire N__17827;
    wire N__17824;
    wire N__17823;
    wire N__17820;
    wire N__17817;
    wire N__17812;
    wire N__17809;
    wire N__17806;
    wire N__17805;
    wire N__17804;
    wire N__17803;
    wire N__17802;
    wire N__17799;
    wire N__17796;
    wire N__17789;
    wire N__17782;
    wire N__17781;
    wire N__17780;
    wire N__17779;
    wire N__17778;
    wire N__17773;
    wire N__17766;
    wire N__17761;
    wire N__17760;
    wire N__17757;
    wire N__17754;
    wire N__17749;
    wire N__17748;
    wire N__17745;
    wire N__17744;
    wire N__17739;
    wire N__17736;
    wire N__17731;
    wire N__17728;
    wire N__17725;
    wire N__17724;
    wire N__17723;
    wire N__17718;
    wire N__17715;
    wire N__17710;
    wire N__17707;
    wire N__17704;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17692;
    wire N__17689;
    wire N__17686;
    wire N__17683;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17673;
    wire N__17672;
    wire N__17669;
    wire N__17664;
    wire N__17659;
    wire N__17658;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17641;
    wire N__17638;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17605;
    wire N__17602;
    wire N__17599;
    wire N__17596;
    wire N__17593;
    wire N__17590;
    wire N__17587;
    wire N__17584;
    wire N__17583;
    wire N__17578;
    wire N__17577;
    wire N__17574;
    wire N__17571;
    wire N__17566;
    wire N__17563;
    wire N__17562;
    wire N__17561;
    wire N__17556;
    wire N__17553;
    wire N__17548;
    wire N__17545;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17533;
    wire N__17530;
    wire N__17527;
    wire N__17524;
    wire N__17521;
    wire N__17518;
    wire N__17515;
    wire N__17512;
    wire N__17509;
    wire N__17506;
    wire N__17503;
    wire N__17500;
    wire N__17497;
    wire N__17494;
    wire N__17491;
    wire N__17488;
    wire N__17485;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17473;
    wire N__17470;
    wire N__17467;
    wire N__17464;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17440;
    wire N__17437;
    wire N__17434;
    wire N__17431;
    wire N__17428;
    wire N__17425;
    wire N__17422;
    wire N__17419;
    wire N__17416;
    wire N__17413;
    wire N__17412;
    wire N__17411;
    wire N__17404;
    wire N__17401;
    wire N__17398;
    wire N__17395;
    wire N__17392;
    wire N__17391;
    wire N__17390;
    wire N__17387;
    wire N__17382;
    wire N__17377;
    wire N__17374;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17362;
    wire N__17361;
    wire N__17358;
    wire N__17353;
    wire N__17352;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17338;
    wire N__17335;
    wire N__17332;
    wire N__17329;
    wire N__17326;
    wire N__17323;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17311;
    wire N__17308;
    wire N__17305;
    wire N__17302;
    wire N__17301;
    wire N__17296;
    wire N__17293;
    wire N__17290;
    wire N__17287;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17251;
    wire N__17248;
    wire N__17247;
    wire N__17246;
    wire N__17243;
    wire N__17240;
    wire N__17237;
    wire N__17230;
    wire N__17227;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17212;
    wire N__17209;
    wire N__17206;
    wire N__17203;
    wire N__17200;
    wire N__17197;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17185;
    wire N__17182;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17161;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire n17299_cascade_;
    wire LED_c;
    wire tx2_enable;
    wire n17298;
    wire bfn_1_28_0_;
    wire \c0.tx2.n15675 ;
    wire \c0.tx2.n15676 ;
    wire n17457;
    wire \c0.tx2.n15677 ;
    wire \c0.tx2.n15678 ;
    wire \c0.tx2.n15679 ;
    wire \c0.tx2.n15680 ;
    wire \c0.tx2.n15681 ;
    wire \c0.tx2.n15682 ;
    wire bfn_1_29_0_;
    wire n17640;
    wire n16824;
    wire n10_adj_2412;
    wire n17458;
    wire bfn_1_30_0_;
    wire \c0.tx.n15660 ;
    wire \c0.tx.n15661 ;
    wire \c0.tx.n15662 ;
    wire \c0.tx.n15663 ;
    wire \c0.tx.n15664 ;
    wire \c0.tx.n15665 ;
    wire \c0.tx.n15666 ;
    wire \c0.tx.n15667 ;
    wire bfn_1_31_0_;
    wire n17537_cascade_;
    wire \c0.rx.r_SM_Main_2_N_2090_2_cascade_ ;
    wire n17631;
    wire n16810_cascade_;
    wire \c0.rx.n13452_cascade_ ;
    wire n16867;
    wire n17222;
    wire \c0.rx.n16850 ;
    wire \c0.FRAME_MATCHER_state_7 ;
    wire \c0.n16443 ;
    wire \c0.FRAME_MATCHER_state_13 ;
    wire \c0.n16447 ;
    wire \c0.FRAME_MATCHER_state_11 ;
    wire \c0.n16451 ;
    wire \c0.n16445 ;
    wire n26;
    wire bfn_2_25_0_;
    wire n25;
    wire n15590;
    wire n24;
    wire n15591;
    wire n23;
    wire n15592;
    wire n22;
    wire n15593;
    wire n21;
    wire n15594;
    wire n20;
    wire n15595;
    wire n19;
    wire n15596;
    wire n15597;
    wire n18;
    wire bfn_2_26_0_;
    wire n17_adj_2422;
    wire n15598;
    wire n16;
    wire n15599;
    wire n15;
    wire n15600;
    wire n14_adj_2424;
    wire n15601;
    wire n13;
    wire n15602;
    wire n12_adj_2419;
    wire n15603;
    wire n11;
    wire n15604;
    wire n15605;
    wire n10_adj_2420;
    wire bfn_2_27_0_;
    wire n9;
    wire n15606;
    wire n8;
    wire n15607;
    wire n7;
    wire n15608;
    wire n6_adj_2421;
    wire n15609;
    wire blink_counter_21;
    wire n15610;
    wire blink_counter_22;
    wire n15611;
    wire blink_counter_23;
    wire n15612;
    wire n15613;
    wire blink_counter_24;
    wire bfn_2_28_0_;
    wire n15614;
    wire blink_counter_25;
    wire n17570;
    wire n17629;
    wire n17504;
    wire r_Clock_Count_2_adj_2452;
    wire r_Clock_Count_3_adj_2451;
    wire n9403;
    wire n17140_cascade_;
    wire n16817;
    wire n12_adj_2410;
    wire r_Clock_Count_5_adj_2449;
    wire r_Clock_Count_1_adj_2453;
    wire \c0.tx2.n10 ;
    wire n15837;
    wire n15837_cascade_;
    wire r_SM_Main_2_N_2033_1_cascade_;
    wire r_Clock_Count_7_adj_2447;
    wire r_Clock_Count_8_adj_2446;
    wire n9929;
    wire n17494;
    wire n17542;
    wire n17484;
    wire n17_adj_2416_cascade_;
    wire r_Clock_Count_2;
    wire r_Clock_Count_3;
    wire r_Clock_Count_0;
    wire r_Clock_Count_5;
    wire \c0.tx.n10_cascade_ ;
    wire n16863;
    wire n16863_cascade_;
    wire \c0.rx.r_SM_Main_2_N_2096_0_cascade_ ;
    wire n6_adj_2461;
    wire n17641;
    wire n17144_cascade_;
    wire n16828;
    wire bfn_2_32_0_;
    wire \c0.rx.n15668 ;
    wire r_Clock_Count_2_adj_2435;
    wire n16860;
    wire \c0.rx.n15669 ;
    wire \c0.rx.n15670 ;
    wire n16854;
    wire \c0.rx.n15671 ;
    wire \c0.rx.n15672 ;
    wire \c0.rx.n15673 ;
    wire r_Clock_Count_7_adj_2430;
    wire n16852;
    wire \c0.rx.n15674 ;
    wire n16855;
    wire \c0.FRAME_MATCHER_state_15 ;
    wire \c0.n16349 ;
    wire n1651_cascade_;
    wire n1651;
    wire n6_cascade_;
    wire n4;
    wire n8_adj_2459_cascade_;
    wire FRAME_MATCHER_state_31_N_1440_1;
    wire n3_adj_2408;
    wire \c0.FRAME_MATCHER_i_31_N_1312_5_cascade_ ;
    wire \c0.n3_adj_2256 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_4_cascade_ ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_3_cascade_ ;
    wire \c0.n3_adj_2258 ;
    wire \c0.n16379 ;
    wire \c0.n3_adj_2242 ;
    wire \c0.n3_adj_2243 ;
    wire \c0.n3_adj_2244 ;
    wire \c0.n17172_cascade_ ;
    wire data_in_0_7;
    wire data_in_1_5;
    wire data_in_0_4;
    wire n9472_cascade_;
    wire \c0.rx.n10086_cascade_ ;
    wire \c0.rx.r_SM_Main_2_N_2090_2 ;
    wire n14060_cascade_;
    wire n7866_cascade_;
    wire n10425_cascade_;
    wire n12;
    wire n13276;
    wire n10_adj_2415_cascade_;
    wire n15701;
    wire n16844;
    wire n17461;
    wire r_Clock_Count_1;
    wire n17601;
    wire n17602;
    wire r_Clock_Count_4_adj_2433;
    wire \c0.rx.n6 ;
    wire n16853;
    wire r_Clock_Count_1_adj_2436;
    wire n4_adj_2411;
    wire n17260;
    wire n10425;
    wire n16857;
    wire r_Clock_Count_5_adj_2432;
    wire n16858;
    wire r_Clock_Count_3_adj_2434;
    wire n9406;
    wire \c0.n3_adj_2217 ;
    wire \c0.n3_adj_2215 ;
    wire \c0.n3_adj_2210 ;
    wire \c0.n3_adj_2249 ;
    wire \c0.n9393 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_2_cascade_ ;
    wire \c0.n3_adj_2259 ;
    wire \c0.n10_adj_2329 ;
    wire \c0.n16895 ;
    wire \c0.n16895_cascade_ ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_1_cascade_ ;
    wire \c0.n3_adj_2260 ;
    wire bfn_4_22_0_;
    wire \c0.FRAME_MATCHER_i_31_N_1312_1 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_1 ;
    wire \c0.n15622 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_2 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_2 ;
    wire \c0.n15623 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_3 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_3 ;
    wire \c0.n15624 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_4 ;
    wire \c0.n15625 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_5 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_5 ;
    wire \c0.n15626 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_6 ;
    wire \c0.n15627 ;
    wire \c0.n15628 ;
    wire \c0.n15629 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_8 ;
    wire bfn_4_23_0_;
    wire \c0.FRAME_MATCHER_i_31_N_1280_9 ;
    wire \c0.n15630 ;
    wire \c0.n15631 ;
    wire \c0.n15632 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_12 ;
    wire \c0.n15633 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_13 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_13 ;
    wire \c0.n15634 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_14 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_14 ;
    wire \c0.n15635 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_15 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_15 ;
    wire \c0.n15636 ;
    wire \c0.n15637 ;
    wire bfn_4_24_0_;
    wire \c0.n15638 ;
    wire \c0.n15639 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_19 ;
    wire \c0.n15640 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_20 ;
    wire \c0.n15641 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_21 ;
    wire \c0.n15642 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_22 ;
    wire \c0.n15643 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_23 ;
    wire \c0.n15644 ;
    wire \c0.n15645 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_24 ;
    wire bfn_4_25_0_;
    wire \c0.FRAME_MATCHER_i_31_N_1280_25 ;
    wire \c0.n15646 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_26 ;
    wire \c0.n15647 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_27 ;
    wire \c0.n15648 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_28 ;
    wire \c0.n15649 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_29 ;
    wire \c0.n15650 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_30 ;
    wire \c0.n15651 ;
    wire \c0.n15652 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_31 ;
    wire data_in_0_6;
    wire \c0.n17274_cascade_ ;
    wire \c0.n17889 ;
    wire data_in_3_1;
    wire data_in_2_1;
    wire data_in_2_4;
    wire data_in_1_4;
    wire n17567;
    wire r_Clock_Count_4_adj_2450;
    wire data_in_2_3;
    wire n16856;
    wire r_Clock_Count_6_adj_2431;
    wire n16893_cascade_;
    wire n5;
    wire n17636;
    wire r_SM_Main_2_N_2033_1;
    wire r_Bit_Index_2;
    wire r_Bit_Index_1_adj_2438;
    wire r_Clock_Count_7;
    wire r_Clock_Count_6;
    wire r_Clock_Count_8;
    wire n9937;
    wire \c0.tx.n15683_cascade_ ;
    wire \c0.tx.n14082 ;
    wire n17573;
    wire r_Clock_Count_4;
    wire \c0.n12993_cascade_ ;
    wire \c0.n12993 ;
    wire \c0.n13298 ;
    wire \c0.n20_adj_2267 ;
    wire \c0.n21_adj_2271_cascade_ ;
    wire n29_cascade_;
    wire tx_enable;
    wire \c0.n12991 ;
    wire \c0.n12991_cascade_ ;
    wire \c0.n19_adj_2270 ;
    wire n16859;
    wire n17_adj_2416;
    wire r_Clock_Count_0_adj_2437;
    wire tx_o;
    wire data_in_1_0;
    wire n3977_cascade_;
    wire \c0.n3_adj_2233 ;
    wire \c0.n3_adj_2219 ;
    wire \c0.n16441 ;
    wire \c0.n3_adj_2229 ;
    wire \c0.n3_adj_2231 ;
    wire \c0.n3_adj_2227 ;
    wire \c0.n3_adj_2223 ;
    wire \c0.n3_adj_2225 ;
    wire \c0.n1439_cascade_ ;
    wire \c0.n3_adj_2221 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_7 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_7 ;
    wire \c0.n3_adj_2250 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_6 ;
    wire \c0.n3_adj_2253 ;
    wire \c0.n3_adj_2237 ;
    wire \c0.n3_adj_2235 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_11 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_11 ;
    wire \c0.n3_adj_2246 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_10 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_9 ;
    wire \c0.n3_adj_2248 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_8 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_19 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_20 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_21 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_23 ;
    wire \c0.n18_adj_2198_cascade_ ;
    wire \c0.n127_adj_2136_cascade_ ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_27 ;
    wire n9472;
    wire \c0.FRAME_MATCHER_i_31_N_1312_30 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_25 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_28 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_24 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_26 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_22 ;
    wire \c0.n12_adj_2200 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_31 ;
    wire n4_adj_2460;
    wire n4_adj_2417;
    wire data_in_0_2;
    wire data_in_1_3;
    wire n13082;
    wire \c0.n16891_cascade_ ;
    wire r_Bit_Index_0;
    wire \c0.rx.n9323 ;
    wire n9477;
    wire n4_adj_2409;
    wire n9477_cascade_;
    wire n16893;
    wire \c0.tx.n17462 ;
    wire \c0.tx.r_Bit_Index_0 ;
    wire n17397;
    wire \c0.tx.r_Bit_Index_2 ;
    wire \c0.tx.n17975_cascade_ ;
    wire \c0.tx.o_Tx_Serial_N_2064_cascade_ ;
    wire n3_adj_2406;
    wire \c0.n1419_cascade_ ;
    wire \c0.n1419 ;
    wire n53;
    wire \c0.delay_counter_0 ;
    wire \c0.n17637 ;
    wire bfn_5_31_0_;
    wire \c0.delay_counter_1 ;
    wire \c0.n6531 ;
    wire \c0.n15514 ;
    wire \c0.n6530 ;
    wire \c0.n15515 ;
    wire \c0.delay_counter_3 ;
    wire \c0.n6529 ;
    wire \c0.n15516 ;
    wire \c0.n6528 ;
    wire \c0.n15517 ;
    wire \c0.delay_counter_5 ;
    wire \c0.n17574 ;
    wire \c0.n15518 ;
    wire \c0.delay_counter_6 ;
    wire \c0.n6526 ;
    wire \c0.n15519 ;
    wire \c0.delay_counter_7 ;
    wire \c0.n17638 ;
    wire \c0.n15520 ;
    wire \c0.n15521 ;
    wire \c0.n6524 ;
    wire bfn_5_32_0_;
    wire \c0.delay_counter_9 ;
    wire \c0.n6523 ;
    wire \c0.n15522 ;
    wire \c0.delay_counter_10 ;
    wire \c0.n6522 ;
    wire \c0.n15523 ;
    wire \c0.delay_counter_11 ;
    wire \c0.n6521 ;
    wire \c0.n15524 ;
    wire \c0.delay_counter_12 ;
    wire \c0.n17575 ;
    wire \c0.n15525 ;
    wire \c0.n17639 ;
    wire \c0.n15526 ;
    wire \c0.delay_counter_14 ;
    wire \c0.n15527 ;
    wire \c0.n17635 ;
    wire \c0.n16331 ;
    wire \c0.n16381 ;
    wire \c0.FRAME_MATCHER_i_19 ;
    wire \c0.FRAME_MATCHER_i_24 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_16 ;
    wire n1716_cascade_;
    wire n14;
    wire n16775;
    wire n3977;
    wire n16775_cascade_;
    wire n9453;
    wire \c0.FRAME_MATCHER_i_1 ;
    wire n2275;
    wire n2275_cascade_;
    wire \c0.n7212_cascade_ ;
    wire \c0.n17452_cascade_ ;
    wire \c0.n17454 ;
    wire \c0.n7_cascade_ ;
    wire \c0.n16335 ;
    wire \c0.FRAME_MATCHER_state_5 ;
    wire \c0.FRAME_MATCHER_state_6 ;
    wire \c0.FRAME_MATCHER_state_29 ;
    wire \c0.n59_cascade_ ;
    wire \c0.n5_adj_2262_cascade_ ;
    wire \c0.n16876_cascade_ ;
    wire \c0.n60_cascade_ ;
    wire \c0.n16363 ;
    wire \c0.FRAME_MATCHER_state_30 ;
    wire \c0.FRAME_MATCHER_state_23 ;
    wire \c0.n9451_cascade_ ;
    wire n12933_cascade_;
    wire \c0.n9451 ;
    wire \c0.n9 ;
    wire \c0.n17258 ;
    wire \c0.n28_cascade_ ;
    wire \c0.n60 ;
    wire \c0.n16879 ;
    wire \c0.n33 ;
    wire \c0.n16879_cascade_ ;
    wire \c0.FRAME_MATCHER_i_6 ;
    wire \c0.FRAME_MATCHER_i_7 ;
    wire \c0.FRAME_MATCHER_i_9 ;
    wire n9445;
    wire \c0.n9488 ;
    wire \c0.n12_adj_2158 ;
    wire \c0.n9488_cascade_ ;
    wire \c0.n17262 ;
    wire \c0.n17256 ;
    wire data_in_0_0;
    wire \c0.n9485 ;
    wire \c0.n10_adj_2149_cascade_ ;
    wire \c0.FRAME_MATCHER_i_29 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_29 ;
    wire data_in_3_0;
    wire data_in_0_5;
    wire data_in_3_4;
    wire \c0.n17264 ;
    wire \c0.n9493 ;
    wire \c0.n12_cascade_ ;
    wire \c0.FRAME_MATCHER_i_31 ;
    wire n127_adj_2418_cascade_;
    wire \c0.n17240 ;
    wire data_in_1_1;
    wire \c0.n9482 ;
    wire \c0.n9490 ;
    wire n16795;
    wire n127_cascade_;
    wire \c0.n2 ;
    wire \c0.n2_cascade_ ;
    wire n9435;
    wire n7198;
    wire \c0.FRAME_MATCHER_i_31_N_1312_18 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_18 ;
    wire \c0.FRAME_MATCHER_i_18 ;
    wire \c0.n3_adj_2239 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_17 ;
    wire \c0.n127_adj_2136 ;
    wire n127;
    wire \c0.FRAME_MATCHER_i_31_N_1312_16 ;
    wire n127_adj_2418;
    wire \c0.FRAME_MATCHER_i_16 ;
    wire \c0.n7212 ;
    wire \c0.n3_adj_2241 ;
    wire \c0.data_in_frame_9_2 ;
    wire \c0.n15939 ;
    wire \c0.data_in_frame_10_0 ;
    wire \c0.n17013_cascade_ ;
    wire \c0.n17013 ;
    wire \c0.data_in_frame_9_7 ;
    wire data_in_3_6;
    wire data_in_2_0;
    wire \c0.n17268 ;
    wire data_in_1_7;
    wire data_in_0_3;
    wire \c0.n19_adj_2199 ;
    wire \c0.data_in_frame_10_1 ;
    wire \c0.n9743 ;
    wire \c0.n16954_cascade_ ;
    wire \c0.data_in_frame_10_6 ;
    wire \c0.n18_adj_2174_cascade_ ;
    wire \c0.n17015 ;
    wire \c0.data_in_frame_9_4 ;
    wire \c0.n6_adj_2152 ;
    wire \c0.n13272 ;
    wire \c0.n16882_cascade_ ;
    wire \c0.data_in_frame_10_4 ;
    wire \c0.data_in_frame_9_6 ;
    wire \c0.data_in_frame_2_7 ;
    wire \c0.n25_adj_2324 ;
    wire n4_adj_2458_cascade_;
    wire r_SM_Main_0;
    wire n14060;
    wire r_SM_Main_1;
    wire r_SM_Main_2;
    wire n17395;
    wire \c0.tx_active_prev ;
    wire \c0.n65 ;
    wire bfn_6_30_0_;
    wire \c0.n15653 ;
    wire \c0.n15654 ;
    wire \c0.n15655 ;
    wire \c0.n15656 ;
    wire \c0.n15657 ;
    wire \c0.n15658 ;
    wire \c0.n15659 ;
    wire \c0.n8938_cascade_ ;
    wire \c0.n22_adj_2164 ;
    wire \c0.n22_adj_2164_cascade_ ;
    wire \c0.tx_transmit_N_1949_1 ;
    wire \c0.n15868_cascade_ ;
    wire \c0.n8631 ;
    wire n10141_cascade_;
    wire \c0.n446 ;
    wire \c0.n446_cascade_ ;
    wire \c0.n456 ;
    wire \c0.n16371 ;
    wire \c0.n16453 ;
    wire \c0.n59 ;
    wire \c0.n61_cascade_ ;
    wire \c0.n10_adj_2336 ;
    wire \c0.n16133_cascade_ ;
    wire \c0.n16898 ;
    wire \c0.FRAME_MATCHER_state_19 ;
    wire \c0.n52 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_4 ;
    wire \c0.n3_adj_2257 ;
    wire \c0.FRAME_MATCHER_i_20 ;
    wire \c0.FRAME_MATCHER_i_4 ;
    wire \c0.FRAME_MATCHER_i_5 ;
    wire \c0.FRAME_MATCHER_i_21 ;
    wire \c0.n30_cascade_ ;
    wire \c0.FRAME_MATCHER_i_13 ;
    wire \c0.n56 ;
    wire \c0.FRAME_MATCHER_state_10 ;
    wire \c0.n6_adj_2213 ;
    wire \c0.n16869 ;
    wire \c0.n16869_cascade_ ;
    wire \c0.n16871_cascade_ ;
    wire \c0.n16876 ;
    wire \c0.n50 ;
    wire \c0.n46 ;
    wire \c0.n56_adj_2146_cascade_ ;
    wire \c0.n51 ;
    wire \c0.n9346 ;
    wire \c0.FRAME_MATCHER_i_3 ;
    wire \c0.FRAME_MATCHER_i_2 ;
    wire \c0.FRAME_MATCHER_i_28 ;
    wire \c0.n45 ;
    wire \c0.FRAME_MATCHER_i_27 ;
    wire \c0.FRAME_MATCHER_i_30 ;
    wire \c0.FRAME_MATCHER_i_8 ;
    wire \c0.FRAME_MATCHER_i_26 ;
    wire \c0.n47_adj_2144 ;
    wire \c0.FRAME_MATCHER_i_22 ;
    wire \c0.FRAME_MATCHER_i_23 ;
    wire \c0.FRAME_MATCHER_i_25 ;
    wire \c0.n49 ;
    wire \c0.FRAME_MATCHER_state_22 ;
    wire \c0.n16365 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_12 ;
    wire \c0.FRAME_MATCHER_i_12 ;
    wire \c0.n3_adj_2245 ;
    wire \c0.n16351 ;
    wire \c0.FRAME_MATCHER_state_21 ;
    wire \c0.n16367 ;
    wire \c0.FRAME_MATCHER_state_26 ;
    wire \c0.n16357 ;
    wire \c0.FRAME_MATCHER_state_27 ;
    wire \c0.n16355 ;
    wire data_in_0_1;
    wire \c0.n17266 ;
    wire data_in_3_5;
    wire data_in_2_5;
    wire data_in_2_7;
    wire \c0.n8_adj_2157 ;
    wire data_in_3_7;
    wire data_in_3_3;
    wire data_in_frame_7_0;
    wire data_in_frame_7_6;
    wire n16896;
    wire rx_data_6;
    wire rx_data_0;
    wire \c0.n2351_cascade_ ;
    wire data_in_frame_6_7;
    wire data_in_frame_6_1;
    wire \c0.n2352_cascade_ ;
    wire data_in_frame_6_3;
    wire data_in_frame_6_4;
    wire \c0.n23_adj_2145 ;
    wire \c0.n9541_cascade_ ;
    wire \c0.n16943 ;
    wire data_in_frame_0_2;
    wire \c0.data_in_frame_2_5 ;
    wire \c0.data_in_frame_2_3 ;
    wire \c0.n2336_cascade_ ;
    wire \c0.data_in_frame_1_5 ;
    wire \c0.n20_adj_2340_cascade_ ;
    wire data_in_3_2;
    wire data_in_2_2;
    wire data_in_1_2;
    wire \c0.data_in_frame_10_3 ;
    wire data_in_frame_6_6;
    wire data_in_frame_7_7;
    wire data_in_frame_7_2;
    wire data_in_frame_6_2;
    wire \c0.n22_cascade_ ;
    wire \c0.n27 ;
    wire rx_data_7;
    wire \c0.data_in_frame_1_0 ;
    wire n17634;
    wire r_Clock_Count_6_adj_2448;
    wire \c0.n9585 ;
    wire \c0.data_in_frame_2_2 ;
    wire \c0.n22_adj_2301 ;
    wire \c0.n9585_cascade_ ;
    wire data_in_frame_7_1;
    wire data_in_frame_7_4;
    wire rx_data_2;
    wire data_in_frame_0_0;
    wire \c0.data_in_frame_1_6 ;
    wire \c0.data_in_frame_10_2 ;
    wire data_in_frame_0_1;
    wire \c0.n17460 ;
    wire r_Tx_Data_3;
    wire \c0.delay_counter_13 ;
    wire \c0.delay_counter_8 ;
    wire \c0.delay_counter_4 ;
    wire \c0.delay_counter_2 ;
    wire \c0.n17236 ;
    wire \c0.n42_adj_2165 ;
    wire \c0.byte_transmit_counter_5 ;
    wire \c0.n17254 ;
    wire \c0.n17254_cascade_ ;
    wire \c0.n17290 ;
    wire \c0.tx_transmit_N_1949_5 ;
    wire \c0.n5_adj_2319 ;
    wire \c0.tx_transmit_N_1949_6 ;
    wire \c0.byte_transmit_counter_6 ;
    wire \c0.n23_adj_2309 ;
    wire \c0.n17278 ;
    wire \c0.n17276 ;
    wire \c0.tx_transmit_N_1949_0 ;
    wire \c0.n16839_cascade_ ;
    wire \c0.tx_transmit_N_1949_4 ;
    wire \c0.n8938 ;
    wire \c0.tx_transmit_N_1949_3 ;
    wire \c0.n16839 ;
    wire \c0.tx_transmit_N_1949_7 ;
    wire \c0.byte_transmit_counter_7 ;
    wire n17834_cascade_;
    wire n17162;
    wire n9358_cascade_;
    wire n41_cascade_;
    wire n35;
    wire n29;
    wire n445;
    wire n10031;
    wire n17479_cascade_;
    wire n16886;
    wire n38;
    wire \c0.n44_adj_2163 ;
    wire n9357;
    wire \c0.tx_transmit_N_1949_2 ;
    wire \c0.n4_adj_2311 ;
    wire \c0.n17475 ;
    wire \c0.tx2_transmit_N_1997_cascade_ ;
    wire \c0.tx2.n113 ;
    wire \c0.tx2.n113_cascade_ ;
    wire \c0.r_SM_Main_2_N_2036_0_adj_2261 ;
    wire n491;
    wire n491_cascade_;
    wire n17;
    wire \c0.n16369 ;
    wire \c0.n12_adj_2189 ;
    wire \c0.FRAME_MATCHER_state_20 ;
    wire n9460;
    wire n9460_cascade_;
    wire n9462;
    wire \c0.FRAME_MATCHER_state_18 ;
    wire \c0.n16343 ;
    wire data_in_2_6;
    wire rx_data_ready;
    wire data_in_1_6;
    wire \c0.n8603 ;
    wire \c0.FRAME_MATCHER_i_11 ;
    wire \c0.FRAME_MATCHER_i_14 ;
    wire \c0.FRAME_MATCHER_i_15 ;
    wire \c0.n48 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_10 ;
    wire \c0.FRAME_MATCHER_i_10 ;
    wire \c0.n3_adj_2247 ;
    wire \c0.n9819_cascade_ ;
    wire \c0.FRAME_MATCHER_state_25 ;
    wire \c0.n16359 ;
    wire \c0.FRAME_MATCHER_i_31_N_1280_17 ;
    wire \c0.FRAME_MATCHER_i_17 ;
    wire \c0.n3_adj_2240 ;
    wire data_in_frame_0_7;
    wire \c0.data_in_frame_1_7 ;
    wire \c0.data_in_frame_1_4 ;
    wire \c0.n27_adj_2342 ;
    wire \c0.n23_adj_2341_cascade_ ;
    wire \c0.data_in_frame_1_3 ;
    wire \c0.n21_adj_2171 ;
    wire \c0.n15930 ;
    wire \c0.data_in_frame_10_7 ;
    wire \c0.n17352_cascade_ ;
    wire \c0.n27_adj_2196 ;
    wire \c0.n25 ;
    wire \c0.n15846_cascade_ ;
    wire \c0.n15929 ;
    wire \c0.n26_adj_2184 ;
    wire \c0.n15938 ;
    wire \c0.data_in_frame_1_2 ;
    wire \c0.data_in_frame_9_3 ;
    wire \c0.data_in_frame_1_1 ;
    wire \c0.n17014 ;
    wire \c0.n23_adj_2156_cascade_ ;
    wire \c0.n17001 ;
    wire \c0.n28_adj_2183 ;
    wire data_in_frame_0_6;
    wire \c0.n2340 ;
    wire \c0.data_in_frame_9_0 ;
    wire \c0.n17004 ;
    wire \c0.n19 ;
    wire data_in_frame_7_3;
    wire \c0.n2336 ;
    wire data_in_frame_7_5;
    wire \c0.n9541 ;
    wire data_in_frame_6_0;
    wire data_in_frame_6_5;
    wire \c0.n20_cascade_ ;
    wire \c0.n2342 ;
    wire \c0.data_in_frame_9_1 ;
    wire \c0.n8_adj_2310 ;
    wire \c0.data_in_frame_9_5 ;
    wire tx2_o;
    wire \c0.tx2.n18113_cascade_ ;
    wire n10398;
    wire n17194;
    wire n10398_cascade_;
    wire \c0.tx2.n17906 ;
    wire \c0.tx2.n18116 ;
    wire \c0.tx2.o_Tx_Serial_N_2064_cascade_ ;
    wire r_SM_Main_0_adj_2445;
    wire n3;
    wire n5029;
    wire r_Bit_Index_2_adj_2455;
    wire \c0.tx2.n13281 ;
    wire \c0.n2_adj_2266_cascade_ ;
    wire \c0.n18098_cascade_ ;
    wire \c0.n10_adj_2139_cascade_ ;
    wire \c0.rx.r_Rx_Data_R ;
    wire r_Tx_Data_0;
    wire n17394;
    wire \c0.n8_adj_2160 ;
    wire \c0.n15_cascade_ ;
    wire \c0.n12_adj_2150_cascade_ ;
    wire r_Tx_Data_2;
    wire n10_adj_2426;
    wire n10_adj_2407_cascade_;
    wire r_Tx_Data_4;
    wire \c0.n17590_cascade_ ;
    wire n18026;
    wire \c0.n16347 ;
    wire \c0.n16761 ;
    wire \c0.FRAME_MATCHER_state_28 ;
    wire \c0.n16353 ;
    wire \c0.FRAME_MATCHER_state_24 ;
    wire \c0.n16361 ;
    wire \c0.FRAME_MATCHER_state_17 ;
    wire \c0.n16345 ;
    wire \c0.FRAME_MATCHER_state_4 ;
    wire \c0.n4 ;
    wire \c0.n16339 ;
    wire \c0.FRAME_MATCHER_state_14 ;
    wire \c0.n16871 ;
    wire \c0.n16772 ;
    wire \c0.n17349_cascade_ ;
    wire \c0.n1439 ;
    wire \c0.FRAME_MATCHER_i_31_N_1312_0 ;
    wire \c0.n5_adj_2322 ;
    wire \c0.n5_cascade_ ;
    wire \c0.n17328_cascade_ ;
    wire \c0.FRAME_MATCHER_state_8 ;
    wire \c0.n16905 ;
    wire \c0.n17337_cascade_ ;
    wire data_in_frame_0_4;
    wire data_in_frame_0_5;
    wire \c0.n2338 ;
    wire \c0.data_in_frame_2_6 ;
    wire \c0.data_in_frame_2_0 ;
    wire \c0.n2338_cascade_ ;
    wire \c0.n2352 ;
    wire \c0.n26_adj_2344 ;
    wire \c0.n17_adj_2346_cascade_ ;
    wire \c0.n30_adj_2345 ;
    wire n31_cascade_;
    wire \c0.tx2.tx2_active ;
    wire \c0.n17334_cascade_ ;
    wire \c0.n2334 ;
    wire \c0.n2351 ;
    wire \c0.n18_adj_2343 ;
    wire rx_data_3;
    wire n16897;
    wire data_in_frame_0_3;
    wire \c0.n17918_cascade_ ;
    wire \c0.n17343 ;
    wire \c0.n17769 ;
    wire \c0.n18 ;
    wire \c0.n17 ;
    wire \c0.n26_adj_2147 ;
    wire \c0.n30_adj_2148 ;
    wire rx_data_5;
    wire \c0.n16882 ;
    wire \c0.data_in_frame_10_5 ;
    wire r_SM_Main_1_adj_2444;
    wire \c0.tx2.n6480 ;
    wire \c0.tx2.n1 ;
    wire \c0.tx2.n10101 ;
    wire data_out_frame2_18_5;
    wire r_SM_Main_2_adj_2439;
    wire n13440;
    wire r_SM_Main_1_adj_2440;
    wire rx_data_1;
    wire \c0.data_in_frame_2_1 ;
    wire \c0.n16891 ;
    wire \c0.n8 ;
    wire rx_data_4;
    wire \c0.data_in_frame_2_4 ;
    wire \c0.r_SM_Main_2_N_2036_0 ;
    wire tx_active;
    wire n17230;
    wire data_out_1_7;
    wire \c0.n10 ;
    wire r_SM_Main_2_adj_2443;
    wire n17544;
    wire r_Clock_Count_0_adj_2454;
    wire r_Bit_Index_1;
    wire n17398;
    wire \c0.n29_cascade_ ;
    wire r_Tx_Data_1;
    wire r_Tx_Data_5;
    wire \c0.data_out_0_6 ;
    wire \c0.n9_adj_2143_cascade_ ;
    wire \c0.n23 ;
    wire \c0.n17547 ;
    wire \c0.n5_adj_2326_cascade_ ;
    wire \c0.n18023 ;
    wire r_Tx_Data_7;
    wire \c0.n18014 ;
    wire \c0.n17585 ;
    wire n10_adj_2423;
    wire n18044_cascade_;
    wire n10_adj_2414;
    wire data_out_0_1;
    wire \c0.n18080 ;
    wire data_out_3_7;
    wire \c0.n2_adj_2137 ;
    wire \c0.data_out_1_4 ;
    wire n16776;
    wire n17208;
    wire n8828;
    wire \c0.FRAME_MATCHER_state_16 ;
    wire \c0.n47 ;
    wire \c0.n6_adj_2140 ;
    wire FRAME_MATCHER_state_1;
    wire \c0.n5_adj_2339 ;
    wire \c0.n16814_cascade_ ;
    wire \c0.tx2.n89 ;
    wire \c0.FRAME_MATCHER_state_31 ;
    wire \c0.n16377 ;
    wire n9452;
    wire n12933;
    wire \c0.FRAME_MATCHER_i_31_N_1280_0 ;
    wire \c0.FRAME_MATCHER_i_0 ;
    wire \c0.n3 ;
    wire \c0.FRAME_MATCHER_state_12 ;
    wire \c0.n4_adj_2360 ;
    wire \c0.n16449 ;
    wire data_out_frame2_18_2;
    wire \c0.n18119_cascade_ ;
    wire \c0.n18122_cascade_ ;
    wire \c0.tx2.r_Tx_Data_2 ;
    wire \c0.n17340 ;
    wire \c0.n13496 ;
    wire data_out_frame2_7_3;
    wire FRAME_MATCHER_state_2;
    wire \c0.FRAME_MATCHER_state_3 ;
    wire \c0.n62 ;
    wire \c0.n13464 ;
    wire \c0.n2_adj_2330_cascade_ ;
    wire \c0.n9758 ;
    wire \c0.n17915 ;
    wire data_out_frame2_18_1;
    wire \c0.n17909_cascade_ ;
    wire \c0.n6 ;
    wire \c0.n18107 ;
    wire \c0.n17579 ;
    wire \c0.n17912 ;
    wire \c0.n18110 ;
    wire \c0.n22_adj_2359_cascade_ ;
    wire \c0.tx2.r_Tx_Data_1 ;
    wire \c0.n17548 ;
    wire \c0.n17589 ;
    wire \c0.n2_adj_2298 ;
    wire \c0.n18029_cascade_ ;
    wire \c0.n8_adj_2138 ;
    wire \c0.n5_adj_2299 ;
    wire r_SM_Main_0_adj_2441;
    wire \c0.rx.r_SM_Main_2_N_2096_0 ;
    wire r_Rx_Data;
    wire n1;
    wire data_out_3_5;
    wire data_out_2_5;
    wire \c0.n9530 ;
    wire data_out_1_6;
    wire data_out_2_0;
    wire \c0.n9509 ;
    wire \c0.data_out_7_5 ;
    wire \c0.n26 ;
    wire n18032;
    wire n10;
    wire \c0.n5_adj_2142 ;
    wire data_out_3_0;
    wire \c0.data_out_3_6 ;
    wire \c0.n10054_cascade_ ;
    wire \c0.data_out_7_7 ;
    wire \c0.n5_adj_2188_cascade_ ;
    wire \c0.n18041 ;
    wire \c0.n5_adj_2208 ;
    wire \c0.n17543_cascade_ ;
    wire \c0.n18011 ;
    wire \c0.n17445 ;
    wire \c0.n17456_cascade_ ;
    wire \c0.n10054 ;
    wire n9361;
    wire n17154;
    wire FRAME_MATCHER_state_0;
    wire \c0.tx2_transmit_N_1997 ;
    wire bfn_12_18_0_;
    wire \c0.n15615 ;
    wire \c0.n15616 ;
    wire \c0.n15617 ;
    wire \c0.n15618 ;
    wire \c0.byte_transmit_counter2_5 ;
    wire \c0.n15619 ;
    wire \c0.byte_transmit_counter2_6 ;
    wire \c0.n15620 ;
    wire \c0.n15621 ;
    wire \c0.byte_transmit_counter2_7 ;
    wire \c0.n10052 ;
    wire \c0.n10297 ;
    wire \c0.n7 ;
    wire \c0.FRAME_MATCHER_state_9 ;
    wire \c0.n16455 ;
    wire \c0.n17927 ;
    wire data_out_frame2_17_2;
    wire \c0.n17930_cascade_ ;
    wire \c0.n22_adj_2358 ;
    wire \c0.n17936 ;
    wire \c0.n6_adj_2201 ;
    wire \c0.n17942 ;
    wire \c0.n17560 ;
    wire \c0.n17301_cascade_ ;
    wire \c0.n17303_cascade_ ;
    wire \c0.tx2.r_Tx_Data_0 ;
    wire data_out_frame2_18_0;
    wire data_out_frame2_17_0;
    wire \c0.n18101_cascade_ ;
    wire \c0.n18104_cascade_ ;
    wire \c0.n22_adj_2337 ;
    wire \c0.n17939 ;
    wire data_out_frame2_6_3;
    wire \c0.n16_adj_2197 ;
    wire \c0.n22_adj_2194 ;
    wire \c0.n9754 ;
    wire \c0.n9901_cascade_ ;
    wire data_out_frame2_5_3;
    wire \c0.n16148 ;
    wire \c0.n17331_cascade_ ;
    wire \c0.n15846 ;
    wire \c0.n17891 ;
    wire data_out_frame2_10_2;
    wire \c0.n12_adj_2305 ;
    wire \c0.n17990 ;
    wire \c0.n17993_cascade_ ;
    wire \c0.n17894 ;
    wire \c0.n17393_cascade_ ;
    wire \c0.n17571 ;
    wire \c0.n17963_cascade_ ;
    wire \c0.n17966_cascade_ ;
    wire \c0.tx2.r_Tx_Data_5 ;
    wire data_out_0_5;
    wire data_out_0_3;
    wire data_out_2_2;
    wire \c0.n2_adj_2291 ;
    wire data_out_3_2;
    wire data_out_frame2_9_4;
    wire \c0.n9_adj_2347 ;
    wire \c0.n17897 ;
    wire \c0.n8_adj_2348_cascade_ ;
    wire \c0.n17900 ;
    wire r_Bit_Index_1_adj_2456;
    wire r_Bit_Index_0_adj_2457;
    wire \c0.tx2.n17903 ;
    wire \c0.n16975 ;
    wire \c0.n16978_cascade_ ;
    wire \c0.n16912 ;
    wire \c0.n21 ;
    wire \c0.n17588 ;
    wire \c0.n1 ;
    wire n18038_cascade_;
    wire n8730;
    wire n10_adj_2413_cascade_;
    wire byte_transmit_counter_4;
    wire r_Tx_Data_6;
    wire \c0.data_out_1_1 ;
    wire \c0.n10181 ;
    wire \c0.data_out_6_6 ;
    wire \c0.n5_adj_2300 ;
    wire \c0.n17555_cascade_ ;
    wire \c0.n18035 ;
    wire \c0.n17569 ;
    wire \c0.data_out_frame2_0_2 ;
    wire \c0.n17578 ;
    wire \c0.data_out_frame2_0_4 ;
    wire \c0.n6_adj_2335 ;
    wire \c0.n5_adj_2317 ;
    wire \c0.n16957 ;
    wire \c0.n17106 ;
    wire \c0.n16957_cascade_ ;
    wire \c0.n15_adj_2269 ;
    wire \c0.data_out_frame2_20_1 ;
    wire \c0.n17061 ;
    wire \c0.data_out_frame2_20_0 ;
    wire \c0.n9810 ;
    wire \c0.n17_adj_2193 ;
    wire \c0.n16_cascade_ ;
    wire \c0.n17112_cascade_ ;
    wire \c0.n14_adj_2308_cascade_ ;
    wire \c0.data_out_frame2_19_5 ;
    wire \c0.n17933 ;
    wire data_out_frame2_15_3;
    wire data_out_frame2_13_4;
    wire \c0.n11 ;
    wire \c0.n17981 ;
    wire \c0.n17984_cascade_ ;
    wire \c0.n22_adj_2354 ;
    wire data_out_frame2_17_5;
    wire bfn_13_25_0_;
    wire n15528;
    wire n15529;
    wire n15530;
    wire n15531;
    wire n15532;
    wire n15533;
    wire n15534;
    wire n15535;
    wire bfn_13_26_0_;
    wire n15536;
    wire n15537;
    wire n15538;
    wire n15539;
    wire n15540;
    wire n15541;
    wire n15542;
    wire n15543;
    wire bfn_13_27_0_;
    wire n15544;
    wire n15545;
    wire n15546;
    wire n15547;
    wire n15548;
    wire n15549;
    wire n15550;
    wire n15551;
    wire bfn_13_28_0_;
    wire n15552;
    wire n15553;
    wire n15554;
    wire n15555;
    wire n15556;
    wire n15557;
    wire n15558;
    wire rand_setpoint_0;
    wire bfn_13_29_0_;
    wire rand_data_1;
    wire n15559;
    wire rand_data_2;
    wire n15560;
    wire rand_setpoint_3;
    wire n15561;
    wire rand_setpoint_4;
    wire n15562;
    wire n15563;
    wire n15564;
    wire n15565;
    wire n15566;
    wire rand_setpoint_8;
    wire bfn_13_30_0_;
    wire rand_setpoint_9;
    wire n15567;
    wire rand_data_10;
    wire n15568;
    wire rand_setpoint_11;
    wire n15569;
    wire rand_setpoint_12;
    wire n15570;
    wire rand_setpoint_13;
    wire n15571;
    wire rand_setpoint_14;
    wire n15572;
    wire rand_setpoint_15;
    wire n15573;
    wire n15574;
    wire bfn_13_31_0_;
    wire n15575;
    wire n15576;
    wire rand_data_19;
    wire n15577;
    wire n15578;
    wire n15579;
    wire rand_setpoint_22;
    wire n15580;
    wire n15581;
    wire n15582;
    wire bfn_13_32_0_;
    wire rand_setpoint_25;
    wire n15583;
    wire n15584;
    wire n15585;
    wire n15586;
    wire n15587;
    wire rand_setpoint_30;
    wire n15588;
    wire n15589;
    wire rand_setpoint_31;
    wire \c0.data_out_7_4 ;
    wire \c0.n22_adj_2357_cascade_ ;
    wire \c0.tx2.r_Tx_Data_3 ;
    wire \c0.n6_adj_2187 ;
    wire \c0.n18128 ;
    wire \c0.n16936 ;
    wire \c0.n18_adj_2331 ;
    wire \c0.n17100_cascade_ ;
    wire \c0.n16_adj_2332_cascade_ ;
    wire \c0.n20_adj_2333 ;
    wire \c0.data_out_frame2_19_0 ;
    wire \c0.n9886 ;
    wire \c0.n12_adj_2263_cascade_ ;
    wire \c0.data_out_frame2_20_2 ;
    wire \c0.n17112 ;
    wire \c0.n16_adj_2312_cascade_ ;
    wire \c0.n17097 ;
    wire data_out_frame2_6_0;
    wire \c0.n5_adj_2334 ;
    wire \c0.data_out_frame2_0_1 ;
    wire \c0.n17124 ;
    wire \c0.n14_adj_2264 ;
    wire data_out_frame2_16_2;
    wire \c0.n17031 ;
    wire \c0.n17091 ;
    wire \c0.n17031_cascade_ ;
    wire \c0.n9692 ;
    wire \c0.n17085 ;
    wire data_out_frame2_9_3;
    wire \c0.n17085_cascade_ ;
    wire \c0.n17073 ;
    wire data_out_frame2_18_4;
    wire \c0.data_out_frame2_19_4 ;
    wire \c0.n9707 ;
    wire \c0.n16963 ;
    wire \c0.n9579 ;
    wire \c0.n9579_cascade_ ;
    wire \c0.n10_adj_2307 ;
    wire \c0.n17957 ;
    wire \c0.n16908 ;
    wire \c0.n16908_cascade_ ;
    wire \c0.n6_adj_2286 ;
    wire data_out_frame2_14_4;
    wire \c0.n5543 ;
    wire \c0.n5545 ;
    wire n31;
    wire rand_data_4;
    wire n10197_cascade_;
    wire data_out_frame2_15_4;
    wire data_out_frame2_12_5;
    wire \c0.n17049 ;
    wire data_out_frame2_5_2;
    wire \c0.n9865 ;
    wire \c0.n6_adj_2306_cascade_ ;
    wire rand_data_27;
    wire rand_data_9;
    wire data_out_frame2_17_1;
    wire data_out_frame2_10_4;
    wire \c0.n10_adj_2191 ;
    wire \c0.n14 ;
    wire \c0.n17528 ;
    wire data_out_9_2;
    wire \c0.n17064 ;
    wire \c0.n12_adj_2289_cascade_ ;
    wire \c0.data_out_7_6 ;
    wire \c0.n9716_cascade_ ;
    wire \c0.n9728 ;
    wire \c0.n10_adj_2162_cascade_ ;
    wire data_out_9__2__N_367;
    wire data_out_9__2__N_367_cascade_;
    wire rand_setpoint_7;
    wire \c0.n8_adj_2169_cascade_ ;
    wire n10_adj_2427;
    wire \c0.n9496 ;
    wire \c0.n9716 ;
    wire rand_setpoint_2;
    wire \c0.n17594 ;
    wire \c0.n8_adj_2176 ;
    wire \c0.data_out_1_2 ;
    wire data_out_2_7;
    wire rand_setpoint_20;
    wire \c0.n17518 ;
    wire rand_setpoint_19;
    wire \c0.n17514 ;
    wire rand_setpoint_18;
    wire \c0.n17507 ;
    wire rand_setpoint_17;
    wire \c0.n17506_cascade_ ;
    wire rand_setpoint_26;
    wire rand_setpoint_29;
    wire rand_setpoint_24;
    wire rand_setpoint_27;
    wire rand_setpoint_28;
    wire data_out_frame2_7_1;
    wire data_out_frame2_10_5;
    wire \c0.n9763 ;
    wire data_out_frame2_8_2;
    wire \c0.n9916 ;
    wire data_out_frame2_12_4;
    wire \c0.n17037 ;
    wire \c0.n16933_cascade_ ;
    wire \c0.n17_adj_2313 ;
    wire \c0.n17960 ;
    wire \c0.n18125 ;
    wire \c0.n15_adj_2320_cascade_ ;
    wire \c0.n17088 ;
    wire \c0.data_out_frame2_19_2 ;
    wire \c0.n14_adj_2323 ;
    wire \c0.n17052 ;
    wire \c0.n17121 ;
    wire \c0.n19_adj_2254 ;
    wire \c0.n21_adj_2255_cascade_ ;
    wire \c0.data_out_frame2_20_3 ;
    wire data_out_frame2_14_5;
    wire \c0.n17022 ;
    wire \c0.n26_adj_2273 ;
    wire \c0.data_out_frame2_0_5 ;
    wire \c0.n17103 ;
    wire \c0.n17067 ;
    wire \c0.n17100 ;
    wire \c0.n9749 ;
    wire data_out_frame2_5_1;
    wire \c0.n9776 ;
    wire \c0.n9555 ;
    wire \c0.n16946 ;
    wire \c0.n22_adj_2207_cascade_ ;
    wire \c0.n18_adj_2251 ;
    wire \c0.n9892_cascade_ ;
    wire \c0.n17079 ;
    wire \c0.n20_adj_2202 ;
    wire \c0.n17079_cascade_ ;
    wire \c0.n24 ;
    wire \c0.data_out_frame2_20_5 ;
    wire data_out_frame2_10_7;
    wire rand_data_28;
    wire data_out_frame2_15_2;
    wire data_out_frame2_16_1;
    wire rand_data_20;
    wire \c0.n9814 ;
    wire \c0.n16987 ;
    wire \c0.n25_adj_2275 ;
    wire rand_data_17;
    wire data_out_frame2_6_4;
    wire \c0.n5_adj_2141_cascade_ ;
    wire \c0.n17987 ;
    wire \c0.n17951 ;
    wire data_out_frame2_13_3;
    wire \c0.n17954 ;
    wire \c0.n18056 ;
    wire data_out_frame2_7_0;
    wire \c0.n17346 ;
    wire rand_data_26;
    wire data_out_frame2_14_2;
    wire rand_data_0;
    wire data_out_frame2_9_0;
    wire \c0.n32_adj_2297 ;
    wire \c0.data_out_6_4 ;
    wire \c0.data_out_10_0 ;
    wire \c0.n16966 ;
    wire \c0.n16966_cascade_ ;
    wire \c0.n16918 ;
    wire \c0.n10_adj_2288_cascade_ ;
    wire \c0.n17109 ;
    wire \c0.n16990 ;
    wire \c0.data_out_6_1 ;
    wire rand_setpoint_5;
    wire data_out_8_5;
    wire \c0.n28_adj_2287 ;
    wire rand_setpoint_6;
    wire data_out_8_6;
    wire \c0.data_out_10_7 ;
    wire \c0.n8_adj_2166 ;
    wire n10_adj_2425;
    wire \c0.n17055 ;
    wire \c0.data_out_9_5 ;
    wire \c0.data_out_10_1 ;
    wire \c0.data_out_8_2 ;
    wire \c0.data_out_10_5 ;
    wire rand_setpoint_1;
    wire \c0.data_out_7_1 ;
    wire \c0.data_out_9_0 ;
    wire \c0.data_out_5_2 ;
    wire \c0.n9522 ;
    wire data_out_8_1;
    wire \c0.n18077 ;
    wire \c0.data_out_7__2__N_447 ;
    wire rand_setpoint_23;
    wire \c0.n17532_cascade_ ;
    wire \c0.data_out_6_7 ;
    wire \c0.data_out_5_5 ;
    wire \c0.n17025 ;
    wire \c0.n17534 ;
    wire \c0.data_out_frame2_0_3 ;
    wire \c0.n17576 ;
    wire data_out_frame2_8_3;
    wire \c0.n9839 ;
    wire data_out_frame2_18_6;
    wire \c0.n16994 ;
    wire rand_data_21;
    wire \c0.n28_adj_2294 ;
    wire \c0.n32_cascade_ ;
    wire \c0.n31 ;
    wire \c0.n29_adj_2296 ;
    wire \c0.n16933 ;
    wire \c0.n16915_cascade_ ;
    wire data_out_frame2_7_2;
    wire \c0.n19_adj_2303 ;
    wire \c0.n20_adj_2302_cascade_ ;
    wire \c0.n21_adj_2304 ;
    wire \c0.data_out_frame2_19_6 ;
    wire \c0.data_out_frame2_0_0 ;
    wire \c0.n16972_cascade_ ;
    wire data_out_frame2_11_2;
    wire \c0.n10_adj_2281 ;
    wire \c0.n17969 ;
    wire data_out_frame2_16_4;
    wire \c0.data_out_frame2_20_4 ;
    wire \c0.n17972_cascade_ ;
    wire \c0.n17040 ;
    wire \c0.n16972 ;
    wire \c0.n30_adj_2295 ;
    wire data_out_frame2_7_7;
    wire \c0.n5_adj_2351 ;
    wire data_out_frame2_11_3;
    wire \c0.n9695 ;
    wire \c0.n9695_cascade_ ;
    wire rand_data_22;
    wire data_out_frame2_11_7;
    wire data_out_frame2_11_5;
    wire \c0.n9919 ;
    wire \c0.n9901 ;
    wire \c0.n10_adj_2292 ;
    wire data_out_frame2_7_4;
    wire \c0.n9913 ;
    wire \c0.n17034 ;
    wire \c0.n17034_cascade_ ;
    wire \c0.n9688 ;
    wire data_out_frame2_12_1;
    wire \c0.n9688_cascade_ ;
    wire \c0.n6_adj_2325 ;
    wire data_out_frame2_11_1;
    wire data_out_frame2_6_1;
    wire \c0.n17115 ;
    wire rand_data_5;
    wire data_out_frame2_16_5;
    wire data_out_frame2_8_5;
    wire data_out_frame2_10_3;
    wire \c0.n20_adj_2252 ;
    wire \c0.n17322 ;
    wire \c0.n17323_cascade_ ;
    wire \c0.n18053 ;
    wire rand_data_16;
    wire data_out_frame2_9_1;
    wire \c0.n17921 ;
    wire \c0.n17924 ;
    wire data_out_frame2_18_7;
    wire \c0.data_out_frame2_19_7 ;
    wire \c0.n18059_cascade_ ;
    wire \c0.data_out_frame2_20_7 ;
    wire \c0.n18062_cascade_ ;
    wire data_out_frame2_11_4;
    wire data_out_frame2_17_7;
    wire data_out_frame2_14_0;
    wire \c0.n9853 ;
    wire \c0.n9589 ;
    wire \c0.n9853_cascade_ ;
    wire data_out_frame2_13_0;
    wire \c0.n17046 ;
    wire \c0.n17581 ;
    wire \c0.n10259 ;
    wire \c0.data_out_7_3 ;
    wire \c0.n8_adj_2153 ;
    wire \c0.n17070 ;
    wire \c0.n9737 ;
    wire \c0.n12_adj_2285 ;
    wire \c0.data_out_6_3 ;
    wire \c0.data_out_2_3 ;
    wire n2652;
    wire \c0.n5_adj_2350 ;
    wire \c0.n17546_cascade_ ;
    wire \c0.n17592 ;
    wire \c0.n18017_cascade_ ;
    wire \c0.n17593 ;
    wire \c0.n10_adj_2154 ;
    wire \c0.n18020_cascade_ ;
    wire byte_transmit_counter_3;
    wire \c0.n10_adj_2155 ;
    wire \c0.n10_adj_2268 ;
    wire \c0.data_out_8_3 ;
    wire data_out_8_4;
    wire \c0.data_out_9_1 ;
    wire data_out_3_4;
    wire \c0.n17591 ;
    wire rand_setpoint_16;
    wire n2547;
    wire UART_TRANSMITTER_state_2;
    wire \c0.data_out_5_3 ;
    wire \c0.data_out_5_4 ;
    wire \c0.n9783 ;
    wire data_out_frame2_10_6;
    wire data_out_frame2_5_4;
    wire \c0.n17495 ;
    wire data_out_frame2_9_6;
    wire \c0.n18047 ;
    wire \c0.n9859 ;
    wire data_out_frame2_13_2;
    wire \c0.n17133 ;
    wire \c0.n27_adj_2277 ;
    wire data_out_frame2_8_6;
    wire data_out_frame2_6_6;
    wire \c0.n18050 ;
    wire \c0.n9671 ;
    wire \c0.n17016 ;
    wire \c0.n6_adj_2293 ;
    wire \c0.n16960 ;
    wire \c0.n24_adj_2272 ;
    wire data_out_frame2_9_2;
    wire data_out_frame2_16_0;
    wire \c0.n9892 ;
    wire \c0.n20_adj_2205 ;
    wire \c0.n18071 ;
    wire \c0.n18074_cascade_ ;
    wire data_out_frame2_12_7;
    wire data_out_frame2_13_7;
    wire \c0.n18065_cascade_ ;
    wire \c0.n18068 ;
    wire data_out_frame2_14_6;
    wire data_out_frame2_12_6;
    wire \c0.n18005_cascade_ ;
    wire \c0.n18008 ;
    wire data_out_frame2_10_0;
    wire \c0.n17347 ;
    wire rand_data_18;
    wire data_out_frame2_6_2;
    wire data_out_frame2_15_6;
    wire data_out_frame2_7_6;
    wire \c0.n17127 ;
    wire data_out_frame2_8_7;
    wire data_out_frame2_11_6;
    wire data_out_frame2_14_7;
    wire rand_data_12;
    wire data_out_frame2_17_4;
    wire rand_data_23;
    wire data_out_frame2_6_7;
    wire rand_data_31;
    wire data_out_frame2_5_7;
    wire rand_data_15;
    wire data_out_frame2_9_7;
    wire data_out_frame2_9_5;
    wire \c0.n16926 ;
    wire rand_data_24;
    wire data_out_frame2_5_0;
    wire rand_data_25;
    wire data_out_frame2_6_5;
    wire data_out_frame2_5_5;
    wire \c0.n5_adj_2349_cascade_ ;
    wire \c0.n6_adj_2280 ;
    wire rand_data_13;
    wire \c0.n6_adj_2278 ;
    wire \c0.n18089 ;
    wire \c0.n17561 ;
    wire data_out_frame2_7_5;
    wire \c0.n9678 ;
    wire \c0.n18092 ;
    wire \c0.n22_adj_2352 ;
    wire \c0.tx2.r_Tx_Data_7 ;
    wire n4445;
    wire data_out_0_0;
    wire data_out_frame2_12_3;
    wire rand_data_29;
    wire data_out_frame2_13_5;
    wire \c0.data_out_5_1 ;
    wire \c0.n17043 ;
    wire \c0.n16949 ;
    wire data_out_8_7;
    wire \c0.data_out_7__3__N_441 ;
    wire \c0.n10_adj_2276 ;
    wire \c0.data_out_9_3 ;
    wire \c0.n16981 ;
    wire \c0.n16969 ;
    wire \c0.n6_adj_2274 ;
    wire \c0.data_out_9_4 ;
    wire \c0.data_out_10_4 ;
    wire \c0.data_out_7_2 ;
    wire \c0.n17058 ;
    wire \c0.n17028 ;
    wire \c0.n17058_cascade_ ;
    wire \c0.n17094 ;
    wire \c0.n19_adj_2283 ;
    wire \c0.n21_adj_2284_cascade_ ;
    wire \c0.n20_adj_2282 ;
    wire \c0.data_out_9_7 ;
    wire \c0.n17007 ;
    wire \c0.n9505 ;
    wire \c0.n17076 ;
    wire data_out_8_0;
    wire \c0.data_out_10_3 ;
    wire \c0.data_out_9_6 ;
    wire \c0.data_out_10_2 ;
    wire \c0.n16998 ;
    wire \c0.data_out_6_2 ;
    wire \c0.data_out_10_6 ;
    wire data_out_10__7__N_110;
    wire rand_setpoint_21;
    wire \c0.n17522 ;
    wire UART_TRANSMITTER_state_1;
    wire \c0.data_out_6_5 ;
    wire n10055;
    wire rand_setpoint_10;
    wire UART_TRANSMITTER_state_0;
    wire \c0.n17450 ;
    wire \c0.n17999 ;
    wire \c0.n8621 ;
    wire \c0.n18002 ;
    wire \c0.data_out_frame2_20_6 ;
    wire \c0.byte_transmit_counter2_2 ;
    wire \c0.n22_adj_2353 ;
    wire \c0.tx2.r_Tx_Data_6 ;
    wire \c0.n16915 ;
    wire \c0.n17082 ;
    wire \c0.n17118 ;
    wire \c0.n17019 ;
    wire \c0.n5_adj_2321 ;
    wire \c0.n18083 ;
    wire \c0.n6_adj_2290_cascade_ ;
    wire \c0.n18086 ;
    wire data_out_frame2_10_1;
    wire data_out_frame2_12_0;
    wire data_out_frame2_8_1;
    wire data_out_frame2_14_3;
    wire \c0.n9895_cascade_ ;
    wire data_out_frame2_15_1;
    wire \c0.n26_adj_2314 ;
    wire \c0.n25_adj_2316 ;
    wire \c0.n23_adj_2318_cascade_ ;
    wire \c0.n24_adj_2315 ;
    wire rand_data_14;
    wire data_out_frame2_17_6;
    wire \c0.data_out_frame2_19_3 ;
    wire \c0.n17945_cascade_ ;
    wire data_out_frame2_16_3;
    wire \c0.n17948 ;
    wire rand_data_30;
    wire data_out_frame2_5_6;
    wire rand_data_11;
    wire data_out_frame2_17_3;
    wire rand_data_8;
    wire \c0.data_out_frame2_0_6 ;
    wire \c0.byte_transmit_counter2_1 ;
    wire \c0.byte_transmit_counter2_0 ;
    wire \c0.n17563 ;
    wire rand_data_6;
    wire data_out_frame2_16_6;
    wire rand_data_3;
    wire data_out_frame2_18_3;
    wire data_out_frame2_15_5;
    wire data_out_frame2_11_0;
    wire data_out_frame2_13_6;
    wire \c0.n16923 ;
    wire data_out_frame2_13_1;
    wire \c0.n9910 ;
    wire \c0.n9826 ;
    wire \c0.data_out_frame2_0_7 ;
    wire \c0.n9910_cascade_ ;
    wire \c0.n9843 ;
    wire data_out_frame2_14_1;
    wire data_out_frame2_8_0;
    wire data_out_frame2_15_0;
    wire data_out_frame2_8_4;
    wire \c0.n16_adj_2327 ;
    wire data_out_frame2_12_2;
    wire \c0.n17_adj_2328_cascade_ ;
    wire \c0.n17010 ;
    wire \c0.data_out_frame2_19_1 ;
    wire data_out_frame2_15_7;
    wire \c0.n16940 ;
    wire \c0.data_out_7_0 ;
    wire data_out_6_0;
    wire byte_transmit_counter_2;
    wire \c0.n5_adj_2265_cascade_ ;
    wire \c0.byte_transmit_counter_1 ;
    wire \c0.n18095 ;
    wire \c0.data_out_6__1__N_537 ;
    wire \c0.byte_transmit_counter_0 ;
    wire \c0.n17632 ;
    wire \c0.byte_transmit_counter2_4 ;
    wire \c0.n15_adj_2356 ;
    wire \c0.byte_transmit_counter2_3 ;
    wire \c0.n22_adj_2355 ;
    wire \c0.tx2.r_Tx_Data_4 ;
    wire \c0.tx2.n8737 ;
    wire rand_data_7;
    wire n10197;
    wire data_out_frame2_16_7;
    wire CLK_c;
    wire _gnd_net_;

    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__52613),
            .DIN(N__52612),
            .DOUT(N__52611),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__52613),
            .PADOUT(N__52612),
            .PADIN(N__52611),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__17170),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__52604),
            .DIN(N__52603),
            .DOUT(N__52602),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__52604),
            .PADOUT(N__52603),
            .PADIN(N__52602),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rx_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_input_iopad.PULLUP=1'b1;
    IO_PAD rx_input_iopad (
            .OE(N__52595),
            .DIN(N__52594),
            .DOUT(N__52593),
            .PACKAGEPIN(PIN_2));
    defparam rx_input_preio.PIN_TYPE=6'b000000;
    defparam rx_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_input_preio (
            .PADOEN(N__52595),
            .PADOUT(N__52594),
            .PADIN(N__52593),
            .CLOCKENABLE(VCCG0),
            .DIN0(\c0.rx.r_Rx_Data_R ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__50505),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam tx2_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx2_output_iopad.PULLUP=1'b1;
    IO_PAD tx2_output_iopad (
            .OE(N__52586),
            .DIN(N__52585),
            .DOUT(N__52584),
            .PACKAGEPIN(PIN_3));
    defparam tx2_output_preio.PIN_TYPE=6'b101001;
    defparam tx2_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx2_output_preio (
            .PADOEN(N__52586),
            .PADOUT(N__52585),
            .PADIN(N__52584),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__28696),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__17155));
    defparam tx_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_output_iopad.PULLUP=1'b1;
    IO_PAD tx_output_iopad (
            .OE(N__52577),
            .DIN(N__52576),
            .DOUT(N__52575),
            .PACKAGEPIN(PIN_1));
    defparam tx_output_preio.PIN_TYPE=6'b101001;
    defparam tx_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_output_preio (
            .PADOEN(N__52577),
            .PADOUT(N__52576),
            .PADIN(N__52575),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__20074),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20191));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__52568),
            .DIN(N__52567),
            .DOUT(N__52566),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__52568),
            .PADOUT(N__52567),
            .PADIN(N__52566),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__13232 (
            .O(N__52549),
            .I(N__52545));
    InMux I__13231 (
            .O(N__52548),
            .I(N__52541));
    LocalMux I__13230 (
            .O(N__52545),
            .I(N__52538));
    InMux I__13229 (
            .O(N__52544),
            .I(N__52535));
    LocalMux I__13228 (
            .O(N__52541),
            .I(N__52532));
    Span4Mux_h I__13227 (
            .O(N__52538),
            .I(N__52527));
    LocalMux I__13226 (
            .O(N__52535),
            .I(N__52527));
    Span4Mux_h I__13225 (
            .O(N__52532),
            .I(N__52524));
    Span4Mux_h I__13224 (
            .O(N__52527),
            .I(N__52521));
    Span4Mux_h I__13223 (
            .O(N__52524),
            .I(N__52518));
    Odrv4 I__13222 (
            .O(N__52521),
            .I(\c0.data_out_7_0 ));
    Odrv4 I__13221 (
            .O(N__52518),
            .I(\c0.data_out_7_0 ));
    InMux I__13220 (
            .O(N__52513),
            .I(N__52508));
    InMux I__13219 (
            .O(N__52512),
            .I(N__52505));
    InMux I__13218 (
            .O(N__52511),
            .I(N__52502));
    LocalMux I__13217 (
            .O(N__52508),
            .I(N__52499));
    LocalMux I__13216 (
            .O(N__52505),
            .I(N__52494));
    LocalMux I__13215 (
            .O(N__52502),
            .I(N__52491));
    Span4Mux_h I__13214 (
            .O(N__52499),
            .I(N__52488));
    InMux I__13213 (
            .O(N__52498),
            .I(N__52483));
    InMux I__13212 (
            .O(N__52497),
            .I(N__52483));
    Span4Mux_v I__13211 (
            .O(N__52494),
            .I(N__52480));
    Span4Mux_h I__13210 (
            .O(N__52491),
            .I(N__52477));
    Sp12to4 I__13209 (
            .O(N__52488),
            .I(N__52474));
    LocalMux I__13208 (
            .O(N__52483),
            .I(data_out_6_0));
    Odrv4 I__13207 (
            .O(N__52480),
            .I(data_out_6_0));
    Odrv4 I__13206 (
            .O(N__52477),
            .I(data_out_6_0));
    Odrv12 I__13205 (
            .O(N__52474),
            .I(data_out_6_0));
    InMux I__13204 (
            .O(N__52465),
            .I(N__52448));
    InMux I__13203 (
            .O(N__52464),
            .I(N__52445));
    InMux I__13202 (
            .O(N__52463),
            .I(N__52438));
    InMux I__13201 (
            .O(N__52462),
            .I(N__52438));
    InMux I__13200 (
            .O(N__52461),
            .I(N__52438));
    InMux I__13199 (
            .O(N__52460),
            .I(N__52434));
    InMux I__13198 (
            .O(N__52459),
            .I(N__52429));
    InMux I__13197 (
            .O(N__52458),
            .I(N__52429));
    InMux I__13196 (
            .O(N__52457),
            .I(N__52426));
    InMux I__13195 (
            .O(N__52456),
            .I(N__52419));
    InMux I__13194 (
            .O(N__52455),
            .I(N__52419));
    InMux I__13193 (
            .O(N__52454),
            .I(N__52419));
    InMux I__13192 (
            .O(N__52453),
            .I(N__52416));
    InMux I__13191 (
            .O(N__52452),
            .I(N__52410));
    InMux I__13190 (
            .O(N__52451),
            .I(N__52410));
    LocalMux I__13189 (
            .O(N__52448),
            .I(N__52399));
    LocalMux I__13188 (
            .O(N__52445),
            .I(N__52399));
    LocalMux I__13187 (
            .O(N__52438),
            .I(N__52396));
    CascadeMux I__13186 (
            .O(N__52437),
            .I(N__52393));
    LocalMux I__13185 (
            .O(N__52434),
            .I(N__52388));
    LocalMux I__13184 (
            .O(N__52429),
            .I(N__52388));
    LocalMux I__13183 (
            .O(N__52426),
            .I(N__52385));
    LocalMux I__13182 (
            .O(N__52419),
            .I(N__52380));
    LocalMux I__13181 (
            .O(N__52416),
            .I(N__52380));
    InMux I__13180 (
            .O(N__52415),
            .I(N__52377));
    LocalMux I__13179 (
            .O(N__52410),
            .I(N__52374));
    InMux I__13178 (
            .O(N__52409),
            .I(N__52369));
    InMux I__13177 (
            .O(N__52408),
            .I(N__52369));
    InMux I__13176 (
            .O(N__52407),
            .I(N__52364));
    InMux I__13175 (
            .O(N__52406),
            .I(N__52364));
    InMux I__13174 (
            .O(N__52405),
            .I(N__52361));
    InMux I__13173 (
            .O(N__52404),
            .I(N__52358));
    Span4Mux_s2_v I__13172 (
            .O(N__52399),
            .I(N__52355));
    Span4Mux_v I__13171 (
            .O(N__52396),
            .I(N__52352));
    InMux I__13170 (
            .O(N__52393),
            .I(N__52348));
    Span4Mux_s2_v I__13169 (
            .O(N__52388),
            .I(N__52345));
    Span4Mux_v I__13168 (
            .O(N__52385),
            .I(N__52338));
    Span4Mux_s2_v I__13167 (
            .O(N__52380),
            .I(N__52338));
    LocalMux I__13166 (
            .O(N__52377),
            .I(N__52338));
    Span4Mux_h I__13165 (
            .O(N__52374),
            .I(N__52335));
    LocalMux I__13164 (
            .O(N__52369),
            .I(N__52322));
    LocalMux I__13163 (
            .O(N__52364),
            .I(N__52322));
    LocalMux I__13162 (
            .O(N__52361),
            .I(N__52322));
    LocalMux I__13161 (
            .O(N__52358),
            .I(N__52322));
    Sp12to4 I__13160 (
            .O(N__52355),
            .I(N__52322));
    Sp12to4 I__13159 (
            .O(N__52352),
            .I(N__52322));
    InMux I__13158 (
            .O(N__52351),
            .I(N__52319));
    LocalMux I__13157 (
            .O(N__52348),
            .I(byte_transmit_counter_2));
    Odrv4 I__13156 (
            .O(N__52345),
            .I(byte_transmit_counter_2));
    Odrv4 I__13155 (
            .O(N__52338),
            .I(byte_transmit_counter_2));
    Odrv4 I__13154 (
            .O(N__52335),
            .I(byte_transmit_counter_2));
    Odrv12 I__13153 (
            .O(N__52322),
            .I(byte_transmit_counter_2));
    LocalMux I__13152 (
            .O(N__52319),
            .I(byte_transmit_counter_2));
    CascadeMux I__13151 (
            .O(N__52306),
            .I(\c0.n5_adj_2265_cascade_ ));
    InMux I__13150 (
            .O(N__52303),
            .I(N__52297));
    InMux I__13149 (
            .O(N__52302),
            .I(N__52291));
    InMux I__13148 (
            .O(N__52301),
            .I(N__52285));
    CascadeMux I__13147 (
            .O(N__52300),
            .I(N__52282));
    LocalMux I__13146 (
            .O(N__52297),
            .I(N__52279));
    InMux I__13145 (
            .O(N__52296),
            .I(N__52272));
    InMux I__13144 (
            .O(N__52295),
            .I(N__52272));
    InMux I__13143 (
            .O(N__52294),
            .I(N__52272));
    LocalMux I__13142 (
            .O(N__52291),
            .I(N__52269));
    InMux I__13141 (
            .O(N__52290),
            .I(N__52266));
    InMux I__13140 (
            .O(N__52289),
            .I(N__52261));
    InMux I__13139 (
            .O(N__52288),
            .I(N__52258));
    LocalMux I__13138 (
            .O(N__52285),
            .I(N__52254));
    InMux I__13137 (
            .O(N__52282),
            .I(N__52251));
    Span4Mux_h I__13136 (
            .O(N__52279),
            .I(N__52246));
    LocalMux I__13135 (
            .O(N__52272),
            .I(N__52246));
    Span4Mux_v I__13134 (
            .O(N__52269),
            .I(N__52243));
    LocalMux I__13133 (
            .O(N__52266),
            .I(N__52240));
    InMux I__13132 (
            .O(N__52265),
            .I(N__52237));
    CascadeMux I__13131 (
            .O(N__52264),
            .I(N__52233));
    LocalMux I__13130 (
            .O(N__52261),
            .I(N__52227));
    LocalMux I__13129 (
            .O(N__52258),
            .I(N__52224));
    InMux I__13128 (
            .O(N__52257),
            .I(N__52221));
    Span4Mux_v I__13127 (
            .O(N__52254),
            .I(N__52216));
    LocalMux I__13126 (
            .O(N__52251),
            .I(N__52216));
    Span4Mux_v I__13125 (
            .O(N__52246),
            .I(N__52213));
    Span4Mux_h I__13124 (
            .O(N__52243),
            .I(N__52208));
    Span4Mux_v I__13123 (
            .O(N__52240),
            .I(N__52208));
    LocalMux I__13122 (
            .O(N__52237),
            .I(N__52205));
    CascadeMux I__13121 (
            .O(N__52236),
            .I(N__52202));
    InMux I__13120 (
            .O(N__52233),
            .I(N__52197));
    InMux I__13119 (
            .O(N__52232),
            .I(N__52197));
    InMux I__13118 (
            .O(N__52231),
            .I(N__52192));
    InMux I__13117 (
            .O(N__52230),
            .I(N__52192));
    Span4Mux_v I__13116 (
            .O(N__52227),
            .I(N__52187));
    Span4Mux_v I__13115 (
            .O(N__52224),
            .I(N__52187));
    LocalMux I__13114 (
            .O(N__52221),
            .I(N__52176));
    Sp12to4 I__13113 (
            .O(N__52216),
            .I(N__52176));
    Sp12to4 I__13112 (
            .O(N__52213),
            .I(N__52176));
    Sp12to4 I__13111 (
            .O(N__52208),
            .I(N__52176));
    Span12Mux_s4_v I__13110 (
            .O(N__52205),
            .I(N__52176));
    InMux I__13109 (
            .O(N__52202),
            .I(N__52172));
    LocalMux I__13108 (
            .O(N__52197),
            .I(N__52165));
    LocalMux I__13107 (
            .O(N__52192),
            .I(N__52165));
    Sp12to4 I__13106 (
            .O(N__52187),
            .I(N__52165));
    Span12Mux_h I__13105 (
            .O(N__52176),
            .I(N__52162));
    InMux I__13104 (
            .O(N__52175),
            .I(N__52159));
    LocalMux I__13103 (
            .O(N__52172),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv12 I__13102 (
            .O(N__52165),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv12 I__13101 (
            .O(N__52162),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__13100 (
            .O(N__52159),
            .I(\c0.byte_transmit_counter_1 ));
    InMux I__13099 (
            .O(N__52150),
            .I(N__52147));
    LocalMux I__13098 (
            .O(N__52147),
            .I(N__52144));
    Odrv12 I__13097 (
            .O(N__52144),
            .I(\c0.n18095 ));
    InMux I__13096 (
            .O(N__52141),
            .I(N__52137));
    InMux I__13095 (
            .O(N__52140),
            .I(N__52132));
    LocalMux I__13094 (
            .O(N__52137),
            .I(N__52128));
    InMux I__13093 (
            .O(N__52136),
            .I(N__52125));
    InMux I__13092 (
            .O(N__52135),
            .I(N__52122));
    LocalMux I__13091 (
            .O(N__52132),
            .I(N__52119));
    InMux I__13090 (
            .O(N__52131),
            .I(N__52116));
    Span4Mux_h I__13089 (
            .O(N__52128),
            .I(N__52113));
    LocalMux I__13088 (
            .O(N__52125),
            .I(N__52110));
    LocalMux I__13087 (
            .O(N__52122),
            .I(\c0.data_out_6__1__N_537 ));
    Odrv12 I__13086 (
            .O(N__52119),
            .I(\c0.data_out_6__1__N_537 ));
    LocalMux I__13085 (
            .O(N__52116),
            .I(\c0.data_out_6__1__N_537 ));
    Odrv4 I__13084 (
            .O(N__52113),
            .I(\c0.data_out_6__1__N_537 ));
    Odrv4 I__13083 (
            .O(N__52110),
            .I(\c0.data_out_6__1__N_537 ));
    InMux I__13082 (
            .O(N__52099),
            .I(N__52093));
    CascadeMux I__13081 (
            .O(N__52098),
            .I(N__52077));
    CascadeMux I__13080 (
            .O(N__52097),
            .I(N__52073));
    InMux I__13079 (
            .O(N__52096),
            .I(N__52067));
    LocalMux I__13078 (
            .O(N__52093),
            .I(N__52057));
    InMux I__13077 (
            .O(N__52092),
            .I(N__52045));
    InMux I__13076 (
            .O(N__52091),
            .I(N__52045));
    InMux I__13075 (
            .O(N__52090),
            .I(N__52045));
    InMux I__13074 (
            .O(N__52089),
            .I(N__52045));
    InMux I__13073 (
            .O(N__52088),
            .I(N__52035));
    InMux I__13072 (
            .O(N__52087),
            .I(N__52030));
    InMux I__13071 (
            .O(N__52086),
            .I(N__52030));
    InMux I__13070 (
            .O(N__52085),
            .I(N__52025));
    InMux I__13069 (
            .O(N__52084),
            .I(N__52025));
    InMux I__13068 (
            .O(N__52083),
            .I(N__52022));
    InMux I__13067 (
            .O(N__52082),
            .I(N__52019));
    CascadeMux I__13066 (
            .O(N__52081),
            .I(N__52016));
    InMux I__13065 (
            .O(N__52080),
            .I(N__52013));
    InMux I__13064 (
            .O(N__52077),
            .I(N__52010));
    InMux I__13063 (
            .O(N__52076),
            .I(N__52005));
    InMux I__13062 (
            .O(N__52073),
            .I(N__52005));
    InMux I__13061 (
            .O(N__52072),
            .I(N__51998));
    InMux I__13060 (
            .O(N__52071),
            .I(N__51998));
    InMux I__13059 (
            .O(N__52070),
            .I(N__51998));
    LocalMux I__13058 (
            .O(N__52067),
            .I(N__51990));
    InMux I__13057 (
            .O(N__52066),
            .I(N__51987));
    InMux I__13056 (
            .O(N__52065),
            .I(N__51984));
    InMux I__13055 (
            .O(N__52064),
            .I(N__51979));
    InMux I__13054 (
            .O(N__52063),
            .I(N__51979));
    InMux I__13053 (
            .O(N__52062),
            .I(N__51976));
    InMux I__13052 (
            .O(N__52061),
            .I(N__51973));
    InMux I__13051 (
            .O(N__52060),
            .I(N__51967));
    Span4Mux_v I__13050 (
            .O(N__52057),
            .I(N__51964));
    InMux I__13049 (
            .O(N__52056),
            .I(N__51957));
    InMux I__13048 (
            .O(N__52055),
            .I(N__51957));
    InMux I__13047 (
            .O(N__52054),
            .I(N__51957));
    LocalMux I__13046 (
            .O(N__52045),
            .I(N__51954));
    InMux I__13045 (
            .O(N__52044),
            .I(N__51951));
    InMux I__13044 (
            .O(N__52043),
            .I(N__51948));
    InMux I__13043 (
            .O(N__52042),
            .I(N__51939));
    InMux I__13042 (
            .O(N__52041),
            .I(N__51939));
    InMux I__13041 (
            .O(N__52040),
            .I(N__51939));
    InMux I__13040 (
            .O(N__52039),
            .I(N__51939));
    InMux I__13039 (
            .O(N__52038),
            .I(N__51935));
    LocalMux I__13038 (
            .O(N__52035),
            .I(N__51924));
    LocalMux I__13037 (
            .O(N__52030),
            .I(N__51924));
    LocalMux I__13036 (
            .O(N__52025),
            .I(N__51924));
    LocalMux I__13035 (
            .O(N__52022),
            .I(N__51924));
    LocalMux I__13034 (
            .O(N__52019),
            .I(N__51924));
    InMux I__13033 (
            .O(N__52016),
            .I(N__51921));
    LocalMux I__13032 (
            .O(N__52013),
            .I(N__51918));
    LocalMux I__13031 (
            .O(N__52010),
            .I(N__51913));
    LocalMux I__13030 (
            .O(N__52005),
            .I(N__51913));
    LocalMux I__13029 (
            .O(N__51998),
            .I(N__51910));
    InMux I__13028 (
            .O(N__51997),
            .I(N__51905));
    InMux I__13027 (
            .O(N__51996),
            .I(N__51905));
    InMux I__13026 (
            .O(N__51995),
            .I(N__51898));
    InMux I__13025 (
            .O(N__51994),
            .I(N__51898));
    InMux I__13024 (
            .O(N__51993),
            .I(N__51898));
    Span4Mux_v I__13023 (
            .O(N__51990),
            .I(N__51893));
    LocalMux I__13022 (
            .O(N__51987),
            .I(N__51893));
    LocalMux I__13021 (
            .O(N__51984),
            .I(N__51888));
    LocalMux I__13020 (
            .O(N__51979),
            .I(N__51888));
    LocalMux I__13019 (
            .O(N__51976),
            .I(N__51882));
    LocalMux I__13018 (
            .O(N__51973),
            .I(N__51882));
    InMux I__13017 (
            .O(N__51972),
            .I(N__51879));
    InMux I__13016 (
            .O(N__51971),
            .I(N__51874));
    InMux I__13015 (
            .O(N__51970),
            .I(N__51874));
    LocalMux I__13014 (
            .O(N__51967),
            .I(N__51871));
    Span4Mux_h I__13013 (
            .O(N__51964),
            .I(N__51864));
    LocalMux I__13012 (
            .O(N__51957),
            .I(N__51864));
    Span4Mux_v I__13011 (
            .O(N__51954),
            .I(N__51864));
    LocalMux I__13010 (
            .O(N__51951),
            .I(N__51857));
    LocalMux I__13009 (
            .O(N__51948),
            .I(N__51857));
    LocalMux I__13008 (
            .O(N__51939),
            .I(N__51857));
    InMux I__13007 (
            .O(N__51938),
            .I(N__51854));
    LocalMux I__13006 (
            .O(N__51935),
            .I(N__51851));
    Span4Mux_v I__13005 (
            .O(N__51924),
            .I(N__51846));
    LocalMux I__13004 (
            .O(N__51921),
            .I(N__51846));
    Span12Mux_h I__13003 (
            .O(N__51918),
            .I(N__51843));
    Span4Mux_v I__13002 (
            .O(N__51913),
            .I(N__51836));
    Span4Mux_h I__13001 (
            .O(N__51910),
            .I(N__51836));
    LocalMux I__13000 (
            .O(N__51905),
            .I(N__51836));
    LocalMux I__12999 (
            .O(N__51898),
            .I(N__51829));
    Span4Mux_h I__12998 (
            .O(N__51893),
            .I(N__51829));
    Span4Mux_v I__12997 (
            .O(N__51888),
            .I(N__51829));
    CascadeMux I__12996 (
            .O(N__51887),
            .I(N__51826));
    Span4Mux_h I__12995 (
            .O(N__51882),
            .I(N__51823));
    LocalMux I__12994 (
            .O(N__51879),
            .I(N__51812));
    LocalMux I__12993 (
            .O(N__51874),
            .I(N__51812));
    Span4Mux_s1_v I__12992 (
            .O(N__51871),
            .I(N__51812));
    Span4Mux_h I__12991 (
            .O(N__51864),
            .I(N__51812));
    Span4Mux_v I__12990 (
            .O(N__51857),
            .I(N__51812));
    LocalMux I__12989 (
            .O(N__51854),
            .I(N__51809));
    Span12Mux_h I__12988 (
            .O(N__51851),
            .I(N__51802));
    Sp12to4 I__12987 (
            .O(N__51846),
            .I(N__51802));
    Span12Mux_v I__12986 (
            .O(N__51843),
            .I(N__51802));
    Span4Mux_h I__12985 (
            .O(N__51836),
            .I(N__51797));
    Span4Mux_h I__12984 (
            .O(N__51829),
            .I(N__51797));
    InMux I__12983 (
            .O(N__51826),
            .I(N__51794));
    Odrv4 I__12982 (
            .O(N__51823),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__12981 (
            .O(N__51812),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv12 I__12980 (
            .O(N__51809),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv12 I__12979 (
            .O(N__51802),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__12978 (
            .O(N__51797),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__12977 (
            .O(N__51794),
            .I(\c0.byte_transmit_counter_0 ));
    InMux I__12976 (
            .O(N__51781),
            .I(N__51778));
    LocalMux I__12975 (
            .O(N__51778),
            .I(\c0.n17632 ));
    CascadeMux I__12974 (
            .O(N__51775),
            .I(N__51771));
    CascadeMux I__12973 (
            .O(N__51774),
            .I(N__51767));
    InMux I__12972 (
            .O(N__51771),
            .I(N__51764));
    InMux I__12971 (
            .O(N__51770),
            .I(N__51758));
    InMux I__12970 (
            .O(N__51767),
            .I(N__51755));
    LocalMux I__12969 (
            .O(N__51764),
            .I(N__51752));
    InMux I__12968 (
            .O(N__51763),
            .I(N__51749));
    InMux I__12967 (
            .O(N__51762),
            .I(N__51746));
    InMux I__12966 (
            .O(N__51761),
            .I(N__51743));
    LocalMux I__12965 (
            .O(N__51758),
            .I(N__51740));
    LocalMux I__12964 (
            .O(N__51755),
            .I(N__51733));
    Span4Mux_v I__12963 (
            .O(N__51752),
            .I(N__51733));
    LocalMux I__12962 (
            .O(N__51749),
            .I(N__51730));
    LocalMux I__12961 (
            .O(N__51746),
            .I(N__51727));
    LocalMux I__12960 (
            .O(N__51743),
            .I(N__51724));
    Span4Mux_h I__12959 (
            .O(N__51740),
            .I(N__51721));
    InMux I__12958 (
            .O(N__51739),
            .I(N__51718));
    InMux I__12957 (
            .O(N__51738),
            .I(N__51715));
    Span4Mux_v I__12956 (
            .O(N__51733),
            .I(N__51711));
    Span4Mux_v I__12955 (
            .O(N__51730),
            .I(N__51702));
    Span4Mux_v I__12954 (
            .O(N__51727),
            .I(N__51702));
    Span4Mux_v I__12953 (
            .O(N__51724),
            .I(N__51702));
    Span4Mux_h I__12952 (
            .O(N__51721),
            .I(N__51702));
    LocalMux I__12951 (
            .O(N__51718),
            .I(N__51698));
    LocalMux I__12950 (
            .O(N__51715),
            .I(N__51695));
    InMux I__12949 (
            .O(N__51714),
            .I(N__51692));
    Span4Mux_h I__12948 (
            .O(N__51711),
            .I(N__51689));
    Span4Mux_v I__12947 (
            .O(N__51702),
            .I(N__51686));
    InMux I__12946 (
            .O(N__51701),
            .I(N__51683));
    Odrv4 I__12945 (
            .O(N__51698),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv4 I__12944 (
            .O(N__51695),
            .I(\c0.byte_transmit_counter2_4 ));
    LocalMux I__12943 (
            .O(N__51692),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv4 I__12942 (
            .O(N__51689),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv4 I__12941 (
            .O(N__51686),
            .I(\c0.byte_transmit_counter2_4 ));
    LocalMux I__12940 (
            .O(N__51683),
            .I(\c0.byte_transmit_counter2_4 ));
    InMux I__12939 (
            .O(N__51670),
            .I(N__51667));
    LocalMux I__12938 (
            .O(N__51667),
            .I(N__51664));
    Span4Mux_h I__12937 (
            .O(N__51664),
            .I(N__51661));
    Span4Mux_h I__12936 (
            .O(N__51661),
            .I(N__51658));
    Odrv4 I__12935 (
            .O(N__51658),
            .I(\c0.n15_adj_2356 ));
    CascadeMux I__12934 (
            .O(N__51655),
            .I(N__51652));
    InMux I__12933 (
            .O(N__51652),
            .I(N__51648));
    InMux I__12932 (
            .O(N__51651),
            .I(N__51640));
    LocalMux I__12931 (
            .O(N__51648),
            .I(N__51637));
    InMux I__12930 (
            .O(N__51647),
            .I(N__51634));
    InMux I__12929 (
            .O(N__51646),
            .I(N__51626));
    InMux I__12928 (
            .O(N__51645),
            .I(N__51626));
    InMux I__12927 (
            .O(N__51644),
            .I(N__51623));
    InMux I__12926 (
            .O(N__51643),
            .I(N__51610));
    LocalMux I__12925 (
            .O(N__51640),
            .I(N__51601));
    Span4Mux_v I__12924 (
            .O(N__51637),
            .I(N__51601));
    LocalMux I__12923 (
            .O(N__51634),
            .I(N__51601));
    InMux I__12922 (
            .O(N__51633),
            .I(N__51594));
    InMux I__12921 (
            .O(N__51632),
            .I(N__51594));
    InMux I__12920 (
            .O(N__51631),
            .I(N__51594));
    LocalMux I__12919 (
            .O(N__51626),
            .I(N__51589));
    LocalMux I__12918 (
            .O(N__51623),
            .I(N__51589));
    InMux I__12917 (
            .O(N__51622),
            .I(N__51586));
    InMux I__12916 (
            .O(N__51621),
            .I(N__51583));
    InMux I__12915 (
            .O(N__51620),
            .I(N__51580));
    InMux I__12914 (
            .O(N__51619),
            .I(N__51577));
    InMux I__12913 (
            .O(N__51618),
            .I(N__51571));
    InMux I__12912 (
            .O(N__51617),
            .I(N__51571));
    InMux I__12911 (
            .O(N__51616),
            .I(N__51564));
    InMux I__12910 (
            .O(N__51615),
            .I(N__51564));
    InMux I__12909 (
            .O(N__51614),
            .I(N__51564));
    InMux I__12908 (
            .O(N__51613),
            .I(N__51561));
    LocalMux I__12907 (
            .O(N__51610),
            .I(N__51558));
    InMux I__12906 (
            .O(N__51609),
            .I(N__51553));
    InMux I__12905 (
            .O(N__51608),
            .I(N__51553));
    Span4Mux_v I__12904 (
            .O(N__51601),
            .I(N__51550));
    LocalMux I__12903 (
            .O(N__51594),
            .I(N__51545));
    Span4Mux_v I__12902 (
            .O(N__51589),
            .I(N__51545));
    LocalMux I__12901 (
            .O(N__51586),
            .I(N__51536));
    LocalMux I__12900 (
            .O(N__51583),
            .I(N__51536));
    LocalMux I__12899 (
            .O(N__51580),
            .I(N__51536));
    LocalMux I__12898 (
            .O(N__51577),
            .I(N__51536));
    InMux I__12897 (
            .O(N__51576),
            .I(N__51532));
    LocalMux I__12896 (
            .O(N__51571),
            .I(N__51525));
    LocalMux I__12895 (
            .O(N__51564),
            .I(N__51525));
    LocalMux I__12894 (
            .O(N__51561),
            .I(N__51525));
    Span4Mux_h I__12893 (
            .O(N__51558),
            .I(N__51522));
    LocalMux I__12892 (
            .O(N__51553),
            .I(N__51515));
    Span4Mux_h I__12891 (
            .O(N__51550),
            .I(N__51515));
    Span4Mux_v I__12890 (
            .O(N__51545),
            .I(N__51515));
    Span12Mux_v I__12889 (
            .O(N__51536),
            .I(N__51512));
    InMux I__12888 (
            .O(N__51535),
            .I(N__51509));
    LocalMux I__12887 (
            .O(N__51532),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv12 I__12886 (
            .O(N__51525),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv4 I__12885 (
            .O(N__51522),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv4 I__12884 (
            .O(N__51515),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv12 I__12883 (
            .O(N__51512),
            .I(\c0.byte_transmit_counter2_3 ));
    LocalMux I__12882 (
            .O(N__51509),
            .I(\c0.byte_transmit_counter2_3 ));
    InMux I__12881 (
            .O(N__51496),
            .I(N__51493));
    LocalMux I__12880 (
            .O(N__51493),
            .I(N__51490));
    Span4Mux_v I__12879 (
            .O(N__51490),
            .I(N__51487));
    Odrv4 I__12878 (
            .O(N__51487),
            .I(\c0.n22_adj_2355 ));
    CascadeMux I__12877 (
            .O(N__51484),
            .I(N__51481));
    InMux I__12876 (
            .O(N__51481),
            .I(N__51478));
    LocalMux I__12875 (
            .O(N__51478),
            .I(N__51475));
    Span4Mux_h I__12874 (
            .O(N__51475),
            .I(N__51472));
    Span4Mux_h I__12873 (
            .O(N__51472),
            .I(N__51469));
    Span4Mux_v I__12872 (
            .O(N__51469),
            .I(N__51466));
    Odrv4 I__12871 (
            .O(N__51466),
            .I(\c0.tx2.r_Tx_Data_4 ));
    CEMux I__12870 (
            .O(N__51463),
            .I(N__51459));
    CEMux I__12869 (
            .O(N__51462),
            .I(N__51456));
    LocalMux I__12868 (
            .O(N__51459),
            .I(N__51453));
    LocalMux I__12867 (
            .O(N__51456),
            .I(N__51448));
    Span4Mux_v I__12866 (
            .O(N__51453),
            .I(N__51443));
    CEMux I__12865 (
            .O(N__51452),
            .I(N__51440));
    CEMux I__12864 (
            .O(N__51451),
            .I(N__51437));
    Span4Mux_v I__12863 (
            .O(N__51448),
            .I(N__51434));
    CEMux I__12862 (
            .O(N__51447),
            .I(N__51431));
    CEMux I__12861 (
            .O(N__51446),
            .I(N__51428));
    Span4Mux_h I__12860 (
            .O(N__51443),
            .I(N__51423));
    LocalMux I__12859 (
            .O(N__51440),
            .I(N__51423));
    LocalMux I__12858 (
            .O(N__51437),
            .I(N__51420));
    Span4Mux_h I__12857 (
            .O(N__51434),
            .I(N__51415));
    LocalMux I__12856 (
            .O(N__51431),
            .I(N__51415));
    LocalMux I__12855 (
            .O(N__51428),
            .I(N__51412));
    Span4Mux_h I__12854 (
            .O(N__51423),
            .I(N__51408));
    Span4Mux_v I__12853 (
            .O(N__51420),
            .I(N__51405));
    Span4Mux_v I__12852 (
            .O(N__51415),
            .I(N__51401));
    Span4Mux_v I__12851 (
            .O(N__51412),
            .I(N__51398));
    CEMux I__12850 (
            .O(N__51411),
            .I(N__51395));
    Span4Mux_h I__12849 (
            .O(N__51408),
            .I(N__51390));
    Span4Mux_h I__12848 (
            .O(N__51405),
            .I(N__51390));
    CEMux I__12847 (
            .O(N__51404),
            .I(N__51387));
    Sp12to4 I__12846 (
            .O(N__51401),
            .I(N__51384));
    Span4Mux_h I__12845 (
            .O(N__51398),
            .I(N__51381));
    LocalMux I__12844 (
            .O(N__51395),
            .I(N__51378));
    Span4Mux_v I__12843 (
            .O(N__51390),
            .I(N__51373));
    LocalMux I__12842 (
            .O(N__51387),
            .I(N__51373));
    Span12Mux_h I__12841 (
            .O(N__51384),
            .I(N__51370));
    Span4Mux_h I__12840 (
            .O(N__51381),
            .I(N__51365));
    Span4Mux_h I__12839 (
            .O(N__51378),
            .I(N__51365));
    Span4Mux_h I__12838 (
            .O(N__51373),
            .I(N__51362));
    Span12Mux_v I__12837 (
            .O(N__51370),
            .I(N__51359));
    Span4Mux_h I__12836 (
            .O(N__51365),
            .I(N__51356));
    Span4Mux_h I__12835 (
            .O(N__51362),
            .I(N__51353));
    Odrv12 I__12834 (
            .O(N__51359),
            .I(\c0.tx2.n8737 ));
    Odrv4 I__12833 (
            .O(N__51356),
            .I(\c0.tx2.n8737 ));
    Odrv4 I__12832 (
            .O(N__51353),
            .I(\c0.tx2.n8737 ));
    InMux I__12831 (
            .O(N__51346),
            .I(N__51343));
    LocalMux I__12830 (
            .O(N__51343),
            .I(N__51340));
    Span4Mux_v I__12829 (
            .O(N__51340),
            .I(N__51335));
    InMux I__12828 (
            .O(N__51339),
            .I(N__51332));
    InMux I__12827 (
            .O(N__51338),
            .I(N__51329));
    Span4Mux_h I__12826 (
            .O(N__51335),
            .I(N__51322));
    LocalMux I__12825 (
            .O(N__51332),
            .I(N__51322));
    LocalMux I__12824 (
            .O(N__51329),
            .I(N__51319));
    InMux I__12823 (
            .O(N__51328),
            .I(N__51316));
    CascadeMux I__12822 (
            .O(N__51327),
            .I(N__51313));
    Span4Mux_v I__12821 (
            .O(N__51322),
            .I(N__51310));
    Span4Mux_h I__12820 (
            .O(N__51319),
            .I(N__51305));
    LocalMux I__12819 (
            .O(N__51316),
            .I(N__51305));
    InMux I__12818 (
            .O(N__51313),
            .I(N__51301));
    Span4Mux_h I__12817 (
            .O(N__51310),
            .I(N__51298));
    Span4Mux_h I__12816 (
            .O(N__51305),
            .I(N__51295));
    InMux I__12815 (
            .O(N__51304),
            .I(N__51292));
    LocalMux I__12814 (
            .O(N__51301),
            .I(N__51289));
    Odrv4 I__12813 (
            .O(N__51298),
            .I(rand_data_7));
    Odrv4 I__12812 (
            .O(N__51295),
            .I(rand_data_7));
    LocalMux I__12811 (
            .O(N__51292),
            .I(rand_data_7));
    Odrv12 I__12810 (
            .O(N__51289),
            .I(rand_data_7));
    InMux I__12809 (
            .O(N__51280),
            .I(N__51266));
    InMux I__12808 (
            .O(N__51279),
            .I(N__51266));
    InMux I__12807 (
            .O(N__51278),
            .I(N__51261));
    InMux I__12806 (
            .O(N__51277),
            .I(N__51261));
    InMux I__12805 (
            .O(N__51276),
            .I(N__51256));
    InMux I__12804 (
            .O(N__51275),
            .I(N__51256));
    InMux I__12803 (
            .O(N__51274),
            .I(N__51251));
    InMux I__12802 (
            .O(N__51273),
            .I(N__51251));
    InMux I__12801 (
            .O(N__51272),
            .I(N__51240));
    InMux I__12800 (
            .O(N__51271),
            .I(N__51237));
    LocalMux I__12799 (
            .O(N__51266),
            .I(N__51228));
    LocalMux I__12798 (
            .O(N__51261),
            .I(N__51228));
    LocalMux I__12797 (
            .O(N__51256),
            .I(N__51228));
    LocalMux I__12796 (
            .O(N__51251),
            .I(N__51228));
    InMux I__12795 (
            .O(N__51250),
            .I(N__51225));
    InMux I__12794 (
            .O(N__51249),
            .I(N__51174));
    CascadeMux I__12793 (
            .O(N__51248),
            .I(N__51171));
    CascadeMux I__12792 (
            .O(N__51247),
            .I(N__51165));
    CascadeMux I__12791 (
            .O(N__51246),
            .I(N__51162));
    InMux I__12790 (
            .O(N__51245),
            .I(N__51154));
    InMux I__12789 (
            .O(N__51244),
            .I(N__51154));
    InMux I__12788 (
            .O(N__51243),
            .I(N__51154));
    LocalMux I__12787 (
            .O(N__51240),
            .I(N__51151));
    LocalMux I__12786 (
            .O(N__51237),
            .I(N__51148));
    Span4Mux_v I__12785 (
            .O(N__51228),
            .I(N__51142));
    LocalMux I__12784 (
            .O(N__51225),
            .I(N__51142));
    InMux I__12783 (
            .O(N__51224),
            .I(N__51139));
    InMux I__12782 (
            .O(N__51223),
            .I(N__51132));
    InMux I__12781 (
            .O(N__51222),
            .I(N__51117));
    InMux I__12780 (
            .O(N__51221),
            .I(N__51117));
    InMux I__12779 (
            .O(N__51220),
            .I(N__51117));
    InMux I__12778 (
            .O(N__51219),
            .I(N__51117));
    InMux I__12777 (
            .O(N__51218),
            .I(N__51112));
    InMux I__12776 (
            .O(N__51217),
            .I(N__51112));
    CEMux I__12775 (
            .O(N__51216),
            .I(N__51109));
    CEMux I__12774 (
            .O(N__51215),
            .I(N__51106));
    InMux I__12773 (
            .O(N__51214),
            .I(N__51097));
    InMux I__12772 (
            .O(N__51213),
            .I(N__51097));
    InMux I__12771 (
            .O(N__51212),
            .I(N__51094));
    InMux I__12770 (
            .O(N__51211),
            .I(N__51089));
    InMux I__12769 (
            .O(N__51210),
            .I(N__51089));
    InMux I__12768 (
            .O(N__51209),
            .I(N__51084));
    InMux I__12767 (
            .O(N__51208),
            .I(N__51084));
    InMux I__12766 (
            .O(N__51207),
            .I(N__51081));
    InMux I__12765 (
            .O(N__51206),
            .I(N__51074));
    InMux I__12764 (
            .O(N__51205),
            .I(N__51074));
    InMux I__12763 (
            .O(N__51204),
            .I(N__51074));
    InMux I__12762 (
            .O(N__51203),
            .I(N__51066));
    InMux I__12761 (
            .O(N__51202),
            .I(N__51066));
    InMux I__12760 (
            .O(N__51201),
            .I(N__51066));
    InMux I__12759 (
            .O(N__51200),
            .I(N__51061));
    InMux I__12758 (
            .O(N__51199),
            .I(N__51061));
    InMux I__12757 (
            .O(N__51198),
            .I(N__51054));
    InMux I__12756 (
            .O(N__51197),
            .I(N__51054));
    InMux I__12755 (
            .O(N__51196),
            .I(N__51054));
    InMux I__12754 (
            .O(N__51195),
            .I(N__51043));
    InMux I__12753 (
            .O(N__51194),
            .I(N__51043));
    InMux I__12752 (
            .O(N__51193),
            .I(N__51043));
    InMux I__12751 (
            .O(N__51192),
            .I(N__51043));
    InMux I__12750 (
            .O(N__51191),
            .I(N__51043));
    InMux I__12749 (
            .O(N__51190),
            .I(N__51040));
    InMux I__12748 (
            .O(N__51189),
            .I(N__51033));
    InMux I__12747 (
            .O(N__51188),
            .I(N__51033));
    InMux I__12746 (
            .O(N__51187),
            .I(N__51033));
    InMux I__12745 (
            .O(N__51186),
            .I(N__51030));
    CEMux I__12744 (
            .O(N__51185),
            .I(N__51027));
    CEMux I__12743 (
            .O(N__51184),
            .I(N__51024));
    InMux I__12742 (
            .O(N__51183),
            .I(N__51021));
    CEMux I__12741 (
            .O(N__51182),
            .I(N__51018));
    CEMux I__12740 (
            .O(N__51181),
            .I(N__51015));
    InMux I__12739 (
            .O(N__51180),
            .I(N__51012));
    InMux I__12738 (
            .O(N__51179),
            .I(N__51005));
    InMux I__12737 (
            .O(N__51178),
            .I(N__51005));
    InMux I__12736 (
            .O(N__51177),
            .I(N__51005));
    LocalMux I__12735 (
            .O(N__51174),
            .I(N__51002));
    InMux I__12734 (
            .O(N__51171),
            .I(N__50996));
    InMux I__12733 (
            .O(N__51170),
            .I(N__50996));
    CEMux I__12732 (
            .O(N__51169),
            .I(N__50992));
    CEMux I__12731 (
            .O(N__51168),
            .I(N__50989));
    InMux I__12730 (
            .O(N__51165),
            .I(N__50982));
    InMux I__12729 (
            .O(N__51162),
            .I(N__50982));
    InMux I__12728 (
            .O(N__51161),
            .I(N__50982));
    LocalMux I__12727 (
            .O(N__51154),
            .I(N__50977));
    Span4Mux_v I__12726 (
            .O(N__51151),
            .I(N__50977));
    Span4Mux_h I__12725 (
            .O(N__51148),
            .I(N__50974));
    InMux I__12724 (
            .O(N__51147),
            .I(N__50971));
    Span4Mux_v I__12723 (
            .O(N__51142),
            .I(N__50966));
    LocalMux I__12722 (
            .O(N__51139),
            .I(N__50966));
    InMux I__12721 (
            .O(N__51138),
            .I(N__50956));
    InMux I__12720 (
            .O(N__51137),
            .I(N__50956));
    InMux I__12719 (
            .O(N__51136),
            .I(N__50956));
    InMux I__12718 (
            .O(N__51135),
            .I(N__50956));
    LocalMux I__12717 (
            .O(N__51132),
            .I(N__50953));
    InMux I__12716 (
            .O(N__51131),
            .I(N__50908));
    InMux I__12715 (
            .O(N__51130),
            .I(N__50908));
    InMux I__12714 (
            .O(N__51129),
            .I(N__50908));
    InMux I__12713 (
            .O(N__51128),
            .I(N__50908));
    InMux I__12712 (
            .O(N__51127),
            .I(N__50908));
    InMux I__12711 (
            .O(N__51126),
            .I(N__50908));
    LocalMux I__12710 (
            .O(N__51117),
            .I(N__50901));
    LocalMux I__12709 (
            .O(N__51112),
            .I(N__50901));
    LocalMux I__12708 (
            .O(N__51109),
            .I(N__50901));
    LocalMux I__12707 (
            .O(N__51106),
            .I(N__50898));
    InMux I__12706 (
            .O(N__51105),
            .I(N__50889));
    InMux I__12705 (
            .O(N__51104),
            .I(N__50889));
    InMux I__12704 (
            .O(N__51103),
            .I(N__50889));
    InMux I__12703 (
            .O(N__51102),
            .I(N__50889));
    LocalMux I__12702 (
            .O(N__51097),
            .I(N__50882));
    LocalMux I__12701 (
            .O(N__51094),
            .I(N__50882));
    LocalMux I__12700 (
            .O(N__51089),
            .I(N__50882));
    LocalMux I__12699 (
            .O(N__51084),
            .I(N__50879));
    LocalMux I__12698 (
            .O(N__51081),
            .I(N__50874));
    LocalMux I__12697 (
            .O(N__51074),
            .I(N__50874));
    InMux I__12696 (
            .O(N__51073),
            .I(N__50871));
    LocalMux I__12695 (
            .O(N__51066),
            .I(N__50866));
    LocalMux I__12694 (
            .O(N__51061),
            .I(N__50866));
    LocalMux I__12693 (
            .O(N__51054),
            .I(N__50863));
    LocalMux I__12692 (
            .O(N__51043),
            .I(N__50854));
    LocalMux I__12691 (
            .O(N__51040),
            .I(N__50854));
    LocalMux I__12690 (
            .O(N__51033),
            .I(N__50854));
    LocalMux I__12689 (
            .O(N__51030),
            .I(N__50854));
    LocalMux I__12688 (
            .O(N__51027),
            .I(N__50849));
    LocalMux I__12687 (
            .O(N__51024),
            .I(N__50849));
    LocalMux I__12686 (
            .O(N__51021),
            .I(N__50844));
    LocalMux I__12685 (
            .O(N__51018),
            .I(N__50844));
    LocalMux I__12684 (
            .O(N__51015),
            .I(N__50841));
    LocalMux I__12683 (
            .O(N__51012),
            .I(N__50834));
    LocalMux I__12682 (
            .O(N__51005),
            .I(N__50834));
    Span4Mux_h I__12681 (
            .O(N__51002),
            .I(N__50834));
    InMux I__12680 (
            .O(N__51001),
            .I(N__50831));
    LocalMux I__12679 (
            .O(N__50996),
            .I(N__50828));
    CEMux I__12678 (
            .O(N__50995),
            .I(N__50825));
    LocalMux I__12677 (
            .O(N__50992),
            .I(N__50822));
    LocalMux I__12676 (
            .O(N__50989),
            .I(N__50819));
    LocalMux I__12675 (
            .O(N__50982),
            .I(N__50812));
    Span4Mux_h I__12674 (
            .O(N__50977),
            .I(N__50812));
    Span4Mux_h I__12673 (
            .O(N__50974),
            .I(N__50812));
    LocalMux I__12672 (
            .O(N__50971),
            .I(N__50807));
    Span4Mux_h I__12671 (
            .O(N__50966),
            .I(N__50807));
    CEMux I__12670 (
            .O(N__50965),
            .I(N__50804));
    LocalMux I__12669 (
            .O(N__50956),
            .I(N__50799));
    Span4Mux_h I__12668 (
            .O(N__50953),
            .I(N__50799));
    InMux I__12667 (
            .O(N__50952),
            .I(N__50790));
    InMux I__12666 (
            .O(N__50951),
            .I(N__50790));
    InMux I__12665 (
            .O(N__50950),
            .I(N__50790));
    InMux I__12664 (
            .O(N__50949),
            .I(N__50790));
    InMux I__12663 (
            .O(N__50948),
            .I(N__50775));
    InMux I__12662 (
            .O(N__50947),
            .I(N__50775));
    InMux I__12661 (
            .O(N__50946),
            .I(N__50775));
    InMux I__12660 (
            .O(N__50945),
            .I(N__50775));
    InMux I__12659 (
            .O(N__50944),
            .I(N__50775));
    InMux I__12658 (
            .O(N__50943),
            .I(N__50775));
    InMux I__12657 (
            .O(N__50942),
            .I(N__50775));
    InMux I__12656 (
            .O(N__50941),
            .I(N__50764));
    InMux I__12655 (
            .O(N__50940),
            .I(N__50764));
    InMux I__12654 (
            .O(N__50939),
            .I(N__50764));
    InMux I__12653 (
            .O(N__50938),
            .I(N__50764));
    InMux I__12652 (
            .O(N__50937),
            .I(N__50764));
    InMux I__12651 (
            .O(N__50936),
            .I(N__50753));
    InMux I__12650 (
            .O(N__50935),
            .I(N__50753));
    InMux I__12649 (
            .O(N__50934),
            .I(N__50753));
    InMux I__12648 (
            .O(N__50933),
            .I(N__50753));
    InMux I__12647 (
            .O(N__50932),
            .I(N__50753));
    InMux I__12646 (
            .O(N__50931),
            .I(N__50744));
    InMux I__12645 (
            .O(N__50930),
            .I(N__50744));
    InMux I__12644 (
            .O(N__50929),
            .I(N__50744));
    InMux I__12643 (
            .O(N__50928),
            .I(N__50744));
    InMux I__12642 (
            .O(N__50927),
            .I(N__50737));
    InMux I__12641 (
            .O(N__50926),
            .I(N__50737));
    InMux I__12640 (
            .O(N__50925),
            .I(N__50737));
    InMux I__12639 (
            .O(N__50924),
            .I(N__50728));
    InMux I__12638 (
            .O(N__50923),
            .I(N__50728));
    InMux I__12637 (
            .O(N__50922),
            .I(N__50728));
    InMux I__12636 (
            .O(N__50921),
            .I(N__50728));
    LocalMux I__12635 (
            .O(N__50908),
            .I(N__50721));
    Span4Mux_v I__12634 (
            .O(N__50901),
            .I(N__50721));
    Span4Mux_v I__12633 (
            .O(N__50898),
            .I(N__50721));
    LocalMux I__12632 (
            .O(N__50889),
            .I(N__50712));
    Span4Mux_h I__12631 (
            .O(N__50882),
            .I(N__50712));
    Span4Mux_v I__12630 (
            .O(N__50879),
            .I(N__50712));
    Span4Mux_v I__12629 (
            .O(N__50874),
            .I(N__50712));
    LocalMux I__12628 (
            .O(N__50871),
            .I(N__50703));
    Span4Mux_v I__12627 (
            .O(N__50866),
            .I(N__50703));
    Span4Mux_v I__12626 (
            .O(N__50863),
            .I(N__50703));
    Span4Mux_v I__12625 (
            .O(N__50854),
            .I(N__50703));
    Span4Mux_v I__12624 (
            .O(N__50849),
            .I(N__50694));
    Span4Mux_v I__12623 (
            .O(N__50844),
            .I(N__50694));
    Span4Mux_v I__12622 (
            .O(N__50841),
            .I(N__50694));
    Span4Mux_h I__12621 (
            .O(N__50834),
            .I(N__50694));
    LocalMux I__12620 (
            .O(N__50831),
            .I(N__50689));
    Span4Mux_h I__12619 (
            .O(N__50828),
            .I(N__50689));
    LocalMux I__12618 (
            .O(N__50825),
            .I(N__50678));
    Span4Mux_h I__12617 (
            .O(N__50822),
            .I(N__50678));
    Span4Mux_v I__12616 (
            .O(N__50819),
            .I(N__50678));
    Span4Mux_v I__12615 (
            .O(N__50812),
            .I(N__50678));
    Span4Mux_h I__12614 (
            .O(N__50807),
            .I(N__50678));
    LocalMux I__12613 (
            .O(N__50804),
            .I(N__50673));
    Span4Mux_v I__12612 (
            .O(N__50799),
            .I(N__50673));
    LocalMux I__12611 (
            .O(N__50790),
            .I(n10197));
    LocalMux I__12610 (
            .O(N__50775),
            .I(n10197));
    LocalMux I__12609 (
            .O(N__50764),
            .I(n10197));
    LocalMux I__12608 (
            .O(N__50753),
            .I(n10197));
    LocalMux I__12607 (
            .O(N__50744),
            .I(n10197));
    LocalMux I__12606 (
            .O(N__50737),
            .I(n10197));
    LocalMux I__12605 (
            .O(N__50728),
            .I(n10197));
    Odrv4 I__12604 (
            .O(N__50721),
            .I(n10197));
    Odrv4 I__12603 (
            .O(N__50712),
            .I(n10197));
    Odrv4 I__12602 (
            .O(N__50703),
            .I(n10197));
    Odrv4 I__12601 (
            .O(N__50694),
            .I(n10197));
    Odrv4 I__12600 (
            .O(N__50689),
            .I(n10197));
    Odrv4 I__12599 (
            .O(N__50678),
            .I(n10197));
    Odrv4 I__12598 (
            .O(N__50673),
            .I(n10197));
    CascadeMux I__12597 (
            .O(N__50644),
            .I(N__50641));
    InMux I__12596 (
            .O(N__50641),
            .I(N__50638));
    LocalMux I__12595 (
            .O(N__50638),
            .I(N__50631));
    InMux I__12594 (
            .O(N__50637),
            .I(N__50628));
    InMux I__12593 (
            .O(N__50636),
            .I(N__50623));
    InMux I__12592 (
            .O(N__50635),
            .I(N__50623));
    InMux I__12591 (
            .O(N__50634),
            .I(N__50620));
    Span4Mux_h I__12590 (
            .O(N__50631),
            .I(N__50617));
    LocalMux I__12589 (
            .O(N__50628),
            .I(N__50614));
    LocalMux I__12588 (
            .O(N__50623),
            .I(N__50611));
    LocalMux I__12587 (
            .O(N__50620),
            .I(data_out_frame2_16_7));
    Odrv4 I__12586 (
            .O(N__50617),
            .I(data_out_frame2_16_7));
    Odrv12 I__12585 (
            .O(N__50614),
            .I(data_out_frame2_16_7));
    Odrv4 I__12584 (
            .O(N__50611),
            .I(data_out_frame2_16_7));
    ClkMux I__12583 (
            .O(N__50602),
            .I(N__49924));
    ClkMux I__12582 (
            .O(N__50601),
            .I(N__49924));
    ClkMux I__12581 (
            .O(N__50600),
            .I(N__49924));
    ClkMux I__12580 (
            .O(N__50599),
            .I(N__49924));
    ClkMux I__12579 (
            .O(N__50598),
            .I(N__49924));
    ClkMux I__12578 (
            .O(N__50597),
            .I(N__49924));
    ClkMux I__12577 (
            .O(N__50596),
            .I(N__49924));
    ClkMux I__12576 (
            .O(N__50595),
            .I(N__49924));
    ClkMux I__12575 (
            .O(N__50594),
            .I(N__49924));
    ClkMux I__12574 (
            .O(N__50593),
            .I(N__49924));
    ClkMux I__12573 (
            .O(N__50592),
            .I(N__49924));
    ClkMux I__12572 (
            .O(N__50591),
            .I(N__49924));
    ClkMux I__12571 (
            .O(N__50590),
            .I(N__49924));
    ClkMux I__12570 (
            .O(N__50589),
            .I(N__49924));
    ClkMux I__12569 (
            .O(N__50588),
            .I(N__49924));
    ClkMux I__12568 (
            .O(N__50587),
            .I(N__49924));
    ClkMux I__12567 (
            .O(N__50586),
            .I(N__49924));
    ClkMux I__12566 (
            .O(N__50585),
            .I(N__49924));
    ClkMux I__12565 (
            .O(N__50584),
            .I(N__49924));
    ClkMux I__12564 (
            .O(N__50583),
            .I(N__49924));
    ClkMux I__12563 (
            .O(N__50582),
            .I(N__49924));
    ClkMux I__12562 (
            .O(N__50581),
            .I(N__49924));
    ClkMux I__12561 (
            .O(N__50580),
            .I(N__49924));
    ClkMux I__12560 (
            .O(N__50579),
            .I(N__49924));
    ClkMux I__12559 (
            .O(N__50578),
            .I(N__49924));
    ClkMux I__12558 (
            .O(N__50577),
            .I(N__49924));
    ClkMux I__12557 (
            .O(N__50576),
            .I(N__49924));
    ClkMux I__12556 (
            .O(N__50575),
            .I(N__49924));
    ClkMux I__12555 (
            .O(N__50574),
            .I(N__49924));
    ClkMux I__12554 (
            .O(N__50573),
            .I(N__49924));
    ClkMux I__12553 (
            .O(N__50572),
            .I(N__49924));
    ClkMux I__12552 (
            .O(N__50571),
            .I(N__49924));
    ClkMux I__12551 (
            .O(N__50570),
            .I(N__49924));
    ClkMux I__12550 (
            .O(N__50569),
            .I(N__49924));
    ClkMux I__12549 (
            .O(N__50568),
            .I(N__49924));
    ClkMux I__12548 (
            .O(N__50567),
            .I(N__49924));
    ClkMux I__12547 (
            .O(N__50566),
            .I(N__49924));
    ClkMux I__12546 (
            .O(N__50565),
            .I(N__49924));
    ClkMux I__12545 (
            .O(N__50564),
            .I(N__49924));
    ClkMux I__12544 (
            .O(N__50563),
            .I(N__49924));
    ClkMux I__12543 (
            .O(N__50562),
            .I(N__49924));
    ClkMux I__12542 (
            .O(N__50561),
            .I(N__49924));
    ClkMux I__12541 (
            .O(N__50560),
            .I(N__49924));
    ClkMux I__12540 (
            .O(N__50559),
            .I(N__49924));
    ClkMux I__12539 (
            .O(N__50558),
            .I(N__49924));
    ClkMux I__12538 (
            .O(N__50557),
            .I(N__49924));
    ClkMux I__12537 (
            .O(N__50556),
            .I(N__49924));
    ClkMux I__12536 (
            .O(N__50555),
            .I(N__49924));
    ClkMux I__12535 (
            .O(N__50554),
            .I(N__49924));
    ClkMux I__12534 (
            .O(N__50553),
            .I(N__49924));
    ClkMux I__12533 (
            .O(N__50552),
            .I(N__49924));
    ClkMux I__12532 (
            .O(N__50551),
            .I(N__49924));
    ClkMux I__12531 (
            .O(N__50550),
            .I(N__49924));
    ClkMux I__12530 (
            .O(N__50549),
            .I(N__49924));
    ClkMux I__12529 (
            .O(N__50548),
            .I(N__49924));
    ClkMux I__12528 (
            .O(N__50547),
            .I(N__49924));
    ClkMux I__12527 (
            .O(N__50546),
            .I(N__49924));
    ClkMux I__12526 (
            .O(N__50545),
            .I(N__49924));
    ClkMux I__12525 (
            .O(N__50544),
            .I(N__49924));
    ClkMux I__12524 (
            .O(N__50543),
            .I(N__49924));
    ClkMux I__12523 (
            .O(N__50542),
            .I(N__49924));
    ClkMux I__12522 (
            .O(N__50541),
            .I(N__49924));
    ClkMux I__12521 (
            .O(N__50540),
            .I(N__49924));
    ClkMux I__12520 (
            .O(N__50539),
            .I(N__49924));
    ClkMux I__12519 (
            .O(N__50538),
            .I(N__49924));
    ClkMux I__12518 (
            .O(N__50537),
            .I(N__49924));
    ClkMux I__12517 (
            .O(N__50536),
            .I(N__49924));
    ClkMux I__12516 (
            .O(N__50535),
            .I(N__49924));
    ClkMux I__12515 (
            .O(N__50534),
            .I(N__49924));
    ClkMux I__12514 (
            .O(N__50533),
            .I(N__49924));
    ClkMux I__12513 (
            .O(N__50532),
            .I(N__49924));
    ClkMux I__12512 (
            .O(N__50531),
            .I(N__49924));
    ClkMux I__12511 (
            .O(N__50530),
            .I(N__49924));
    ClkMux I__12510 (
            .O(N__50529),
            .I(N__49924));
    ClkMux I__12509 (
            .O(N__50528),
            .I(N__49924));
    ClkMux I__12508 (
            .O(N__50527),
            .I(N__49924));
    ClkMux I__12507 (
            .O(N__50526),
            .I(N__49924));
    ClkMux I__12506 (
            .O(N__50525),
            .I(N__49924));
    ClkMux I__12505 (
            .O(N__50524),
            .I(N__49924));
    ClkMux I__12504 (
            .O(N__50523),
            .I(N__49924));
    ClkMux I__12503 (
            .O(N__50522),
            .I(N__49924));
    ClkMux I__12502 (
            .O(N__50521),
            .I(N__49924));
    ClkMux I__12501 (
            .O(N__50520),
            .I(N__49924));
    ClkMux I__12500 (
            .O(N__50519),
            .I(N__49924));
    ClkMux I__12499 (
            .O(N__50518),
            .I(N__49924));
    ClkMux I__12498 (
            .O(N__50517),
            .I(N__49924));
    ClkMux I__12497 (
            .O(N__50516),
            .I(N__49924));
    ClkMux I__12496 (
            .O(N__50515),
            .I(N__49924));
    ClkMux I__12495 (
            .O(N__50514),
            .I(N__49924));
    ClkMux I__12494 (
            .O(N__50513),
            .I(N__49924));
    ClkMux I__12493 (
            .O(N__50512),
            .I(N__49924));
    ClkMux I__12492 (
            .O(N__50511),
            .I(N__49924));
    ClkMux I__12491 (
            .O(N__50510),
            .I(N__49924));
    ClkMux I__12490 (
            .O(N__50509),
            .I(N__49924));
    ClkMux I__12489 (
            .O(N__50508),
            .I(N__49924));
    ClkMux I__12488 (
            .O(N__50507),
            .I(N__49924));
    ClkMux I__12487 (
            .O(N__50506),
            .I(N__49924));
    ClkMux I__12486 (
            .O(N__50505),
            .I(N__49924));
    ClkMux I__12485 (
            .O(N__50504),
            .I(N__49924));
    ClkMux I__12484 (
            .O(N__50503),
            .I(N__49924));
    ClkMux I__12483 (
            .O(N__50502),
            .I(N__49924));
    ClkMux I__12482 (
            .O(N__50501),
            .I(N__49924));
    ClkMux I__12481 (
            .O(N__50500),
            .I(N__49924));
    ClkMux I__12480 (
            .O(N__50499),
            .I(N__49924));
    ClkMux I__12479 (
            .O(N__50498),
            .I(N__49924));
    ClkMux I__12478 (
            .O(N__50497),
            .I(N__49924));
    ClkMux I__12477 (
            .O(N__50496),
            .I(N__49924));
    ClkMux I__12476 (
            .O(N__50495),
            .I(N__49924));
    ClkMux I__12475 (
            .O(N__50494),
            .I(N__49924));
    ClkMux I__12474 (
            .O(N__50493),
            .I(N__49924));
    ClkMux I__12473 (
            .O(N__50492),
            .I(N__49924));
    ClkMux I__12472 (
            .O(N__50491),
            .I(N__49924));
    ClkMux I__12471 (
            .O(N__50490),
            .I(N__49924));
    ClkMux I__12470 (
            .O(N__50489),
            .I(N__49924));
    ClkMux I__12469 (
            .O(N__50488),
            .I(N__49924));
    ClkMux I__12468 (
            .O(N__50487),
            .I(N__49924));
    ClkMux I__12467 (
            .O(N__50486),
            .I(N__49924));
    ClkMux I__12466 (
            .O(N__50485),
            .I(N__49924));
    ClkMux I__12465 (
            .O(N__50484),
            .I(N__49924));
    ClkMux I__12464 (
            .O(N__50483),
            .I(N__49924));
    ClkMux I__12463 (
            .O(N__50482),
            .I(N__49924));
    ClkMux I__12462 (
            .O(N__50481),
            .I(N__49924));
    ClkMux I__12461 (
            .O(N__50480),
            .I(N__49924));
    ClkMux I__12460 (
            .O(N__50479),
            .I(N__49924));
    ClkMux I__12459 (
            .O(N__50478),
            .I(N__49924));
    ClkMux I__12458 (
            .O(N__50477),
            .I(N__49924));
    ClkMux I__12457 (
            .O(N__50476),
            .I(N__49924));
    ClkMux I__12456 (
            .O(N__50475),
            .I(N__49924));
    ClkMux I__12455 (
            .O(N__50474),
            .I(N__49924));
    ClkMux I__12454 (
            .O(N__50473),
            .I(N__49924));
    ClkMux I__12453 (
            .O(N__50472),
            .I(N__49924));
    ClkMux I__12452 (
            .O(N__50471),
            .I(N__49924));
    ClkMux I__12451 (
            .O(N__50470),
            .I(N__49924));
    ClkMux I__12450 (
            .O(N__50469),
            .I(N__49924));
    ClkMux I__12449 (
            .O(N__50468),
            .I(N__49924));
    ClkMux I__12448 (
            .O(N__50467),
            .I(N__49924));
    ClkMux I__12447 (
            .O(N__50466),
            .I(N__49924));
    ClkMux I__12446 (
            .O(N__50465),
            .I(N__49924));
    ClkMux I__12445 (
            .O(N__50464),
            .I(N__49924));
    ClkMux I__12444 (
            .O(N__50463),
            .I(N__49924));
    ClkMux I__12443 (
            .O(N__50462),
            .I(N__49924));
    ClkMux I__12442 (
            .O(N__50461),
            .I(N__49924));
    ClkMux I__12441 (
            .O(N__50460),
            .I(N__49924));
    ClkMux I__12440 (
            .O(N__50459),
            .I(N__49924));
    ClkMux I__12439 (
            .O(N__50458),
            .I(N__49924));
    ClkMux I__12438 (
            .O(N__50457),
            .I(N__49924));
    ClkMux I__12437 (
            .O(N__50456),
            .I(N__49924));
    ClkMux I__12436 (
            .O(N__50455),
            .I(N__49924));
    ClkMux I__12435 (
            .O(N__50454),
            .I(N__49924));
    ClkMux I__12434 (
            .O(N__50453),
            .I(N__49924));
    ClkMux I__12433 (
            .O(N__50452),
            .I(N__49924));
    ClkMux I__12432 (
            .O(N__50451),
            .I(N__49924));
    ClkMux I__12431 (
            .O(N__50450),
            .I(N__49924));
    ClkMux I__12430 (
            .O(N__50449),
            .I(N__49924));
    ClkMux I__12429 (
            .O(N__50448),
            .I(N__49924));
    ClkMux I__12428 (
            .O(N__50447),
            .I(N__49924));
    ClkMux I__12427 (
            .O(N__50446),
            .I(N__49924));
    ClkMux I__12426 (
            .O(N__50445),
            .I(N__49924));
    ClkMux I__12425 (
            .O(N__50444),
            .I(N__49924));
    ClkMux I__12424 (
            .O(N__50443),
            .I(N__49924));
    ClkMux I__12423 (
            .O(N__50442),
            .I(N__49924));
    ClkMux I__12422 (
            .O(N__50441),
            .I(N__49924));
    ClkMux I__12421 (
            .O(N__50440),
            .I(N__49924));
    ClkMux I__12420 (
            .O(N__50439),
            .I(N__49924));
    ClkMux I__12419 (
            .O(N__50438),
            .I(N__49924));
    ClkMux I__12418 (
            .O(N__50437),
            .I(N__49924));
    ClkMux I__12417 (
            .O(N__50436),
            .I(N__49924));
    ClkMux I__12416 (
            .O(N__50435),
            .I(N__49924));
    ClkMux I__12415 (
            .O(N__50434),
            .I(N__49924));
    ClkMux I__12414 (
            .O(N__50433),
            .I(N__49924));
    ClkMux I__12413 (
            .O(N__50432),
            .I(N__49924));
    ClkMux I__12412 (
            .O(N__50431),
            .I(N__49924));
    ClkMux I__12411 (
            .O(N__50430),
            .I(N__49924));
    ClkMux I__12410 (
            .O(N__50429),
            .I(N__49924));
    ClkMux I__12409 (
            .O(N__50428),
            .I(N__49924));
    ClkMux I__12408 (
            .O(N__50427),
            .I(N__49924));
    ClkMux I__12407 (
            .O(N__50426),
            .I(N__49924));
    ClkMux I__12406 (
            .O(N__50425),
            .I(N__49924));
    ClkMux I__12405 (
            .O(N__50424),
            .I(N__49924));
    ClkMux I__12404 (
            .O(N__50423),
            .I(N__49924));
    ClkMux I__12403 (
            .O(N__50422),
            .I(N__49924));
    ClkMux I__12402 (
            .O(N__50421),
            .I(N__49924));
    ClkMux I__12401 (
            .O(N__50420),
            .I(N__49924));
    ClkMux I__12400 (
            .O(N__50419),
            .I(N__49924));
    ClkMux I__12399 (
            .O(N__50418),
            .I(N__49924));
    ClkMux I__12398 (
            .O(N__50417),
            .I(N__49924));
    ClkMux I__12397 (
            .O(N__50416),
            .I(N__49924));
    ClkMux I__12396 (
            .O(N__50415),
            .I(N__49924));
    ClkMux I__12395 (
            .O(N__50414),
            .I(N__49924));
    ClkMux I__12394 (
            .O(N__50413),
            .I(N__49924));
    ClkMux I__12393 (
            .O(N__50412),
            .I(N__49924));
    ClkMux I__12392 (
            .O(N__50411),
            .I(N__49924));
    ClkMux I__12391 (
            .O(N__50410),
            .I(N__49924));
    ClkMux I__12390 (
            .O(N__50409),
            .I(N__49924));
    ClkMux I__12389 (
            .O(N__50408),
            .I(N__49924));
    ClkMux I__12388 (
            .O(N__50407),
            .I(N__49924));
    ClkMux I__12387 (
            .O(N__50406),
            .I(N__49924));
    ClkMux I__12386 (
            .O(N__50405),
            .I(N__49924));
    ClkMux I__12385 (
            .O(N__50404),
            .I(N__49924));
    ClkMux I__12384 (
            .O(N__50403),
            .I(N__49924));
    ClkMux I__12383 (
            .O(N__50402),
            .I(N__49924));
    ClkMux I__12382 (
            .O(N__50401),
            .I(N__49924));
    ClkMux I__12381 (
            .O(N__50400),
            .I(N__49924));
    ClkMux I__12380 (
            .O(N__50399),
            .I(N__49924));
    ClkMux I__12379 (
            .O(N__50398),
            .I(N__49924));
    ClkMux I__12378 (
            .O(N__50397),
            .I(N__49924));
    ClkMux I__12377 (
            .O(N__50396),
            .I(N__49924));
    ClkMux I__12376 (
            .O(N__50395),
            .I(N__49924));
    ClkMux I__12375 (
            .O(N__50394),
            .I(N__49924));
    ClkMux I__12374 (
            .O(N__50393),
            .I(N__49924));
    ClkMux I__12373 (
            .O(N__50392),
            .I(N__49924));
    ClkMux I__12372 (
            .O(N__50391),
            .I(N__49924));
    ClkMux I__12371 (
            .O(N__50390),
            .I(N__49924));
    ClkMux I__12370 (
            .O(N__50389),
            .I(N__49924));
    ClkMux I__12369 (
            .O(N__50388),
            .I(N__49924));
    ClkMux I__12368 (
            .O(N__50387),
            .I(N__49924));
    ClkMux I__12367 (
            .O(N__50386),
            .I(N__49924));
    ClkMux I__12366 (
            .O(N__50385),
            .I(N__49924));
    ClkMux I__12365 (
            .O(N__50384),
            .I(N__49924));
    ClkMux I__12364 (
            .O(N__50383),
            .I(N__49924));
    ClkMux I__12363 (
            .O(N__50382),
            .I(N__49924));
    ClkMux I__12362 (
            .O(N__50381),
            .I(N__49924));
    ClkMux I__12361 (
            .O(N__50380),
            .I(N__49924));
    ClkMux I__12360 (
            .O(N__50379),
            .I(N__49924));
    ClkMux I__12359 (
            .O(N__50378),
            .I(N__49924));
    ClkMux I__12358 (
            .O(N__50377),
            .I(N__49924));
    GlobalMux I__12357 (
            .O(N__49924),
            .I(N__49921));
    gio2CtrlBuf I__12356 (
            .O(N__49921),
            .I(CLK_c));
    InMux I__12355 (
            .O(N__49918),
            .I(N__49913));
    InMux I__12354 (
            .O(N__49917),
            .I(N__49910));
    InMux I__12353 (
            .O(N__49916),
            .I(N__49907));
    LocalMux I__12352 (
            .O(N__49913),
            .I(N__49901));
    LocalMux I__12351 (
            .O(N__49910),
            .I(N__49901));
    LocalMux I__12350 (
            .O(N__49907),
            .I(N__49898));
    InMux I__12349 (
            .O(N__49906),
            .I(N__49894));
    Span4Mux_v I__12348 (
            .O(N__49901),
            .I(N__49891));
    Span4Mux_v I__12347 (
            .O(N__49898),
            .I(N__49888));
    InMux I__12346 (
            .O(N__49897),
            .I(N__49885));
    LocalMux I__12345 (
            .O(N__49894),
            .I(N__49882));
    Span4Mux_h I__12344 (
            .O(N__49891),
            .I(N__49879));
    Span4Mux_h I__12343 (
            .O(N__49888),
            .I(N__49873));
    LocalMux I__12342 (
            .O(N__49885),
            .I(N__49873));
    Span4Mux_h I__12341 (
            .O(N__49882),
            .I(N__49868));
    Span4Mux_h I__12340 (
            .O(N__49879),
            .I(N__49868));
    InMux I__12339 (
            .O(N__49878),
            .I(N__49865));
    Span4Mux_v I__12338 (
            .O(N__49873),
            .I(N__49862));
    Odrv4 I__12337 (
            .O(N__49868),
            .I(rand_data_6));
    LocalMux I__12336 (
            .O(N__49865),
            .I(rand_data_6));
    Odrv4 I__12335 (
            .O(N__49862),
            .I(rand_data_6));
    CascadeMux I__12334 (
            .O(N__49855),
            .I(N__49851));
    InMux I__12333 (
            .O(N__49854),
            .I(N__49848));
    InMux I__12332 (
            .O(N__49851),
            .I(N__49844));
    LocalMux I__12331 (
            .O(N__49848),
            .I(N__49840));
    InMux I__12330 (
            .O(N__49847),
            .I(N__49837));
    LocalMux I__12329 (
            .O(N__49844),
            .I(N__49834));
    InMux I__12328 (
            .O(N__49843),
            .I(N__49831));
    Span4Mux_v I__12327 (
            .O(N__49840),
            .I(N__49828));
    LocalMux I__12326 (
            .O(N__49837),
            .I(N__49825));
    Span4Mux_h I__12325 (
            .O(N__49834),
            .I(N__49822));
    LocalMux I__12324 (
            .O(N__49831),
            .I(data_out_frame2_16_6));
    Odrv4 I__12323 (
            .O(N__49828),
            .I(data_out_frame2_16_6));
    Odrv12 I__12322 (
            .O(N__49825),
            .I(data_out_frame2_16_6));
    Odrv4 I__12321 (
            .O(N__49822),
            .I(data_out_frame2_16_6));
    InMux I__12320 (
            .O(N__49813),
            .I(N__49810));
    LocalMux I__12319 (
            .O(N__49810),
            .I(N__49806));
    InMux I__12318 (
            .O(N__49809),
            .I(N__49803));
    Span4Mux_h I__12317 (
            .O(N__49806),
            .I(N__49796));
    LocalMux I__12316 (
            .O(N__49803),
            .I(N__49796));
    InMux I__12315 (
            .O(N__49802),
            .I(N__49793));
    InMux I__12314 (
            .O(N__49801),
            .I(N__49790));
    Span4Mux_v I__12313 (
            .O(N__49796),
            .I(N__49785));
    LocalMux I__12312 (
            .O(N__49793),
            .I(N__49785));
    LocalMux I__12311 (
            .O(N__49790),
            .I(N__49781));
    Span4Mux_h I__12310 (
            .O(N__49785),
            .I(N__49777));
    InMux I__12309 (
            .O(N__49784),
            .I(N__49774));
    Span12Mux_v I__12308 (
            .O(N__49781),
            .I(N__49771));
    InMux I__12307 (
            .O(N__49780),
            .I(N__49768));
    Sp12to4 I__12306 (
            .O(N__49777),
            .I(N__49763));
    LocalMux I__12305 (
            .O(N__49774),
            .I(N__49763));
    Odrv12 I__12304 (
            .O(N__49771),
            .I(rand_data_3));
    LocalMux I__12303 (
            .O(N__49768),
            .I(rand_data_3));
    Odrv12 I__12302 (
            .O(N__49763),
            .I(rand_data_3));
    InMux I__12301 (
            .O(N__49756),
            .I(N__49752));
    InMux I__12300 (
            .O(N__49755),
            .I(N__49749));
    LocalMux I__12299 (
            .O(N__49752),
            .I(data_out_frame2_18_3));
    LocalMux I__12298 (
            .O(N__49749),
            .I(data_out_frame2_18_3));
    CascadeMux I__12297 (
            .O(N__49744),
            .I(N__49739));
    InMux I__12296 (
            .O(N__49743),
            .I(N__49736));
    InMux I__12295 (
            .O(N__49742),
            .I(N__49732));
    InMux I__12294 (
            .O(N__49739),
            .I(N__49729));
    LocalMux I__12293 (
            .O(N__49736),
            .I(N__49726));
    InMux I__12292 (
            .O(N__49735),
            .I(N__49723));
    LocalMux I__12291 (
            .O(N__49732),
            .I(N__49720));
    LocalMux I__12290 (
            .O(N__49729),
            .I(N__49717));
    Span4Mux_v I__12289 (
            .O(N__49726),
            .I(N__49714));
    LocalMux I__12288 (
            .O(N__49723),
            .I(N__49707));
    Span4Mux_v I__12287 (
            .O(N__49720),
            .I(N__49707));
    Span4Mux_h I__12286 (
            .O(N__49717),
            .I(N__49707));
    Odrv4 I__12285 (
            .O(N__49714),
            .I(data_out_frame2_15_5));
    Odrv4 I__12284 (
            .O(N__49707),
            .I(data_out_frame2_15_5));
    InMux I__12283 (
            .O(N__49702),
            .I(N__49699));
    LocalMux I__12282 (
            .O(N__49699),
            .I(N__49695));
    InMux I__12281 (
            .O(N__49698),
            .I(N__49692));
    Span4Mux_h I__12280 (
            .O(N__49695),
            .I(N__49687));
    LocalMux I__12279 (
            .O(N__49692),
            .I(N__49687));
    Span4Mux_v I__12278 (
            .O(N__49687),
            .I(N__49681));
    InMux I__12277 (
            .O(N__49686),
            .I(N__49676));
    InMux I__12276 (
            .O(N__49685),
            .I(N__49676));
    InMux I__12275 (
            .O(N__49684),
            .I(N__49673));
    Span4Mux_h I__12274 (
            .O(N__49681),
            .I(N__49670));
    LocalMux I__12273 (
            .O(N__49676),
            .I(data_out_frame2_11_0));
    LocalMux I__12272 (
            .O(N__49673),
            .I(data_out_frame2_11_0));
    Odrv4 I__12271 (
            .O(N__49670),
            .I(data_out_frame2_11_0));
    InMux I__12270 (
            .O(N__49663),
            .I(N__49660));
    LocalMux I__12269 (
            .O(N__49660),
            .I(N__49655));
    InMux I__12268 (
            .O(N__49659),
            .I(N__49652));
    CascadeMux I__12267 (
            .O(N__49658),
            .I(N__49648));
    Span12Mux_s9_v I__12266 (
            .O(N__49655),
            .I(N__49643));
    LocalMux I__12265 (
            .O(N__49652),
            .I(N__49643));
    InMux I__12264 (
            .O(N__49651),
            .I(N__49638));
    InMux I__12263 (
            .O(N__49648),
            .I(N__49638));
    Odrv12 I__12262 (
            .O(N__49643),
            .I(data_out_frame2_13_6));
    LocalMux I__12261 (
            .O(N__49638),
            .I(data_out_frame2_13_6));
    InMux I__12260 (
            .O(N__49633),
            .I(N__49630));
    LocalMux I__12259 (
            .O(N__49630),
            .I(N__49626));
    InMux I__12258 (
            .O(N__49629),
            .I(N__49623));
    Span4Mux_h I__12257 (
            .O(N__49626),
            .I(N__49620));
    LocalMux I__12256 (
            .O(N__49623),
            .I(N__49617));
    Span4Mux_h I__12255 (
            .O(N__49620),
            .I(N__49614));
    Span4Mux_h I__12254 (
            .O(N__49617),
            .I(N__49611));
    Span4Mux_h I__12253 (
            .O(N__49614),
            .I(N__49608));
    Odrv4 I__12252 (
            .O(N__49611),
            .I(\c0.n16923 ));
    Odrv4 I__12251 (
            .O(N__49608),
            .I(\c0.n16923 ));
    CascadeMux I__12250 (
            .O(N__49603),
            .I(N__49600));
    InMux I__12249 (
            .O(N__49600),
            .I(N__49597));
    LocalMux I__12248 (
            .O(N__49597),
            .I(N__49592));
    InMux I__12247 (
            .O(N__49596),
            .I(N__49589));
    InMux I__12246 (
            .O(N__49595),
            .I(N__49586));
    Span12Mux_h I__12245 (
            .O(N__49592),
            .I(N__49583));
    LocalMux I__12244 (
            .O(N__49589),
            .I(data_out_frame2_13_1));
    LocalMux I__12243 (
            .O(N__49586),
            .I(data_out_frame2_13_1));
    Odrv12 I__12242 (
            .O(N__49583),
            .I(data_out_frame2_13_1));
    InMux I__12241 (
            .O(N__49576),
            .I(N__49573));
    LocalMux I__12240 (
            .O(N__49573),
            .I(N__49570));
    Span4Mux_h I__12239 (
            .O(N__49570),
            .I(N__49567));
    Odrv4 I__12238 (
            .O(N__49567),
            .I(\c0.n9910 ));
    InMux I__12237 (
            .O(N__49564),
            .I(N__49561));
    LocalMux I__12236 (
            .O(N__49561),
            .I(N__49558));
    Span4Mux_v I__12235 (
            .O(N__49558),
            .I(N__49554));
    InMux I__12234 (
            .O(N__49557),
            .I(N__49551));
    Span4Mux_v I__12233 (
            .O(N__49554),
            .I(N__49548));
    LocalMux I__12232 (
            .O(N__49551),
            .I(N__49545));
    Odrv4 I__12231 (
            .O(N__49548),
            .I(\c0.n9826 ));
    Odrv4 I__12230 (
            .O(N__49545),
            .I(\c0.n9826 ));
    InMux I__12229 (
            .O(N__49540),
            .I(N__49537));
    LocalMux I__12228 (
            .O(N__49537),
            .I(N__49532));
    InMux I__12227 (
            .O(N__49536),
            .I(N__49529));
    InMux I__12226 (
            .O(N__49535),
            .I(N__49526));
    Span4Mux_h I__12225 (
            .O(N__49532),
            .I(N__49518));
    LocalMux I__12224 (
            .O(N__49529),
            .I(N__49518));
    LocalMux I__12223 (
            .O(N__49526),
            .I(N__49518));
    InMux I__12222 (
            .O(N__49525),
            .I(N__49515));
    Span4Mux_h I__12221 (
            .O(N__49518),
            .I(N__49512));
    LocalMux I__12220 (
            .O(N__49515),
            .I(\c0.data_out_frame2_0_7 ));
    Odrv4 I__12219 (
            .O(N__49512),
            .I(\c0.data_out_frame2_0_7 ));
    CascadeMux I__12218 (
            .O(N__49507),
            .I(\c0.n9910_cascade_ ));
    InMux I__12217 (
            .O(N__49504),
            .I(N__49500));
    InMux I__12216 (
            .O(N__49503),
            .I(N__49497));
    LocalMux I__12215 (
            .O(N__49500),
            .I(N__49494));
    LocalMux I__12214 (
            .O(N__49497),
            .I(N__49491));
    Span4Mux_v I__12213 (
            .O(N__49494),
            .I(N__49488));
    Span4Mux_v I__12212 (
            .O(N__49491),
            .I(N__49485));
    Span4Mux_v I__12211 (
            .O(N__49488),
            .I(N__49480));
    Span4Mux_v I__12210 (
            .O(N__49485),
            .I(N__49480));
    Odrv4 I__12209 (
            .O(N__49480),
            .I(\c0.n9843 ));
    InMux I__12208 (
            .O(N__49477),
            .I(N__49473));
    CascadeMux I__12207 (
            .O(N__49476),
            .I(N__49470));
    LocalMux I__12206 (
            .O(N__49473),
            .I(N__49466));
    InMux I__12205 (
            .O(N__49470),
            .I(N__49463));
    CascadeMux I__12204 (
            .O(N__49469),
            .I(N__49460));
    Span4Mux_v I__12203 (
            .O(N__49466),
            .I(N__49456));
    LocalMux I__12202 (
            .O(N__49463),
            .I(N__49453));
    InMux I__12201 (
            .O(N__49460),
            .I(N__49450));
    InMux I__12200 (
            .O(N__49459),
            .I(N__49447));
    Span4Mux_h I__12199 (
            .O(N__49456),
            .I(N__49442));
    Span4Mux_v I__12198 (
            .O(N__49453),
            .I(N__49442));
    LocalMux I__12197 (
            .O(N__49450),
            .I(N__49439));
    LocalMux I__12196 (
            .O(N__49447),
            .I(data_out_frame2_14_1));
    Odrv4 I__12195 (
            .O(N__49442),
            .I(data_out_frame2_14_1));
    Odrv12 I__12194 (
            .O(N__49439),
            .I(data_out_frame2_14_1));
    InMux I__12193 (
            .O(N__49432),
            .I(N__49428));
    InMux I__12192 (
            .O(N__49431),
            .I(N__49424));
    LocalMux I__12191 (
            .O(N__49428),
            .I(N__49420));
    InMux I__12190 (
            .O(N__49427),
            .I(N__49417));
    LocalMux I__12189 (
            .O(N__49424),
            .I(N__49412));
    InMux I__12188 (
            .O(N__49423),
            .I(N__49409));
    Span4Mux_h I__12187 (
            .O(N__49420),
            .I(N__49406));
    LocalMux I__12186 (
            .O(N__49417),
            .I(N__49403));
    InMux I__12185 (
            .O(N__49416),
            .I(N__49398));
    InMux I__12184 (
            .O(N__49415),
            .I(N__49398));
    Span4Mux_h I__12183 (
            .O(N__49412),
            .I(N__49393));
    LocalMux I__12182 (
            .O(N__49409),
            .I(N__49393));
    Odrv4 I__12181 (
            .O(N__49406),
            .I(data_out_frame2_8_0));
    Odrv12 I__12180 (
            .O(N__49403),
            .I(data_out_frame2_8_0));
    LocalMux I__12179 (
            .O(N__49398),
            .I(data_out_frame2_8_0));
    Odrv4 I__12178 (
            .O(N__49393),
            .I(data_out_frame2_8_0));
    CascadeMux I__12177 (
            .O(N__49384),
            .I(N__49381));
    InMux I__12176 (
            .O(N__49381),
            .I(N__49375));
    InMux I__12175 (
            .O(N__49380),
            .I(N__49372));
    InMux I__12174 (
            .O(N__49379),
            .I(N__49369));
    CascadeMux I__12173 (
            .O(N__49378),
            .I(N__49366));
    LocalMux I__12172 (
            .O(N__49375),
            .I(N__49362));
    LocalMux I__12171 (
            .O(N__49372),
            .I(N__49357));
    LocalMux I__12170 (
            .O(N__49369),
            .I(N__49357));
    InMux I__12169 (
            .O(N__49366),
            .I(N__49352));
    InMux I__12168 (
            .O(N__49365),
            .I(N__49352));
    Odrv4 I__12167 (
            .O(N__49362),
            .I(data_out_frame2_15_0));
    Odrv12 I__12166 (
            .O(N__49357),
            .I(data_out_frame2_15_0));
    LocalMux I__12165 (
            .O(N__49352),
            .I(data_out_frame2_15_0));
    InMux I__12164 (
            .O(N__49345),
            .I(N__49340));
    InMux I__12163 (
            .O(N__49344),
            .I(N__49337));
    InMux I__12162 (
            .O(N__49343),
            .I(N__49334));
    LocalMux I__12161 (
            .O(N__49340),
            .I(N__49331));
    LocalMux I__12160 (
            .O(N__49337),
            .I(N__49328));
    LocalMux I__12159 (
            .O(N__49334),
            .I(N__49325));
    Span4Mux_h I__12158 (
            .O(N__49331),
            .I(N__49320));
    Span4Mux_v I__12157 (
            .O(N__49328),
            .I(N__49317));
    Span4Mux_h I__12156 (
            .O(N__49325),
            .I(N__49314));
    InMux I__12155 (
            .O(N__49324),
            .I(N__49309));
    InMux I__12154 (
            .O(N__49323),
            .I(N__49309));
    Odrv4 I__12153 (
            .O(N__49320),
            .I(data_out_frame2_8_4));
    Odrv4 I__12152 (
            .O(N__49317),
            .I(data_out_frame2_8_4));
    Odrv4 I__12151 (
            .O(N__49314),
            .I(data_out_frame2_8_4));
    LocalMux I__12150 (
            .O(N__49309),
            .I(data_out_frame2_8_4));
    InMux I__12149 (
            .O(N__49300),
            .I(N__49297));
    LocalMux I__12148 (
            .O(N__49297),
            .I(\c0.n16_adj_2327 ));
    InMux I__12147 (
            .O(N__49294),
            .I(N__49291));
    LocalMux I__12146 (
            .O(N__49291),
            .I(N__49287));
    CascadeMux I__12145 (
            .O(N__49290),
            .I(N__49284));
    Span4Mux_h I__12144 (
            .O(N__49287),
            .I(N__49280));
    InMux I__12143 (
            .O(N__49284),
            .I(N__49277));
    CascadeMux I__12142 (
            .O(N__49283),
            .I(N__49274));
    Span4Mux_h I__12141 (
            .O(N__49280),
            .I(N__49266));
    LocalMux I__12140 (
            .O(N__49277),
            .I(N__49266));
    InMux I__12139 (
            .O(N__49274),
            .I(N__49263));
    InMux I__12138 (
            .O(N__49273),
            .I(N__49260));
    InMux I__12137 (
            .O(N__49272),
            .I(N__49257));
    InMux I__12136 (
            .O(N__49271),
            .I(N__49254));
    Span4Mux_v I__12135 (
            .O(N__49266),
            .I(N__49251));
    LocalMux I__12134 (
            .O(N__49263),
            .I(N__49246));
    LocalMux I__12133 (
            .O(N__49260),
            .I(N__49246));
    LocalMux I__12132 (
            .O(N__49257),
            .I(data_out_frame2_12_2));
    LocalMux I__12131 (
            .O(N__49254),
            .I(data_out_frame2_12_2));
    Odrv4 I__12130 (
            .O(N__49251),
            .I(data_out_frame2_12_2));
    Odrv12 I__12129 (
            .O(N__49246),
            .I(data_out_frame2_12_2));
    CascadeMux I__12128 (
            .O(N__49237),
            .I(\c0.n17_adj_2328_cascade_ ));
    InMux I__12127 (
            .O(N__49234),
            .I(N__49231));
    LocalMux I__12126 (
            .O(N__49231),
            .I(N__49228));
    Span4Mux_h I__12125 (
            .O(N__49228),
            .I(N__49224));
    InMux I__12124 (
            .O(N__49227),
            .I(N__49221));
    Odrv4 I__12123 (
            .O(N__49224),
            .I(\c0.n17010 ));
    LocalMux I__12122 (
            .O(N__49221),
            .I(\c0.n17010 ));
    CascadeMux I__12121 (
            .O(N__49216),
            .I(N__49213));
    InMux I__12120 (
            .O(N__49213),
            .I(N__49210));
    LocalMux I__12119 (
            .O(N__49210),
            .I(N__49207));
    Span4Mux_h I__12118 (
            .O(N__49207),
            .I(N__49204));
    Span4Mux_h I__12117 (
            .O(N__49204),
            .I(N__49201));
    Odrv4 I__12116 (
            .O(N__49201),
            .I(\c0.data_out_frame2_19_1 ));
    InMux I__12115 (
            .O(N__49198),
            .I(N__49195));
    LocalMux I__12114 (
            .O(N__49195),
            .I(N__49191));
    InMux I__12113 (
            .O(N__49194),
            .I(N__49188));
    Span4Mux_h I__12112 (
            .O(N__49191),
            .I(N__49184));
    LocalMux I__12111 (
            .O(N__49188),
            .I(N__49179));
    InMux I__12110 (
            .O(N__49187),
            .I(N__49176));
    Span4Mux_v I__12109 (
            .O(N__49184),
            .I(N__49173));
    InMux I__12108 (
            .O(N__49183),
            .I(N__49168));
    InMux I__12107 (
            .O(N__49182),
            .I(N__49168));
    Span4Mux_h I__12106 (
            .O(N__49179),
            .I(N__49165));
    LocalMux I__12105 (
            .O(N__49176),
            .I(data_out_frame2_15_7));
    Odrv4 I__12104 (
            .O(N__49173),
            .I(data_out_frame2_15_7));
    LocalMux I__12103 (
            .O(N__49168),
            .I(data_out_frame2_15_7));
    Odrv4 I__12102 (
            .O(N__49165),
            .I(data_out_frame2_15_7));
    CascadeMux I__12101 (
            .O(N__49156),
            .I(N__49153));
    InMux I__12100 (
            .O(N__49153),
            .I(N__49150));
    LocalMux I__12099 (
            .O(N__49150),
            .I(N__49147));
    Odrv4 I__12098 (
            .O(N__49147),
            .I(\c0.n16940 ));
    InMux I__12097 (
            .O(N__49144),
            .I(N__49141));
    LocalMux I__12096 (
            .O(N__49141),
            .I(\c0.n26_adj_2314 ));
    InMux I__12095 (
            .O(N__49138),
            .I(N__49135));
    LocalMux I__12094 (
            .O(N__49135),
            .I(N__49132));
    Span4Mux_h I__12093 (
            .O(N__49132),
            .I(N__49129));
    Odrv4 I__12092 (
            .O(N__49129),
            .I(\c0.n25_adj_2316 ));
    CascadeMux I__12091 (
            .O(N__49126),
            .I(\c0.n23_adj_2318_cascade_ ));
    InMux I__12090 (
            .O(N__49123),
            .I(N__49120));
    LocalMux I__12089 (
            .O(N__49120),
            .I(N__49117));
    Span4Mux_v I__12088 (
            .O(N__49117),
            .I(N__49114));
    Odrv4 I__12087 (
            .O(N__49114),
            .I(\c0.n24_adj_2315 ));
    CascadeMux I__12086 (
            .O(N__49111),
            .I(N__49107));
    InMux I__12085 (
            .O(N__49110),
            .I(N__49103));
    InMux I__12084 (
            .O(N__49107),
            .I(N__49099));
    InMux I__12083 (
            .O(N__49106),
            .I(N__49096));
    LocalMux I__12082 (
            .O(N__49103),
            .I(N__49092));
    InMux I__12081 (
            .O(N__49102),
            .I(N__49089));
    LocalMux I__12080 (
            .O(N__49099),
            .I(N__49086));
    LocalMux I__12079 (
            .O(N__49096),
            .I(N__49083));
    InMux I__12078 (
            .O(N__49095),
            .I(N__49080));
    Span4Mux_h I__12077 (
            .O(N__49092),
            .I(N__49077));
    LocalMux I__12076 (
            .O(N__49089),
            .I(N__49074));
    Span4Mux_v I__12075 (
            .O(N__49086),
            .I(N__49068));
    Span4Mux_v I__12074 (
            .O(N__49083),
            .I(N__49068));
    LocalMux I__12073 (
            .O(N__49080),
            .I(N__49065));
    Span4Mux_h I__12072 (
            .O(N__49077),
            .I(N__49062));
    Span4Mux_h I__12071 (
            .O(N__49074),
            .I(N__49059));
    InMux I__12070 (
            .O(N__49073),
            .I(N__49056));
    Span4Mux_h I__12069 (
            .O(N__49068),
            .I(N__49051));
    Span4Mux_s3_v I__12068 (
            .O(N__49065),
            .I(N__49051));
    Odrv4 I__12067 (
            .O(N__49062),
            .I(rand_data_14));
    Odrv4 I__12066 (
            .O(N__49059),
            .I(rand_data_14));
    LocalMux I__12065 (
            .O(N__49056),
            .I(rand_data_14));
    Odrv4 I__12064 (
            .O(N__49051),
            .I(rand_data_14));
    CascadeMux I__12063 (
            .O(N__49042),
            .I(N__49039));
    InMux I__12062 (
            .O(N__49039),
            .I(N__49035));
    InMux I__12061 (
            .O(N__49038),
            .I(N__49032));
    LocalMux I__12060 (
            .O(N__49035),
            .I(N__49029));
    LocalMux I__12059 (
            .O(N__49032),
            .I(data_out_frame2_17_6));
    Odrv12 I__12058 (
            .O(N__49029),
            .I(data_out_frame2_17_6));
    InMux I__12057 (
            .O(N__49024),
            .I(N__49021));
    LocalMux I__12056 (
            .O(N__49021),
            .I(\c0.data_out_frame2_19_3 ));
    CascadeMux I__12055 (
            .O(N__49018),
            .I(\c0.n17945_cascade_ ));
    InMux I__12054 (
            .O(N__49015),
            .I(N__49012));
    LocalMux I__12053 (
            .O(N__49012),
            .I(N__49008));
    InMux I__12052 (
            .O(N__49011),
            .I(N__49004));
    Span4Mux_v I__12051 (
            .O(N__49008),
            .I(N__49000));
    InMux I__12050 (
            .O(N__49007),
            .I(N__48997));
    LocalMux I__12049 (
            .O(N__49004),
            .I(N__48994));
    InMux I__12048 (
            .O(N__49003),
            .I(N__48990));
    Span4Mux_h I__12047 (
            .O(N__49000),
            .I(N__48986));
    LocalMux I__12046 (
            .O(N__48997),
            .I(N__48981));
    Span4Mux_h I__12045 (
            .O(N__48994),
            .I(N__48981));
    InMux I__12044 (
            .O(N__48993),
            .I(N__48978));
    LocalMux I__12043 (
            .O(N__48990),
            .I(N__48975));
    InMux I__12042 (
            .O(N__48989),
            .I(N__48972));
    Span4Mux_h I__12041 (
            .O(N__48986),
            .I(N__48969));
    Span4Mux_h I__12040 (
            .O(N__48981),
            .I(N__48966));
    LocalMux I__12039 (
            .O(N__48978),
            .I(data_out_frame2_16_3));
    Odrv4 I__12038 (
            .O(N__48975),
            .I(data_out_frame2_16_3));
    LocalMux I__12037 (
            .O(N__48972),
            .I(data_out_frame2_16_3));
    Odrv4 I__12036 (
            .O(N__48969),
            .I(data_out_frame2_16_3));
    Odrv4 I__12035 (
            .O(N__48966),
            .I(data_out_frame2_16_3));
    InMux I__12034 (
            .O(N__48955),
            .I(N__48952));
    LocalMux I__12033 (
            .O(N__48952),
            .I(N__48949));
    Span4Mux_h I__12032 (
            .O(N__48949),
            .I(N__48946));
    Span4Mux_v I__12031 (
            .O(N__48946),
            .I(N__48943));
    Odrv4 I__12030 (
            .O(N__48943),
            .I(\c0.n17948 ));
    InMux I__12029 (
            .O(N__48940),
            .I(N__48937));
    LocalMux I__12028 (
            .O(N__48937),
            .I(N__48931));
    InMux I__12027 (
            .O(N__48936),
            .I(N__48928));
    InMux I__12026 (
            .O(N__48935),
            .I(N__48925));
    InMux I__12025 (
            .O(N__48934),
            .I(N__48922));
    Span4Mux_v I__12024 (
            .O(N__48931),
            .I(N__48919));
    LocalMux I__12023 (
            .O(N__48928),
            .I(N__48916));
    LocalMux I__12022 (
            .O(N__48925),
            .I(N__48913));
    LocalMux I__12021 (
            .O(N__48922),
            .I(N__48909));
    Span4Mux_h I__12020 (
            .O(N__48919),
            .I(N__48906));
    Span12Mux_v I__12019 (
            .O(N__48916),
            .I(N__48903));
    Span4Mux_v I__12018 (
            .O(N__48913),
            .I(N__48900));
    InMux I__12017 (
            .O(N__48912),
            .I(N__48897));
    Span4Mux_s1_v I__12016 (
            .O(N__48909),
            .I(N__48894));
    Odrv4 I__12015 (
            .O(N__48906),
            .I(rand_data_30));
    Odrv12 I__12014 (
            .O(N__48903),
            .I(rand_data_30));
    Odrv4 I__12013 (
            .O(N__48900),
            .I(rand_data_30));
    LocalMux I__12012 (
            .O(N__48897),
            .I(rand_data_30));
    Odrv4 I__12011 (
            .O(N__48894),
            .I(rand_data_30));
    InMux I__12010 (
            .O(N__48883),
            .I(N__48877));
    InMux I__12009 (
            .O(N__48882),
            .I(N__48877));
    LocalMux I__12008 (
            .O(N__48877),
            .I(N__48873));
    InMux I__12007 (
            .O(N__48876),
            .I(N__48869));
    Span4Mux_v I__12006 (
            .O(N__48873),
            .I(N__48866));
    InMux I__12005 (
            .O(N__48872),
            .I(N__48862));
    LocalMux I__12004 (
            .O(N__48869),
            .I(N__48859));
    Sp12to4 I__12003 (
            .O(N__48866),
            .I(N__48856));
    InMux I__12002 (
            .O(N__48865),
            .I(N__48853));
    LocalMux I__12001 (
            .O(N__48862),
            .I(data_out_frame2_5_6));
    Odrv4 I__12000 (
            .O(N__48859),
            .I(data_out_frame2_5_6));
    Odrv12 I__11999 (
            .O(N__48856),
            .I(data_out_frame2_5_6));
    LocalMux I__11998 (
            .O(N__48853),
            .I(data_out_frame2_5_6));
    InMux I__11997 (
            .O(N__48844),
            .I(N__48841));
    LocalMux I__11996 (
            .O(N__48841),
            .I(N__48836));
    InMux I__11995 (
            .O(N__48840),
            .I(N__48833));
    InMux I__11994 (
            .O(N__48839),
            .I(N__48830));
    Span4Mux_h I__11993 (
            .O(N__48836),
            .I(N__48825));
    LocalMux I__11992 (
            .O(N__48833),
            .I(N__48822));
    LocalMux I__11991 (
            .O(N__48830),
            .I(N__48819));
    InMux I__11990 (
            .O(N__48829),
            .I(N__48816));
    InMux I__11989 (
            .O(N__48828),
            .I(N__48812));
    Span4Mux_v I__11988 (
            .O(N__48825),
            .I(N__48809));
    Span12Mux_v I__11987 (
            .O(N__48822),
            .I(N__48806));
    Span4Mux_v I__11986 (
            .O(N__48819),
            .I(N__48803));
    LocalMux I__11985 (
            .O(N__48816),
            .I(N__48800));
    InMux I__11984 (
            .O(N__48815),
            .I(N__48797));
    LocalMux I__11983 (
            .O(N__48812),
            .I(N__48794));
    Odrv4 I__11982 (
            .O(N__48809),
            .I(rand_data_11));
    Odrv12 I__11981 (
            .O(N__48806),
            .I(rand_data_11));
    Odrv4 I__11980 (
            .O(N__48803),
            .I(rand_data_11));
    Odrv4 I__11979 (
            .O(N__48800),
            .I(rand_data_11));
    LocalMux I__11978 (
            .O(N__48797),
            .I(rand_data_11));
    Odrv12 I__11977 (
            .O(N__48794),
            .I(rand_data_11));
    InMux I__11976 (
            .O(N__48781),
            .I(N__48777));
    InMux I__11975 (
            .O(N__48780),
            .I(N__48774));
    LocalMux I__11974 (
            .O(N__48777),
            .I(data_out_frame2_17_3));
    LocalMux I__11973 (
            .O(N__48774),
            .I(data_out_frame2_17_3));
    InMux I__11972 (
            .O(N__48769),
            .I(N__48763));
    InMux I__11971 (
            .O(N__48768),
            .I(N__48760));
    InMux I__11970 (
            .O(N__48767),
            .I(N__48757));
    InMux I__11969 (
            .O(N__48766),
            .I(N__48754));
    LocalMux I__11968 (
            .O(N__48763),
            .I(N__48751));
    LocalMux I__11967 (
            .O(N__48760),
            .I(N__48748));
    LocalMux I__11966 (
            .O(N__48757),
            .I(N__48745));
    LocalMux I__11965 (
            .O(N__48754),
            .I(N__48741));
    Span4Mux_h I__11964 (
            .O(N__48751),
            .I(N__48738));
    Span4Mux_v I__11963 (
            .O(N__48748),
            .I(N__48733));
    Span4Mux_v I__11962 (
            .O(N__48745),
            .I(N__48733));
    InMux I__11961 (
            .O(N__48744),
            .I(N__48729));
    Span4Mux_v I__11960 (
            .O(N__48741),
            .I(N__48724));
    Span4Mux_h I__11959 (
            .O(N__48738),
            .I(N__48724));
    Span4Mux_h I__11958 (
            .O(N__48733),
            .I(N__48721));
    InMux I__11957 (
            .O(N__48732),
            .I(N__48718));
    LocalMux I__11956 (
            .O(N__48729),
            .I(N__48715));
    Odrv4 I__11955 (
            .O(N__48724),
            .I(rand_data_8));
    Odrv4 I__11954 (
            .O(N__48721),
            .I(rand_data_8));
    LocalMux I__11953 (
            .O(N__48718),
            .I(rand_data_8));
    Odrv12 I__11952 (
            .O(N__48715),
            .I(rand_data_8));
    InMux I__11951 (
            .O(N__48706),
            .I(N__48702));
    InMux I__11950 (
            .O(N__48705),
            .I(N__48698));
    LocalMux I__11949 (
            .O(N__48702),
            .I(N__48695));
    InMux I__11948 (
            .O(N__48701),
            .I(N__48691));
    LocalMux I__11947 (
            .O(N__48698),
            .I(N__48688));
    Span4Mux_h I__11946 (
            .O(N__48695),
            .I(N__48685));
    InMux I__11945 (
            .O(N__48694),
            .I(N__48682));
    LocalMux I__11944 (
            .O(N__48691),
            .I(N__48679));
    Span4Mux_h I__11943 (
            .O(N__48688),
            .I(N__48676));
    Odrv4 I__11942 (
            .O(N__48685),
            .I(\c0.data_out_frame2_0_6 ));
    LocalMux I__11941 (
            .O(N__48682),
            .I(\c0.data_out_frame2_0_6 ));
    Odrv12 I__11940 (
            .O(N__48679),
            .I(\c0.data_out_frame2_0_6 ));
    Odrv4 I__11939 (
            .O(N__48676),
            .I(\c0.data_out_frame2_0_6 ));
    InMux I__11938 (
            .O(N__48667),
            .I(N__48662));
    InMux I__11937 (
            .O(N__48666),
            .I(N__48659));
    InMux I__11936 (
            .O(N__48665),
            .I(N__48656));
    LocalMux I__11935 (
            .O(N__48662),
            .I(N__48642));
    LocalMux I__11934 (
            .O(N__48659),
            .I(N__48642));
    LocalMux I__11933 (
            .O(N__48656),
            .I(N__48642));
    InMux I__11932 (
            .O(N__48655),
            .I(N__48631));
    InMux I__11931 (
            .O(N__48654),
            .I(N__48631));
    CascadeMux I__11930 (
            .O(N__48653),
            .I(N__48626));
    InMux I__11929 (
            .O(N__48652),
            .I(N__48618));
    InMux I__11928 (
            .O(N__48651),
            .I(N__48618));
    InMux I__11927 (
            .O(N__48650),
            .I(N__48615));
    CascadeMux I__11926 (
            .O(N__48649),
            .I(N__48611));
    Span4Mux_v I__11925 (
            .O(N__48642),
            .I(N__48608));
    InMux I__11924 (
            .O(N__48641),
            .I(N__48605));
    InMux I__11923 (
            .O(N__48640),
            .I(N__48601));
    InMux I__11922 (
            .O(N__48639),
            .I(N__48596));
    InMux I__11921 (
            .O(N__48638),
            .I(N__48596));
    CascadeMux I__11920 (
            .O(N__48637),
            .I(N__48590));
    CascadeMux I__11919 (
            .O(N__48636),
            .I(N__48587));
    LocalMux I__11918 (
            .O(N__48631),
            .I(N__48575));
    InMux I__11917 (
            .O(N__48630),
            .I(N__48572));
    CascadeMux I__11916 (
            .O(N__48629),
            .I(N__48569));
    InMux I__11915 (
            .O(N__48626),
            .I(N__48565));
    InMux I__11914 (
            .O(N__48625),
            .I(N__48561));
    InMux I__11913 (
            .O(N__48624),
            .I(N__48558));
    InMux I__11912 (
            .O(N__48623),
            .I(N__48555));
    LocalMux I__11911 (
            .O(N__48618),
            .I(N__48552));
    LocalMux I__11910 (
            .O(N__48615),
            .I(N__48549));
    InMux I__11909 (
            .O(N__48614),
            .I(N__48546));
    InMux I__11908 (
            .O(N__48611),
            .I(N__48543));
    Span4Mux_h I__11907 (
            .O(N__48608),
            .I(N__48536));
    LocalMux I__11906 (
            .O(N__48605),
            .I(N__48536));
    InMux I__11905 (
            .O(N__48604),
            .I(N__48532));
    LocalMux I__11904 (
            .O(N__48601),
            .I(N__48527));
    LocalMux I__11903 (
            .O(N__48596),
            .I(N__48527));
    InMux I__11902 (
            .O(N__48595),
            .I(N__48524));
    InMux I__11901 (
            .O(N__48594),
            .I(N__48517));
    InMux I__11900 (
            .O(N__48593),
            .I(N__48517));
    InMux I__11899 (
            .O(N__48590),
            .I(N__48517));
    InMux I__11898 (
            .O(N__48587),
            .I(N__48514));
    InMux I__11897 (
            .O(N__48586),
            .I(N__48509));
    InMux I__11896 (
            .O(N__48585),
            .I(N__48506));
    InMux I__11895 (
            .O(N__48584),
            .I(N__48503));
    CascadeMux I__11894 (
            .O(N__48583),
            .I(N__48500));
    CascadeMux I__11893 (
            .O(N__48582),
            .I(N__48497));
    CascadeMux I__11892 (
            .O(N__48581),
            .I(N__48494));
    CascadeMux I__11891 (
            .O(N__48580),
            .I(N__48486));
    InMux I__11890 (
            .O(N__48579),
            .I(N__48481));
    InMux I__11889 (
            .O(N__48578),
            .I(N__48481));
    Span4Mux_v I__11888 (
            .O(N__48575),
            .I(N__48478));
    LocalMux I__11887 (
            .O(N__48572),
            .I(N__48475));
    InMux I__11886 (
            .O(N__48569),
            .I(N__48472));
    InMux I__11885 (
            .O(N__48568),
            .I(N__48469));
    LocalMux I__11884 (
            .O(N__48565),
            .I(N__48466));
    CascadeMux I__11883 (
            .O(N__48564),
            .I(N__48462));
    LocalMux I__11882 (
            .O(N__48561),
            .I(N__48453));
    LocalMux I__11881 (
            .O(N__48558),
            .I(N__48450));
    LocalMux I__11880 (
            .O(N__48555),
            .I(N__48447));
    Span4Mux_v I__11879 (
            .O(N__48552),
            .I(N__48438));
    Span4Mux_v I__11878 (
            .O(N__48549),
            .I(N__48438));
    LocalMux I__11877 (
            .O(N__48546),
            .I(N__48438));
    LocalMux I__11876 (
            .O(N__48543),
            .I(N__48438));
    InMux I__11875 (
            .O(N__48542),
            .I(N__48433));
    InMux I__11874 (
            .O(N__48541),
            .I(N__48433));
    Span4Mux_v I__11873 (
            .O(N__48536),
            .I(N__48430));
    InMux I__11872 (
            .O(N__48535),
            .I(N__48427));
    LocalMux I__11871 (
            .O(N__48532),
            .I(N__48418));
    Span4Mux_v I__11870 (
            .O(N__48527),
            .I(N__48418));
    LocalMux I__11869 (
            .O(N__48524),
            .I(N__48418));
    LocalMux I__11868 (
            .O(N__48517),
            .I(N__48418));
    LocalMux I__11867 (
            .O(N__48514),
            .I(N__48415));
    InMux I__11866 (
            .O(N__48513),
            .I(N__48412));
    InMux I__11865 (
            .O(N__48512),
            .I(N__48409));
    LocalMux I__11864 (
            .O(N__48509),
            .I(N__48402));
    LocalMux I__11863 (
            .O(N__48506),
            .I(N__48402));
    LocalMux I__11862 (
            .O(N__48503),
            .I(N__48402));
    InMux I__11861 (
            .O(N__48500),
            .I(N__48397));
    InMux I__11860 (
            .O(N__48497),
            .I(N__48397));
    InMux I__11859 (
            .O(N__48494),
            .I(N__48394));
    InMux I__11858 (
            .O(N__48493),
            .I(N__48388));
    InMux I__11857 (
            .O(N__48492),
            .I(N__48381));
    InMux I__11856 (
            .O(N__48491),
            .I(N__48381));
    InMux I__11855 (
            .O(N__48490),
            .I(N__48381));
    InMux I__11854 (
            .O(N__48489),
            .I(N__48378));
    InMux I__11853 (
            .O(N__48486),
            .I(N__48375));
    LocalMux I__11852 (
            .O(N__48481),
            .I(N__48372));
    Span4Mux_h I__11851 (
            .O(N__48478),
            .I(N__48365));
    Span4Mux_h I__11850 (
            .O(N__48475),
            .I(N__48365));
    LocalMux I__11849 (
            .O(N__48472),
            .I(N__48365));
    LocalMux I__11848 (
            .O(N__48469),
            .I(N__48360));
    Span4Mux_h I__11847 (
            .O(N__48466),
            .I(N__48360));
    InMux I__11846 (
            .O(N__48465),
            .I(N__48355));
    InMux I__11845 (
            .O(N__48462),
            .I(N__48355));
    InMux I__11844 (
            .O(N__48461),
            .I(N__48350));
    InMux I__11843 (
            .O(N__48460),
            .I(N__48341));
    InMux I__11842 (
            .O(N__48459),
            .I(N__48341));
    InMux I__11841 (
            .O(N__48458),
            .I(N__48341));
    InMux I__11840 (
            .O(N__48457),
            .I(N__48341));
    InMux I__11839 (
            .O(N__48456),
            .I(N__48338));
    Span4Mux_v I__11838 (
            .O(N__48453),
            .I(N__48331));
    Span4Mux_v I__11837 (
            .O(N__48450),
            .I(N__48331));
    Span4Mux_v I__11836 (
            .O(N__48447),
            .I(N__48331));
    Span4Mux_v I__11835 (
            .O(N__48438),
            .I(N__48328));
    LocalMux I__11834 (
            .O(N__48433),
            .I(N__48323));
    Span4Mux_v I__11833 (
            .O(N__48430),
            .I(N__48323));
    LocalMux I__11832 (
            .O(N__48427),
            .I(N__48318));
    Span4Mux_v I__11831 (
            .O(N__48418),
            .I(N__48318));
    Span4Mux_v I__11830 (
            .O(N__48415),
            .I(N__48315));
    LocalMux I__11829 (
            .O(N__48412),
            .I(N__48304));
    LocalMux I__11828 (
            .O(N__48409),
            .I(N__48304));
    Span4Mux_v I__11827 (
            .O(N__48402),
            .I(N__48304));
    LocalMux I__11826 (
            .O(N__48397),
            .I(N__48304));
    LocalMux I__11825 (
            .O(N__48394),
            .I(N__48304));
    InMux I__11824 (
            .O(N__48393),
            .I(N__48299));
    InMux I__11823 (
            .O(N__48392),
            .I(N__48299));
    InMux I__11822 (
            .O(N__48391),
            .I(N__48296));
    LocalMux I__11821 (
            .O(N__48388),
            .I(N__48279));
    LocalMux I__11820 (
            .O(N__48381),
            .I(N__48279));
    LocalMux I__11819 (
            .O(N__48378),
            .I(N__48279));
    LocalMux I__11818 (
            .O(N__48375),
            .I(N__48279));
    Span4Mux_h I__11817 (
            .O(N__48372),
            .I(N__48279));
    Span4Mux_v I__11816 (
            .O(N__48365),
            .I(N__48279));
    Span4Mux_h I__11815 (
            .O(N__48360),
            .I(N__48279));
    LocalMux I__11814 (
            .O(N__48355),
            .I(N__48279));
    InMux I__11813 (
            .O(N__48354),
            .I(N__48276));
    InMux I__11812 (
            .O(N__48353),
            .I(N__48273));
    LocalMux I__11811 (
            .O(N__48350),
            .I(N__48270));
    LocalMux I__11810 (
            .O(N__48341),
            .I(N__48265));
    LocalMux I__11809 (
            .O(N__48338),
            .I(N__48265));
    Span4Mux_h I__11808 (
            .O(N__48331),
            .I(N__48260));
    Span4Mux_h I__11807 (
            .O(N__48328),
            .I(N__48260));
    Span4Mux_v I__11806 (
            .O(N__48323),
            .I(N__48251));
    Span4Mux_h I__11805 (
            .O(N__48318),
            .I(N__48251));
    Span4Mux_h I__11804 (
            .O(N__48315),
            .I(N__48251));
    Span4Mux_v I__11803 (
            .O(N__48304),
            .I(N__48251));
    LocalMux I__11802 (
            .O(N__48299),
            .I(N__48244));
    LocalMux I__11801 (
            .O(N__48296),
            .I(N__48244));
    Sp12to4 I__11800 (
            .O(N__48279),
            .I(N__48244));
    LocalMux I__11799 (
            .O(N__48276),
            .I(\c0.byte_transmit_counter2_1 ));
    LocalMux I__11798 (
            .O(N__48273),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv12 I__11797 (
            .O(N__48270),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__11796 (
            .O(N__48265),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__11795 (
            .O(N__48260),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__11794 (
            .O(N__48251),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv12 I__11793 (
            .O(N__48244),
            .I(\c0.byte_transmit_counter2_1 ));
    InMux I__11792 (
            .O(N__48229),
            .I(N__48216));
    InMux I__11791 (
            .O(N__48228),
            .I(N__48216));
    InMux I__11790 (
            .O(N__48227),
            .I(N__48202));
    InMux I__11789 (
            .O(N__48226),
            .I(N__48202));
    InMux I__11788 (
            .O(N__48225),
            .I(N__48195));
    InMux I__11787 (
            .O(N__48224),
            .I(N__48195));
    InMux I__11786 (
            .O(N__48223),
            .I(N__48195));
    CascadeMux I__11785 (
            .O(N__48222),
            .I(N__48191));
    InMux I__11784 (
            .O(N__48221),
            .I(N__48183));
    LocalMux I__11783 (
            .O(N__48216),
            .I(N__48180));
    InMux I__11782 (
            .O(N__48215),
            .I(N__48177));
    InMux I__11781 (
            .O(N__48214),
            .I(N__48172));
    InMux I__11780 (
            .O(N__48213),
            .I(N__48172));
    InMux I__11779 (
            .O(N__48212),
            .I(N__48168));
    InMux I__11778 (
            .O(N__48211),
            .I(N__48161));
    InMux I__11777 (
            .O(N__48210),
            .I(N__48154));
    InMux I__11776 (
            .O(N__48209),
            .I(N__48154));
    InMux I__11775 (
            .O(N__48208),
            .I(N__48154));
    InMux I__11774 (
            .O(N__48207),
            .I(N__48151));
    LocalMux I__11773 (
            .O(N__48202),
            .I(N__48146));
    LocalMux I__11772 (
            .O(N__48195),
            .I(N__48146));
    InMux I__11771 (
            .O(N__48194),
            .I(N__48143));
    InMux I__11770 (
            .O(N__48191),
            .I(N__48137));
    InMux I__11769 (
            .O(N__48190),
            .I(N__48134));
    InMux I__11768 (
            .O(N__48189),
            .I(N__48131));
    InMux I__11767 (
            .O(N__48188),
            .I(N__48128));
    InMux I__11766 (
            .O(N__48187),
            .I(N__48125));
    InMux I__11765 (
            .O(N__48186),
            .I(N__48122));
    LocalMux I__11764 (
            .O(N__48183),
            .I(N__48111));
    Span4Mux_v I__11763 (
            .O(N__48180),
            .I(N__48111));
    LocalMux I__11762 (
            .O(N__48177),
            .I(N__48111));
    LocalMux I__11761 (
            .O(N__48172),
            .I(N__48111));
    InMux I__11760 (
            .O(N__48171),
            .I(N__48108));
    LocalMux I__11759 (
            .O(N__48168),
            .I(N__48101));
    InMux I__11758 (
            .O(N__48167),
            .I(N__48098));
    InMux I__11757 (
            .O(N__48166),
            .I(N__48093));
    InMux I__11756 (
            .O(N__48165),
            .I(N__48089));
    InMux I__11755 (
            .O(N__48164),
            .I(N__48086));
    LocalMux I__11754 (
            .O(N__48161),
            .I(N__48081));
    LocalMux I__11753 (
            .O(N__48154),
            .I(N__48081));
    LocalMux I__11752 (
            .O(N__48151),
            .I(N__48074));
    Span4Mux_v I__11751 (
            .O(N__48146),
            .I(N__48074));
    LocalMux I__11750 (
            .O(N__48143),
            .I(N__48074));
    InMux I__11749 (
            .O(N__48142),
            .I(N__48067));
    InMux I__11748 (
            .O(N__48141),
            .I(N__48067));
    InMux I__11747 (
            .O(N__48140),
            .I(N__48067));
    LocalMux I__11746 (
            .O(N__48137),
            .I(N__48060));
    LocalMux I__11745 (
            .O(N__48134),
            .I(N__48060));
    LocalMux I__11744 (
            .O(N__48131),
            .I(N__48053));
    LocalMux I__11743 (
            .O(N__48128),
            .I(N__48053));
    LocalMux I__11742 (
            .O(N__48125),
            .I(N__48053));
    LocalMux I__11741 (
            .O(N__48122),
            .I(N__48048));
    InMux I__11740 (
            .O(N__48121),
            .I(N__48045));
    InMux I__11739 (
            .O(N__48120),
            .I(N__48039));
    Span4Mux_v I__11738 (
            .O(N__48111),
            .I(N__48034));
    LocalMux I__11737 (
            .O(N__48108),
            .I(N__48034));
    InMux I__11736 (
            .O(N__48107),
            .I(N__48031));
    InMux I__11735 (
            .O(N__48106),
            .I(N__48027));
    InMux I__11734 (
            .O(N__48105),
            .I(N__48024));
    InMux I__11733 (
            .O(N__48104),
            .I(N__48021));
    Span4Mux_h I__11732 (
            .O(N__48101),
            .I(N__48016));
    LocalMux I__11731 (
            .O(N__48098),
            .I(N__48016));
    InMux I__11730 (
            .O(N__48097),
            .I(N__48013));
    CascadeMux I__11729 (
            .O(N__48096),
            .I(N__48010));
    LocalMux I__11728 (
            .O(N__48093),
            .I(N__48006));
    InMux I__11727 (
            .O(N__48092),
            .I(N__48003));
    LocalMux I__11726 (
            .O(N__48089),
            .I(N__47998));
    LocalMux I__11725 (
            .O(N__48086),
            .I(N__47998));
    Span4Mux_h I__11724 (
            .O(N__48081),
            .I(N__47991));
    Span4Mux_v I__11723 (
            .O(N__48074),
            .I(N__47991));
    LocalMux I__11722 (
            .O(N__48067),
            .I(N__47991));
    InMux I__11721 (
            .O(N__48066),
            .I(N__47988));
    InMux I__11720 (
            .O(N__48065),
            .I(N__47985));
    Span4Mux_h I__11719 (
            .O(N__48060),
            .I(N__47980));
    Span4Mux_v I__11718 (
            .O(N__48053),
            .I(N__47980));
    InMux I__11717 (
            .O(N__48052),
            .I(N__47977));
    InMux I__11716 (
            .O(N__48051),
            .I(N__47974));
    Span4Mux_h I__11715 (
            .O(N__48048),
            .I(N__47969));
    LocalMux I__11714 (
            .O(N__48045),
            .I(N__47969));
    InMux I__11713 (
            .O(N__48044),
            .I(N__47964));
    InMux I__11712 (
            .O(N__48043),
            .I(N__47964));
    InMux I__11711 (
            .O(N__48042),
            .I(N__47957));
    LocalMux I__11710 (
            .O(N__48039),
            .I(N__47954));
    Span4Mux_h I__11709 (
            .O(N__48034),
            .I(N__47949));
    LocalMux I__11708 (
            .O(N__48031),
            .I(N__47949));
    InMux I__11707 (
            .O(N__48030),
            .I(N__47946));
    LocalMux I__11706 (
            .O(N__48027),
            .I(N__47943));
    LocalMux I__11705 (
            .O(N__48024),
            .I(N__47938));
    LocalMux I__11704 (
            .O(N__48021),
            .I(N__47938));
    Span4Mux_v I__11703 (
            .O(N__48016),
            .I(N__47933));
    LocalMux I__11702 (
            .O(N__48013),
            .I(N__47933));
    InMux I__11701 (
            .O(N__48010),
            .I(N__47930));
    InMux I__11700 (
            .O(N__48009),
            .I(N__47927));
    Span4Mux_v I__11699 (
            .O(N__48006),
            .I(N__47924));
    LocalMux I__11698 (
            .O(N__48003),
            .I(N__47917));
    Span4Mux_v I__11697 (
            .O(N__47998),
            .I(N__47917));
    Span4Mux_h I__11696 (
            .O(N__47991),
            .I(N__47917));
    LocalMux I__11695 (
            .O(N__47988),
            .I(N__47910));
    LocalMux I__11694 (
            .O(N__47985),
            .I(N__47910));
    Span4Mux_h I__11693 (
            .O(N__47980),
            .I(N__47910));
    LocalMux I__11692 (
            .O(N__47977),
            .I(N__47901));
    LocalMux I__11691 (
            .O(N__47974),
            .I(N__47901));
    Span4Mux_v I__11690 (
            .O(N__47969),
            .I(N__47901));
    LocalMux I__11689 (
            .O(N__47964),
            .I(N__47901));
    InMux I__11688 (
            .O(N__47963),
            .I(N__47898));
    InMux I__11687 (
            .O(N__47962),
            .I(N__47895));
    InMux I__11686 (
            .O(N__47961),
            .I(N__47890));
    InMux I__11685 (
            .O(N__47960),
            .I(N__47890));
    LocalMux I__11684 (
            .O(N__47957),
            .I(N__47881));
    Span4Mux_h I__11683 (
            .O(N__47954),
            .I(N__47881));
    Span4Mux_v I__11682 (
            .O(N__47949),
            .I(N__47881));
    LocalMux I__11681 (
            .O(N__47946),
            .I(N__47881));
    Span4Mux_v I__11680 (
            .O(N__47943),
            .I(N__47874));
    Span4Mux_v I__11679 (
            .O(N__47938),
            .I(N__47874));
    Span4Mux_h I__11678 (
            .O(N__47933),
            .I(N__47874));
    LocalMux I__11677 (
            .O(N__47930),
            .I(N__47865));
    LocalMux I__11676 (
            .O(N__47927),
            .I(N__47865));
    Span4Mux_h I__11675 (
            .O(N__47924),
            .I(N__47865));
    Span4Mux_v I__11674 (
            .O(N__47917),
            .I(N__47865));
    Span4Mux_v I__11673 (
            .O(N__47910),
            .I(N__47860));
    Span4Mux_v I__11672 (
            .O(N__47901),
            .I(N__47860));
    LocalMux I__11671 (
            .O(N__47898),
            .I(N__47855));
    LocalMux I__11670 (
            .O(N__47895),
            .I(N__47855));
    LocalMux I__11669 (
            .O(N__47890),
            .I(N__47848));
    Span4Mux_v I__11668 (
            .O(N__47881),
            .I(N__47848));
    Span4Mux_h I__11667 (
            .O(N__47874),
            .I(N__47848));
    Odrv4 I__11666 (
            .O(N__47865),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__11665 (
            .O(N__47860),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv12 I__11664 (
            .O(N__47855),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__11663 (
            .O(N__47848),
            .I(\c0.byte_transmit_counter2_0 ));
    InMux I__11662 (
            .O(N__47839),
            .I(N__47836));
    LocalMux I__11661 (
            .O(N__47836),
            .I(N__47833));
    Odrv4 I__11660 (
            .O(N__47833),
            .I(\c0.n17563 ));
    InMux I__11659 (
            .O(N__47830),
            .I(N__47827));
    LocalMux I__11658 (
            .O(N__47827),
            .I(N__47824));
    Odrv4 I__11657 (
            .O(N__47824),
            .I(\c0.n17999 ));
    InMux I__11656 (
            .O(N__47821),
            .I(N__47818));
    LocalMux I__11655 (
            .O(N__47818),
            .I(N__47811));
    InMux I__11654 (
            .O(N__47817),
            .I(N__47808));
    InMux I__11653 (
            .O(N__47816),
            .I(N__47805));
    InMux I__11652 (
            .O(N__47815),
            .I(N__47801));
    InMux I__11651 (
            .O(N__47814),
            .I(N__47798));
    Span4Mux_h I__11650 (
            .O(N__47811),
            .I(N__47791));
    LocalMux I__11649 (
            .O(N__47808),
            .I(N__47791));
    LocalMux I__11648 (
            .O(N__47805),
            .I(N__47791));
    InMux I__11647 (
            .O(N__47804),
            .I(N__47788));
    LocalMux I__11646 (
            .O(N__47801),
            .I(N__47784));
    LocalMux I__11645 (
            .O(N__47798),
            .I(N__47781));
    Span4Mux_v I__11644 (
            .O(N__47791),
            .I(N__47776));
    LocalMux I__11643 (
            .O(N__47788),
            .I(N__47776));
    InMux I__11642 (
            .O(N__47787),
            .I(N__47773));
    Span4Mux_h I__11641 (
            .O(N__47784),
            .I(N__47770));
    Span4Mux_h I__11640 (
            .O(N__47781),
            .I(N__47767));
    Span4Mux_v I__11639 (
            .O(N__47776),
            .I(N__47762));
    LocalMux I__11638 (
            .O(N__47773),
            .I(N__47762));
    Span4Mux_h I__11637 (
            .O(N__47770),
            .I(N__47758));
    Span4Mux_v I__11636 (
            .O(N__47767),
            .I(N__47755));
    Span4Mux_h I__11635 (
            .O(N__47762),
            .I(N__47752));
    InMux I__11634 (
            .O(N__47761),
            .I(N__47749));
    Odrv4 I__11633 (
            .O(N__47758),
            .I(\c0.n8621 ));
    Odrv4 I__11632 (
            .O(N__47755),
            .I(\c0.n8621 ));
    Odrv4 I__11631 (
            .O(N__47752),
            .I(\c0.n8621 ));
    LocalMux I__11630 (
            .O(N__47749),
            .I(\c0.n8621 ));
    InMux I__11629 (
            .O(N__47740),
            .I(N__47737));
    LocalMux I__11628 (
            .O(N__47737),
            .I(\c0.n18002 ));
    CascadeMux I__11627 (
            .O(N__47734),
            .I(N__47731));
    InMux I__11626 (
            .O(N__47731),
            .I(N__47728));
    LocalMux I__11625 (
            .O(N__47728),
            .I(N__47725));
    Span4Mux_v I__11624 (
            .O(N__47725),
            .I(N__47722));
    Sp12to4 I__11623 (
            .O(N__47722),
            .I(N__47719));
    Odrv12 I__11622 (
            .O(N__47719),
            .I(\c0.data_out_frame2_20_6 ));
    InMux I__11621 (
            .O(N__47716),
            .I(N__47702));
    InMux I__11620 (
            .O(N__47715),
            .I(N__47699));
    InMux I__11619 (
            .O(N__47714),
            .I(N__47696));
    InMux I__11618 (
            .O(N__47713),
            .I(N__47693));
    InMux I__11617 (
            .O(N__47712),
            .I(N__47690));
    InMux I__11616 (
            .O(N__47711),
            .I(N__47687));
    InMux I__11615 (
            .O(N__47710),
            .I(N__47684));
    InMux I__11614 (
            .O(N__47709),
            .I(N__47681));
    InMux I__11613 (
            .O(N__47708),
            .I(N__47678));
    InMux I__11612 (
            .O(N__47707),
            .I(N__47675));
    InMux I__11611 (
            .O(N__47706),
            .I(N__47671));
    InMux I__11610 (
            .O(N__47705),
            .I(N__47668));
    LocalMux I__11609 (
            .O(N__47702),
            .I(N__47661));
    LocalMux I__11608 (
            .O(N__47699),
            .I(N__47661));
    LocalMux I__11607 (
            .O(N__47696),
            .I(N__47661));
    LocalMux I__11606 (
            .O(N__47693),
            .I(N__47651));
    LocalMux I__11605 (
            .O(N__47690),
            .I(N__47651));
    LocalMux I__11604 (
            .O(N__47687),
            .I(N__47651));
    LocalMux I__11603 (
            .O(N__47684),
            .I(N__47646));
    LocalMux I__11602 (
            .O(N__47681),
            .I(N__47646));
    LocalMux I__11601 (
            .O(N__47678),
            .I(N__47639));
    LocalMux I__11600 (
            .O(N__47675),
            .I(N__47636));
    InMux I__11599 (
            .O(N__47674),
            .I(N__47633));
    LocalMux I__11598 (
            .O(N__47671),
            .I(N__47624));
    LocalMux I__11597 (
            .O(N__47668),
            .I(N__47624));
    Span4Mux_v I__11596 (
            .O(N__47661),
            .I(N__47624));
    InMux I__11595 (
            .O(N__47660),
            .I(N__47621));
    InMux I__11594 (
            .O(N__47659),
            .I(N__47618));
    InMux I__11593 (
            .O(N__47658),
            .I(N__47615));
    Span4Mux_v I__11592 (
            .O(N__47651),
            .I(N__47612));
    Span4Mux_h I__11591 (
            .O(N__47646),
            .I(N__47609));
    InMux I__11590 (
            .O(N__47645),
            .I(N__47606));
    InMux I__11589 (
            .O(N__47644),
            .I(N__47601));
    InMux I__11588 (
            .O(N__47643),
            .I(N__47601));
    InMux I__11587 (
            .O(N__47642),
            .I(N__47598));
    Span4Mux_h I__11586 (
            .O(N__47639),
            .I(N__47595));
    Span4Mux_h I__11585 (
            .O(N__47636),
            .I(N__47590));
    LocalMux I__11584 (
            .O(N__47633),
            .I(N__47590));
    InMux I__11583 (
            .O(N__47632),
            .I(N__47587));
    InMux I__11582 (
            .O(N__47631),
            .I(N__47584));
    Span4Mux_h I__11581 (
            .O(N__47624),
            .I(N__47579));
    LocalMux I__11580 (
            .O(N__47621),
            .I(N__47579));
    LocalMux I__11579 (
            .O(N__47618),
            .I(N__47569));
    LocalMux I__11578 (
            .O(N__47615),
            .I(N__47569));
    Span4Mux_v I__11577 (
            .O(N__47612),
            .I(N__47569));
    Span4Mux_v I__11576 (
            .O(N__47609),
            .I(N__47569));
    LocalMux I__11575 (
            .O(N__47606),
            .I(N__47560));
    LocalMux I__11574 (
            .O(N__47601),
            .I(N__47560));
    LocalMux I__11573 (
            .O(N__47598),
            .I(N__47560));
    Span4Mux_h I__11572 (
            .O(N__47595),
            .I(N__47560));
    Span4Mux_h I__11571 (
            .O(N__47590),
            .I(N__47557));
    LocalMux I__11570 (
            .O(N__47587),
            .I(N__47550));
    LocalMux I__11569 (
            .O(N__47584),
            .I(N__47550));
    Sp12to4 I__11568 (
            .O(N__47579),
            .I(N__47550));
    InMux I__11567 (
            .O(N__47578),
            .I(N__47547));
    Odrv4 I__11566 (
            .O(N__47569),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv4 I__11565 (
            .O(N__47560),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv4 I__11564 (
            .O(N__47557),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv12 I__11563 (
            .O(N__47550),
            .I(\c0.byte_transmit_counter2_2 ));
    LocalMux I__11562 (
            .O(N__47547),
            .I(\c0.byte_transmit_counter2_2 ));
    InMux I__11561 (
            .O(N__47536),
            .I(N__47533));
    LocalMux I__11560 (
            .O(N__47533),
            .I(\c0.n22_adj_2353 ));
    InMux I__11559 (
            .O(N__47530),
            .I(N__47527));
    LocalMux I__11558 (
            .O(N__47527),
            .I(N__47524));
    Span12Mux_h I__11557 (
            .O(N__47524),
            .I(N__47521));
    Odrv12 I__11556 (
            .O(N__47521),
            .I(\c0.tx2.r_Tx_Data_6 ));
    InMux I__11555 (
            .O(N__47518),
            .I(N__47515));
    LocalMux I__11554 (
            .O(N__47515),
            .I(N__47512));
    Odrv4 I__11553 (
            .O(N__47512),
            .I(\c0.n16915 ));
    InMux I__11552 (
            .O(N__47509),
            .I(N__47506));
    LocalMux I__11551 (
            .O(N__47506),
            .I(N__47502));
    InMux I__11550 (
            .O(N__47505),
            .I(N__47499));
    Span4Mux_h I__11549 (
            .O(N__47502),
            .I(N__47496));
    LocalMux I__11548 (
            .O(N__47499),
            .I(N__47493));
    Odrv4 I__11547 (
            .O(N__47496),
            .I(\c0.n17082 ));
    Odrv4 I__11546 (
            .O(N__47493),
            .I(\c0.n17082 ));
    CascadeMux I__11545 (
            .O(N__47488),
            .I(N__47485));
    InMux I__11544 (
            .O(N__47485),
            .I(N__47481));
    CascadeMux I__11543 (
            .O(N__47484),
            .I(N__47478));
    LocalMux I__11542 (
            .O(N__47481),
            .I(N__47475));
    InMux I__11541 (
            .O(N__47478),
            .I(N__47472));
    Span4Mux_h I__11540 (
            .O(N__47475),
            .I(N__47467));
    LocalMux I__11539 (
            .O(N__47472),
            .I(N__47467));
    Span4Mux_h I__11538 (
            .O(N__47467),
            .I(N__47464));
    Span4Mux_h I__11537 (
            .O(N__47464),
            .I(N__47461));
    Odrv4 I__11536 (
            .O(N__47461),
            .I(\c0.n17118 ));
    InMux I__11535 (
            .O(N__47458),
            .I(N__47455));
    LocalMux I__11534 (
            .O(N__47455),
            .I(N__47452));
    Span4Mux_v I__11533 (
            .O(N__47452),
            .I(N__47448));
    InMux I__11532 (
            .O(N__47451),
            .I(N__47445));
    Odrv4 I__11531 (
            .O(N__47448),
            .I(\c0.n17019 ));
    LocalMux I__11530 (
            .O(N__47445),
            .I(\c0.n17019 ));
    CascadeMux I__11529 (
            .O(N__47440),
            .I(N__47437));
    InMux I__11528 (
            .O(N__47437),
            .I(N__47434));
    LocalMux I__11527 (
            .O(N__47434),
            .I(\c0.n5_adj_2321 ));
    InMux I__11526 (
            .O(N__47431),
            .I(N__47428));
    LocalMux I__11525 (
            .O(N__47428),
            .I(\c0.n18083 ));
    CascadeMux I__11524 (
            .O(N__47425),
            .I(\c0.n6_adj_2290_cascade_ ));
    InMux I__11523 (
            .O(N__47422),
            .I(N__47419));
    LocalMux I__11522 (
            .O(N__47419),
            .I(\c0.n18086 ));
    InMux I__11521 (
            .O(N__47416),
            .I(N__47412));
    InMux I__11520 (
            .O(N__47415),
            .I(N__47406));
    LocalMux I__11519 (
            .O(N__47412),
            .I(N__47403));
    InMux I__11518 (
            .O(N__47411),
            .I(N__47398));
    InMux I__11517 (
            .O(N__47410),
            .I(N__47398));
    InMux I__11516 (
            .O(N__47409),
            .I(N__47395));
    LocalMux I__11515 (
            .O(N__47406),
            .I(N__47392));
    Span4Mux_v I__11514 (
            .O(N__47403),
            .I(N__47389));
    LocalMux I__11513 (
            .O(N__47398),
            .I(N__47386));
    LocalMux I__11512 (
            .O(N__47395),
            .I(data_out_frame2_10_1));
    Odrv4 I__11511 (
            .O(N__47392),
            .I(data_out_frame2_10_1));
    Odrv4 I__11510 (
            .O(N__47389),
            .I(data_out_frame2_10_1));
    Odrv4 I__11509 (
            .O(N__47386),
            .I(data_out_frame2_10_1));
    InMux I__11508 (
            .O(N__47377),
            .I(N__47373));
    InMux I__11507 (
            .O(N__47376),
            .I(N__47368));
    LocalMux I__11506 (
            .O(N__47373),
            .I(N__47365));
    InMux I__11505 (
            .O(N__47372),
            .I(N__47362));
    InMux I__11504 (
            .O(N__47371),
            .I(N__47357));
    LocalMux I__11503 (
            .O(N__47368),
            .I(N__47354));
    Span4Mux_v I__11502 (
            .O(N__47365),
            .I(N__47351));
    LocalMux I__11501 (
            .O(N__47362),
            .I(N__47348));
    InMux I__11500 (
            .O(N__47361),
            .I(N__47345));
    InMux I__11499 (
            .O(N__47360),
            .I(N__47342));
    LocalMux I__11498 (
            .O(N__47357),
            .I(N__47339));
    Span4Mux_v I__11497 (
            .O(N__47354),
            .I(N__47332));
    Span4Mux_h I__11496 (
            .O(N__47351),
            .I(N__47332));
    Span4Mux_v I__11495 (
            .O(N__47348),
            .I(N__47332));
    LocalMux I__11494 (
            .O(N__47345),
            .I(N__47329));
    LocalMux I__11493 (
            .O(N__47342),
            .I(data_out_frame2_12_0));
    Odrv4 I__11492 (
            .O(N__47339),
            .I(data_out_frame2_12_0));
    Odrv4 I__11491 (
            .O(N__47332),
            .I(data_out_frame2_12_0));
    Odrv12 I__11490 (
            .O(N__47329),
            .I(data_out_frame2_12_0));
    CascadeMux I__11489 (
            .O(N__47320),
            .I(N__47317));
    InMux I__11488 (
            .O(N__47317),
            .I(N__47314));
    LocalMux I__11487 (
            .O(N__47314),
            .I(N__47309));
    InMux I__11486 (
            .O(N__47313),
            .I(N__47306));
    CascadeMux I__11485 (
            .O(N__47312),
            .I(N__47303));
    Span4Mux_h I__11484 (
            .O(N__47309),
            .I(N__47296));
    LocalMux I__11483 (
            .O(N__47306),
            .I(N__47296));
    InMux I__11482 (
            .O(N__47303),
            .I(N__47293));
    CascadeMux I__11481 (
            .O(N__47302),
            .I(N__47290));
    InMux I__11480 (
            .O(N__47301),
            .I(N__47287));
    Span4Mux_v I__11479 (
            .O(N__47296),
            .I(N__47282));
    LocalMux I__11478 (
            .O(N__47293),
            .I(N__47282));
    InMux I__11477 (
            .O(N__47290),
            .I(N__47279));
    LocalMux I__11476 (
            .O(N__47287),
            .I(N__47276));
    Span4Mux_h I__11475 (
            .O(N__47282),
            .I(N__47271));
    LocalMux I__11474 (
            .O(N__47279),
            .I(N__47271));
    Span4Mux_h I__11473 (
            .O(N__47276),
            .I(N__47267));
    Span4Mux_v I__11472 (
            .O(N__47271),
            .I(N__47264));
    InMux I__11471 (
            .O(N__47270),
            .I(N__47261));
    Span4Mux_h I__11470 (
            .O(N__47267),
            .I(N__47258));
    Span4Mux_h I__11469 (
            .O(N__47264),
            .I(N__47255));
    LocalMux I__11468 (
            .O(N__47261),
            .I(data_out_frame2_8_1));
    Odrv4 I__11467 (
            .O(N__47258),
            .I(data_out_frame2_8_1));
    Odrv4 I__11466 (
            .O(N__47255),
            .I(data_out_frame2_8_1));
    CascadeMux I__11465 (
            .O(N__47248),
            .I(N__47244));
    InMux I__11464 (
            .O(N__47247),
            .I(N__47241));
    InMux I__11463 (
            .O(N__47244),
            .I(N__47238));
    LocalMux I__11462 (
            .O(N__47241),
            .I(N__47232));
    LocalMux I__11461 (
            .O(N__47238),
            .I(N__47232));
    InMux I__11460 (
            .O(N__47237),
            .I(N__47228));
    Span4Mux_h I__11459 (
            .O(N__47232),
            .I(N__47225));
    InMux I__11458 (
            .O(N__47231),
            .I(N__47221));
    LocalMux I__11457 (
            .O(N__47228),
            .I(N__47216));
    Span4Mux_h I__11456 (
            .O(N__47225),
            .I(N__47216));
    InMux I__11455 (
            .O(N__47224),
            .I(N__47213));
    LocalMux I__11454 (
            .O(N__47221),
            .I(N__47210));
    Odrv4 I__11453 (
            .O(N__47216),
            .I(data_out_frame2_14_3));
    LocalMux I__11452 (
            .O(N__47213),
            .I(data_out_frame2_14_3));
    Odrv4 I__11451 (
            .O(N__47210),
            .I(data_out_frame2_14_3));
    CascadeMux I__11450 (
            .O(N__47203),
            .I(\c0.n9895_cascade_ ));
    InMux I__11449 (
            .O(N__47200),
            .I(N__47195));
    InMux I__11448 (
            .O(N__47199),
            .I(N__47192));
    InMux I__11447 (
            .O(N__47198),
            .I(N__47189));
    LocalMux I__11446 (
            .O(N__47195),
            .I(N__47185));
    LocalMux I__11445 (
            .O(N__47192),
            .I(N__47182));
    LocalMux I__11444 (
            .O(N__47189),
            .I(N__47178));
    InMux I__11443 (
            .O(N__47188),
            .I(N__47175));
    Span4Mux_h I__11442 (
            .O(N__47185),
            .I(N__47172));
    Span12Mux_h I__11441 (
            .O(N__47182),
            .I(N__47169));
    InMux I__11440 (
            .O(N__47181),
            .I(N__47166));
    Span12Mux_s9_v I__11439 (
            .O(N__47178),
            .I(N__47163));
    LocalMux I__11438 (
            .O(N__47175),
            .I(data_out_frame2_15_1));
    Odrv4 I__11437 (
            .O(N__47172),
            .I(data_out_frame2_15_1));
    Odrv12 I__11436 (
            .O(N__47169),
            .I(data_out_frame2_15_1));
    LocalMux I__11435 (
            .O(N__47166),
            .I(data_out_frame2_15_1));
    Odrv12 I__11434 (
            .O(N__47163),
            .I(data_out_frame2_15_1));
    CascadeMux I__11433 (
            .O(N__47152),
            .I(N__47149));
    InMux I__11432 (
            .O(N__47149),
            .I(N__47146));
    LocalMux I__11431 (
            .O(N__47146),
            .I(N__47143));
    Odrv4 I__11430 (
            .O(N__47143),
            .I(\c0.n6_adj_2274 ));
    InMux I__11429 (
            .O(N__47140),
            .I(N__47135));
    InMux I__11428 (
            .O(N__47139),
            .I(N__47132));
    InMux I__11427 (
            .O(N__47138),
            .I(N__47129));
    LocalMux I__11426 (
            .O(N__47135),
            .I(N__47126));
    LocalMux I__11425 (
            .O(N__47132),
            .I(N__47123));
    LocalMux I__11424 (
            .O(N__47129),
            .I(N__47120));
    Span4Mux_v I__11423 (
            .O(N__47126),
            .I(N__47117));
    Span4Mux_v I__11422 (
            .O(N__47123),
            .I(N__47112));
    Span4Mux_h I__11421 (
            .O(N__47120),
            .I(N__47112));
    Span4Mux_h I__11420 (
            .O(N__47117),
            .I(N__47109));
    Span4Mux_h I__11419 (
            .O(N__47112),
            .I(N__47106));
    Odrv4 I__11418 (
            .O(N__47109),
            .I(\c0.data_out_9_4 ));
    Odrv4 I__11417 (
            .O(N__47106),
            .I(\c0.data_out_9_4 ));
    CascadeMux I__11416 (
            .O(N__47101),
            .I(N__47098));
    InMux I__11415 (
            .O(N__47098),
            .I(N__47093));
    InMux I__11414 (
            .O(N__47097),
            .I(N__47090));
    InMux I__11413 (
            .O(N__47096),
            .I(N__47087));
    LocalMux I__11412 (
            .O(N__47093),
            .I(N__47084));
    LocalMux I__11411 (
            .O(N__47090),
            .I(N__47081));
    LocalMux I__11410 (
            .O(N__47087),
            .I(N__47078));
    Span4Mux_h I__11409 (
            .O(N__47084),
            .I(N__47075));
    Span4Mux_v I__11408 (
            .O(N__47081),
            .I(N__47072));
    Span4Mux_v I__11407 (
            .O(N__47078),
            .I(N__47069));
    Span4Mux_v I__11406 (
            .O(N__47075),
            .I(N__47064));
    Span4Mux_h I__11405 (
            .O(N__47072),
            .I(N__47064));
    Span4Mux_h I__11404 (
            .O(N__47069),
            .I(N__47061));
    Odrv4 I__11403 (
            .O(N__47064),
            .I(\c0.data_out_10_4 ));
    Odrv4 I__11402 (
            .O(N__47061),
            .I(\c0.data_out_10_4 ));
    InMux I__11401 (
            .O(N__47056),
            .I(N__47053));
    LocalMux I__11400 (
            .O(N__47053),
            .I(N__47050));
    Span4Mux_h I__11399 (
            .O(N__47050),
            .I(N__47046));
    CascadeMux I__11398 (
            .O(N__47049),
            .I(N__47042));
    Span4Mux_h I__11397 (
            .O(N__47046),
            .I(N__47039));
    InMux I__11396 (
            .O(N__47045),
            .I(N__47034));
    InMux I__11395 (
            .O(N__47042),
            .I(N__47034));
    Odrv4 I__11394 (
            .O(N__47039),
            .I(\c0.data_out_7_2 ));
    LocalMux I__11393 (
            .O(N__47034),
            .I(\c0.data_out_7_2 ));
    InMux I__11392 (
            .O(N__47029),
            .I(N__47026));
    LocalMux I__11391 (
            .O(N__47026),
            .I(\c0.n17058 ));
    InMux I__11390 (
            .O(N__47023),
            .I(N__47019));
    InMux I__11389 (
            .O(N__47022),
            .I(N__47016));
    LocalMux I__11388 (
            .O(N__47019),
            .I(\c0.n17028 ));
    LocalMux I__11387 (
            .O(N__47016),
            .I(\c0.n17028 ));
    CascadeMux I__11386 (
            .O(N__47011),
            .I(\c0.n17058_cascade_ ));
    InMux I__11385 (
            .O(N__47008),
            .I(N__47005));
    LocalMux I__11384 (
            .O(N__47005),
            .I(N__47001));
    InMux I__11383 (
            .O(N__47004),
            .I(N__46998));
    Odrv4 I__11382 (
            .O(N__47001),
            .I(\c0.n17094 ));
    LocalMux I__11381 (
            .O(N__46998),
            .I(\c0.n17094 ));
    InMux I__11380 (
            .O(N__46993),
            .I(N__46990));
    LocalMux I__11379 (
            .O(N__46990),
            .I(N__46987));
    Odrv4 I__11378 (
            .O(N__46987),
            .I(\c0.n19_adj_2283 ));
    CascadeMux I__11377 (
            .O(N__46984),
            .I(\c0.n21_adj_2284_cascade_ ));
    InMux I__11376 (
            .O(N__46981),
            .I(N__46978));
    LocalMux I__11375 (
            .O(N__46978),
            .I(N__46975));
    Span4Mux_h I__11374 (
            .O(N__46975),
            .I(N__46972));
    Odrv4 I__11373 (
            .O(N__46972),
            .I(\c0.n20_adj_2282 ));
    InMux I__11372 (
            .O(N__46969),
            .I(N__46963));
    InMux I__11371 (
            .O(N__46968),
            .I(N__46960));
    InMux I__11370 (
            .O(N__46967),
            .I(N__46955));
    InMux I__11369 (
            .O(N__46966),
            .I(N__46955));
    LocalMux I__11368 (
            .O(N__46963),
            .I(N__46952));
    LocalMux I__11367 (
            .O(N__46960),
            .I(N__46949));
    LocalMux I__11366 (
            .O(N__46955),
            .I(N__46946));
    Span4Mux_s3_v I__11365 (
            .O(N__46952),
            .I(N__46943));
    Span4Mux_h I__11364 (
            .O(N__46949),
            .I(N__46940));
    Span4Mux_h I__11363 (
            .O(N__46946),
            .I(N__46937));
    Span4Mux_h I__11362 (
            .O(N__46943),
            .I(N__46934));
    Odrv4 I__11361 (
            .O(N__46940),
            .I(\c0.data_out_9_7 ));
    Odrv4 I__11360 (
            .O(N__46937),
            .I(\c0.data_out_9_7 ));
    Odrv4 I__11359 (
            .O(N__46934),
            .I(\c0.data_out_9_7 ));
    InMux I__11358 (
            .O(N__46927),
            .I(N__46921));
    InMux I__11357 (
            .O(N__46926),
            .I(N__46921));
    LocalMux I__11356 (
            .O(N__46921),
            .I(N__46918));
    Span4Mux_h I__11355 (
            .O(N__46918),
            .I(N__46915));
    Odrv4 I__11354 (
            .O(N__46915),
            .I(\c0.n17007 ));
    InMux I__11353 (
            .O(N__46912),
            .I(N__46908));
    InMux I__11352 (
            .O(N__46911),
            .I(N__46905));
    LocalMux I__11351 (
            .O(N__46908),
            .I(N__46902));
    LocalMux I__11350 (
            .O(N__46905),
            .I(N__46899));
    Span4Mux_h I__11349 (
            .O(N__46902),
            .I(N__46895));
    Span4Mux_h I__11348 (
            .O(N__46899),
            .I(N__46892));
    InMux I__11347 (
            .O(N__46898),
            .I(N__46889));
    Odrv4 I__11346 (
            .O(N__46895),
            .I(\c0.n9505 ));
    Odrv4 I__11345 (
            .O(N__46892),
            .I(\c0.n9505 ));
    LocalMux I__11344 (
            .O(N__46889),
            .I(\c0.n9505 ));
    CascadeMux I__11343 (
            .O(N__46882),
            .I(N__46879));
    InMux I__11342 (
            .O(N__46879),
            .I(N__46875));
    InMux I__11341 (
            .O(N__46878),
            .I(N__46872));
    LocalMux I__11340 (
            .O(N__46875),
            .I(\c0.n17076 ));
    LocalMux I__11339 (
            .O(N__46872),
            .I(\c0.n17076 ));
    InMux I__11338 (
            .O(N__46867),
            .I(N__46864));
    LocalMux I__11337 (
            .O(N__46864),
            .I(N__46860));
    InMux I__11336 (
            .O(N__46863),
            .I(N__46857));
    Span4Mux_h I__11335 (
            .O(N__46860),
            .I(N__46848));
    LocalMux I__11334 (
            .O(N__46857),
            .I(N__46848));
    InMux I__11333 (
            .O(N__46856),
            .I(N__46845));
    InMux I__11332 (
            .O(N__46855),
            .I(N__46842));
    InMux I__11331 (
            .O(N__46854),
            .I(N__46839));
    InMux I__11330 (
            .O(N__46853),
            .I(N__46836));
    Span4Mux_h I__11329 (
            .O(N__46848),
            .I(N__46831));
    LocalMux I__11328 (
            .O(N__46845),
            .I(N__46831));
    LocalMux I__11327 (
            .O(N__46842),
            .I(data_out_8_0));
    LocalMux I__11326 (
            .O(N__46839),
            .I(data_out_8_0));
    LocalMux I__11325 (
            .O(N__46836),
            .I(data_out_8_0));
    Odrv4 I__11324 (
            .O(N__46831),
            .I(data_out_8_0));
    InMux I__11323 (
            .O(N__46822),
            .I(N__46817));
    InMux I__11322 (
            .O(N__46821),
            .I(N__46812));
    InMux I__11321 (
            .O(N__46820),
            .I(N__46812));
    LocalMux I__11320 (
            .O(N__46817),
            .I(N__46809));
    LocalMux I__11319 (
            .O(N__46812),
            .I(\c0.data_out_10_3 ));
    Odrv12 I__11318 (
            .O(N__46809),
            .I(\c0.data_out_10_3 ));
    InMux I__11317 (
            .O(N__46804),
            .I(N__46800));
    InMux I__11316 (
            .O(N__46803),
            .I(N__46795));
    LocalMux I__11315 (
            .O(N__46800),
            .I(N__46792));
    InMux I__11314 (
            .O(N__46799),
            .I(N__46788));
    InMux I__11313 (
            .O(N__46798),
            .I(N__46785));
    LocalMux I__11312 (
            .O(N__46795),
            .I(N__46780));
    Span4Mux_v I__11311 (
            .O(N__46792),
            .I(N__46780));
    InMux I__11310 (
            .O(N__46791),
            .I(N__46777));
    LocalMux I__11309 (
            .O(N__46788),
            .I(N__46772));
    LocalMux I__11308 (
            .O(N__46785),
            .I(N__46772));
    Span4Mux_h I__11307 (
            .O(N__46780),
            .I(N__46769));
    LocalMux I__11306 (
            .O(N__46777),
            .I(N__46766));
    Span4Mux_h I__11305 (
            .O(N__46772),
            .I(N__46763));
    Odrv4 I__11304 (
            .O(N__46769),
            .I(\c0.data_out_9_6 ));
    Odrv4 I__11303 (
            .O(N__46766),
            .I(\c0.data_out_9_6 ));
    Odrv4 I__11302 (
            .O(N__46763),
            .I(\c0.data_out_9_6 ));
    InMux I__11301 (
            .O(N__46756),
            .I(N__46752));
    InMux I__11300 (
            .O(N__46755),
            .I(N__46749));
    LocalMux I__11299 (
            .O(N__46752),
            .I(N__46746));
    LocalMux I__11298 (
            .O(N__46749),
            .I(N__46743));
    Span4Mux_s2_v I__11297 (
            .O(N__46746),
            .I(N__46740));
    Span4Mux_h I__11296 (
            .O(N__46743),
            .I(N__46734));
    Span4Mux_h I__11295 (
            .O(N__46740),
            .I(N__46734));
    InMux I__11294 (
            .O(N__46739),
            .I(N__46731));
    Odrv4 I__11293 (
            .O(N__46734),
            .I(\c0.data_out_10_2 ));
    LocalMux I__11292 (
            .O(N__46731),
            .I(\c0.data_out_10_2 ));
    CascadeMux I__11291 (
            .O(N__46726),
            .I(N__46723));
    InMux I__11290 (
            .O(N__46723),
            .I(N__46720));
    LocalMux I__11289 (
            .O(N__46720),
            .I(N__46716));
    InMux I__11288 (
            .O(N__46719),
            .I(N__46713));
    Span4Mux_h I__11287 (
            .O(N__46716),
            .I(N__46710));
    LocalMux I__11286 (
            .O(N__46713),
            .I(N__46707));
    Odrv4 I__11285 (
            .O(N__46710),
            .I(\c0.n16998 ));
    Odrv4 I__11284 (
            .O(N__46707),
            .I(\c0.n16998 ));
    CascadeMux I__11283 (
            .O(N__46702),
            .I(N__46698));
    InMux I__11282 (
            .O(N__46701),
            .I(N__46694));
    InMux I__11281 (
            .O(N__46698),
            .I(N__46691));
    InMux I__11280 (
            .O(N__46697),
            .I(N__46686));
    LocalMux I__11279 (
            .O(N__46694),
            .I(N__46683));
    LocalMux I__11278 (
            .O(N__46691),
            .I(N__46680));
    InMux I__11277 (
            .O(N__46690),
            .I(N__46677));
    InMux I__11276 (
            .O(N__46689),
            .I(N__46674));
    LocalMux I__11275 (
            .O(N__46686),
            .I(N__46671));
    Span4Mux_v I__11274 (
            .O(N__46683),
            .I(N__46664));
    Span4Mux_v I__11273 (
            .O(N__46680),
            .I(N__46664));
    LocalMux I__11272 (
            .O(N__46677),
            .I(N__46664));
    LocalMux I__11271 (
            .O(N__46674),
            .I(N__46661));
    Odrv4 I__11270 (
            .O(N__46671),
            .I(\c0.data_out_6_2 ));
    Odrv4 I__11269 (
            .O(N__46664),
            .I(\c0.data_out_6_2 ));
    Odrv4 I__11268 (
            .O(N__46661),
            .I(\c0.data_out_6_2 ));
    InMux I__11267 (
            .O(N__46654),
            .I(N__46651));
    LocalMux I__11266 (
            .O(N__46651),
            .I(N__46648));
    Span4Mux_v I__11265 (
            .O(N__46648),
            .I(N__46643));
    InMux I__11264 (
            .O(N__46647),
            .I(N__46640));
    InMux I__11263 (
            .O(N__46646),
            .I(N__46637));
    Span4Mux_h I__11262 (
            .O(N__46643),
            .I(N__46630));
    LocalMux I__11261 (
            .O(N__46640),
            .I(N__46630));
    LocalMux I__11260 (
            .O(N__46637),
            .I(N__46630));
    Span4Mux_v I__11259 (
            .O(N__46630),
            .I(N__46627));
    Odrv4 I__11258 (
            .O(N__46627),
            .I(\c0.data_out_10_6 ));
    CEMux I__11257 (
            .O(N__46624),
            .I(N__46617));
    CEMux I__11256 (
            .O(N__46623),
            .I(N__46613));
    CEMux I__11255 (
            .O(N__46622),
            .I(N__46610));
    CEMux I__11254 (
            .O(N__46621),
            .I(N__46607));
    CEMux I__11253 (
            .O(N__46620),
            .I(N__46603));
    LocalMux I__11252 (
            .O(N__46617),
            .I(N__46600));
    CEMux I__11251 (
            .O(N__46616),
            .I(N__46597));
    LocalMux I__11250 (
            .O(N__46613),
            .I(N__46590));
    LocalMux I__11249 (
            .O(N__46610),
            .I(N__46590));
    LocalMux I__11248 (
            .O(N__46607),
            .I(N__46590));
    CEMux I__11247 (
            .O(N__46606),
            .I(N__46586));
    LocalMux I__11246 (
            .O(N__46603),
            .I(N__46583));
    Span4Mux_v I__11245 (
            .O(N__46600),
            .I(N__46580));
    LocalMux I__11244 (
            .O(N__46597),
            .I(N__46577));
    Span4Mux_v I__11243 (
            .O(N__46590),
            .I(N__46574));
    CEMux I__11242 (
            .O(N__46589),
            .I(N__46571));
    LocalMux I__11241 (
            .O(N__46586),
            .I(N__46568));
    Span4Mux_h I__11240 (
            .O(N__46583),
            .I(N__46564));
    Span4Mux_h I__11239 (
            .O(N__46580),
            .I(N__46555));
    Span4Mux_h I__11238 (
            .O(N__46577),
            .I(N__46555));
    Span4Mux_h I__11237 (
            .O(N__46574),
            .I(N__46555));
    LocalMux I__11236 (
            .O(N__46571),
            .I(N__46555));
    IoSpan4Mux I__11235 (
            .O(N__46568),
            .I(N__46552));
    InMux I__11234 (
            .O(N__46567),
            .I(N__46549));
    Span4Mux_h I__11233 (
            .O(N__46564),
            .I(N__46546));
    Span4Mux_h I__11232 (
            .O(N__46555),
            .I(N__46543));
    IoSpan4Mux I__11231 (
            .O(N__46552),
            .I(N__46540));
    LocalMux I__11230 (
            .O(N__46549),
            .I(N__46537));
    Span4Mux_h I__11229 (
            .O(N__46546),
            .I(N__46534));
    Span4Mux_v I__11228 (
            .O(N__46543),
            .I(N__46531));
    IoSpan4Mux I__11227 (
            .O(N__46540),
            .I(N__46526));
    Span4Mux_h I__11226 (
            .O(N__46537),
            .I(N__46526));
    Odrv4 I__11225 (
            .O(N__46534),
            .I(data_out_10__7__N_110));
    Odrv4 I__11224 (
            .O(N__46531),
            .I(data_out_10__7__N_110));
    Odrv4 I__11223 (
            .O(N__46526),
            .I(data_out_10__7__N_110));
    InMux I__11222 (
            .O(N__46519),
            .I(N__46515));
    CascadeMux I__11221 (
            .O(N__46518),
            .I(N__46512));
    LocalMux I__11220 (
            .O(N__46515),
            .I(N__46509));
    InMux I__11219 (
            .O(N__46512),
            .I(N__46506));
    Odrv12 I__11218 (
            .O(N__46509),
            .I(rand_setpoint_21));
    LocalMux I__11217 (
            .O(N__46506),
            .I(rand_setpoint_21));
    CascadeMux I__11216 (
            .O(N__46501),
            .I(N__46498));
    InMux I__11215 (
            .O(N__46498),
            .I(N__46495));
    LocalMux I__11214 (
            .O(N__46495),
            .I(\c0.n17522 ));
    InMux I__11213 (
            .O(N__46492),
            .I(N__46482));
    InMux I__11212 (
            .O(N__46491),
            .I(N__46476));
    InMux I__11211 (
            .O(N__46490),
            .I(N__46472));
    InMux I__11210 (
            .O(N__46489),
            .I(N__46467));
    InMux I__11209 (
            .O(N__46488),
            .I(N__46467));
    InMux I__11208 (
            .O(N__46487),
            .I(N__46459));
    InMux I__11207 (
            .O(N__46486),
            .I(N__46459));
    InMux I__11206 (
            .O(N__46485),
            .I(N__46459));
    LocalMux I__11205 (
            .O(N__46482),
            .I(N__46456));
    InMux I__11204 (
            .O(N__46481),
            .I(N__46453));
    InMux I__11203 (
            .O(N__46480),
            .I(N__46450));
    InMux I__11202 (
            .O(N__46479),
            .I(N__46444));
    LocalMux I__11201 (
            .O(N__46476),
            .I(N__46441));
    InMux I__11200 (
            .O(N__46475),
            .I(N__46438));
    LocalMux I__11199 (
            .O(N__46472),
            .I(N__46427));
    LocalMux I__11198 (
            .O(N__46467),
            .I(N__46427));
    InMux I__11197 (
            .O(N__46466),
            .I(N__46424));
    LocalMux I__11196 (
            .O(N__46459),
            .I(N__46408));
    Span4Mux_v I__11195 (
            .O(N__46456),
            .I(N__46408));
    LocalMux I__11194 (
            .O(N__46453),
            .I(N__46408));
    LocalMux I__11193 (
            .O(N__46450),
            .I(N__46405));
    InMux I__11192 (
            .O(N__46449),
            .I(N__46396));
    InMux I__11191 (
            .O(N__46448),
            .I(N__46390));
    InMux I__11190 (
            .O(N__46447),
            .I(N__46390));
    LocalMux I__11189 (
            .O(N__46444),
            .I(N__46383));
    Span4Mux_v I__11188 (
            .O(N__46441),
            .I(N__46383));
    LocalMux I__11187 (
            .O(N__46438),
            .I(N__46383));
    InMux I__11186 (
            .O(N__46437),
            .I(N__46380));
    InMux I__11185 (
            .O(N__46436),
            .I(N__46369));
    InMux I__11184 (
            .O(N__46435),
            .I(N__46369));
    InMux I__11183 (
            .O(N__46434),
            .I(N__46369));
    InMux I__11182 (
            .O(N__46433),
            .I(N__46369));
    InMux I__11181 (
            .O(N__46432),
            .I(N__46369));
    Span4Mux_v I__11180 (
            .O(N__46427),
            .I(N__46366));
    LocalMux I__11179 (
            .O(N__46424),
            .I(N__46363));
    InMux I__11178 (
            .O(N__46423),
            .I(N__46359));
    InMux I__11177 (
            .O(N__46422),
            .I(N__46356));
    InMux I__11176 (
            .O(N__46421),
            .I(N__46353));
    InMux I__11175 (
            .O(N__46420),
            .I(N__46344));
    InMux I__11174 (
            .O(N__46419),
            .I(N__46344));
    InMux I__11173 (
            .O(N__46418),
            .I(N__46344));
    InMux I__11172 (
            .O(N__46417),
            .I(N__46344));
    InMux I__11171 (
            .O(N__46416),
            .I(N__46339));
    InMux I__11170 (
            .O(N__46415),
            .I(N__46339));
    Span4Mux_v I__11169 (
            .O(N__46408),
            .I(N__46336));
    Span4Mux_v I__11168 (
            .O(N__46405),
            .I(N__46333));
    InMux I__11167 (
            .O(N__46404),
            .I(N__46322));
    InMux I__11166 (
            .O(N__46403),
            .I(N__46322));
    InMux I__11165 (
            .O(N__46402),
            .I(N__46322));
    InMux I__11164 (
            .O(N__46401),
            .I(N__46322));
    InMux I__11163 (
            .O(N__46400),
            .I(N__46322));
    CascadeMux I__11162 (
            .O(N__46399),
            .I(N__46318));
    LocalMux I__11161 (
            .O(N__46396),
            .I(N__46315));
    InMux I__11160 (
            .O(N__46395),
            .I(N__46312));
    LocalMux I__11159 (
            .O(N__46390),
            .I(N__46307));
    Span4Mux_h I__11158 (
            .O(N__46383),
            .I(N__46307));
    LocalMux I__11157 (
            .O(N__46380),
            .I(N__46293));
    LocalMux I__11156 (
            .O(N__46369),
            .I(N__46293));
    Span4Mux_h I__11155 (
            .O(N__46366),
            .I(N__46288));
    Span4Mux_v I__11154 (
            .O(N__46363),
            .I(N__46288));
    InMux I__11153 (
            .O(N__46362),
            .I(N__46285));
    LocalMux I__11152 (
            .O(N__46359),
            .I(N__46268));
    LocalMux I__11151 (
            .O(N__46356),
            .I(N__46268));
    LocalMux I__11150 (
            .O(N__46353),
            .I(N__46268));
    LocalMux I__11149 (
            .O(N__46344),
            .I(N__46268));
    LocalMux I__11148 (
            .O(N__46339),
            .I(N__46268));
    Sp12to4 I__11147 (
            .O(N__46336),
            .I(N__46268));
    Sp12to4 I__11146 (
            .O(N__46333),
            .I(N__46268));
    LocalMux I__11145 (
            .O(N__46322),
            .I(N__46268));
    InMux I__11144 (
            .O(N__46321),
            .I(N__46263));
    InMux I__11143 (
            .O(N__46318),
            .I(N__46263));
    Span4Mux_v I__11142 (
            .O(N__46315),
            .I(N__46256));
    LocalMux I__11141 (
            .O(N__46312),
            .I(N__46256));
    Span4Mux_h I__11140 (
            .O(N__46307),
            .I(N__46256));
    InMux I__11139 (
            .O(N__46306),
            .I(N__46253));
    InMux I__11138 (
            .O(N__46305),
            .I(N__46242));
    InMux I__11137 (
            .O(N__46304),
            .I(N__46242));
    InMux I__11136 (
            .O(N__46303),
            .I(N__46242));
    InMux I__11135 (
            .O(N__46302),
            .I(N__46242));
    InMux I__11134 (
            .O(N__46301),
            .I(N__46242));
    InMux I__11133 (
            .O(N__46300),
            .I(N__46235));
    InMux I__11132 (
            .O(N__46299),
            .I(N__46235));
    InMux I__11131 (
            .O(N__46298),
            .I(N__46235));
    Span4Mux_h I__11130 (
            .O(N__46293),
            .I(N__46232));
    Span4Mux_h I__11129 (
            .O(N__46288),
            .I(N__46227));
    LocalMux I__11128 (
            .O(N__46285),
            .I(N__46227));
    Span12Mux_h I__11127 (
            .O(N__46268),
            .I(N__46224));
    LocalMux I__11126 (
            .O(N__46263),
            .I(N__46221));
    Span4Mux_h I__11125 (
            .O(N__46256),
            .I(N__46218));
    LocalMux I__11124 (
            .O(N__46253),
            .I(UART_TRANSMITTER_state_1));
    LocalMux I__11123 (
            .O(N__46242),
            .I(UART_TRANSMITTER_state_1));
    LocalMux I__11122 (
            .O(N__46235),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__11121 (
            .O(N__46232),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__11120 (
            .O(N__46227),
            .I(UART_TRANSMITTER_state_1));
    Odrv12 I__11119 (
            .O(N__46224),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__11118 (
            .O(N__46221),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__11117 (
            .O(N__46218),
            .I(UART_TRANSMITTER_state_1));
    InMux I__11116 (
            .O(N__46201),
            .I(N__46196));
    InMux I__11115 (
            .O(N__46200),
            .I(N__46193));
    InMux I__11114 (
            .O(N__46199),
            .I(N__46189));
    LocalMux I__11113 (
            .O(N__46196),
            .I(N__46186));
    LocalMux I__11112 (
            .O(N__46193),
            .I(N__46183));
    InMux I__11111 (
            .O(N__46192),
            .I(N__46180));
    LocalMux I__11110 (
            .O(N__46189),
            .I(N__46177));
    Span4Mux_v I__11109 (
            .O(N__46186),
            .I(N__46174));
    Span4Mux_v I__11108 (
            .O(N__46183),
            .I(N__46171));
    LocalMux I__11107 (
            .O(N__46180),
            .I(N__46166));
    Span4Mux_v I__11106 (
            .O(N__46177),
            .I(N__46166));
    Span4Mux_v I__11105 (
            .O(N__46174),
            .I(N__46163));
    Span4Mux_s1_v I__11104 (
            .O(N__46171),
            .I(N__46160));
    Span4Mux_v I__11103 (
            .O(N__46166),
            .I(N__46155));
    Span4Mux_h I__11102 (
            .O(N__46163),
            .I(N__46155));
    Odrv4 I__11101 (
            .O(N__46160),
            .I(\c0.data_out_6_5 ));
    Odrv4 I__11100 (
            .O(N__46155),
            .I(\c0.data_out_6_5 ));
    CascadeMux I__11099 (
            .O(N__46150),
            .I(N__46146));
    CascadeMux I__11098 (
            .O(N__46149),
            .I(N__46143));
    InMux I__11097 (
            .O(N__46146),
            .I(N__46140));
    InMux I__11096 (
            .O(N__46143),
            .I(N__46134));
    LocalMux I__11095 (
            .O(N__46140),
            .I(N__46125));
    InMux I__11094 (
            .O(N__46139),
            .I(N__46122));
    CascadeMux I__11093 (
            .O(N__46138),
            .I(N__46119));
    CEMux I__11092 (
            .O(N__46137),
            .I(N__46116));
    LocalMux I__11091 (
            .O(N__46134),
            .I(N__46113));
    CascadeMux I__11090 (
            .O(N__46133),
            .I(N__46110));
    CascadeMux I__11089 (
            .O(N__46132),
            .I(N__46107));
    CEMux I__11088 (
            .O(N__46131),
            .I(N__46103));
    CEMux I__11087 (
            .O(N__46130),
            .I(N__46100));
    CEMux I__11086 (
            .O(N__46129),
            .I(N__46097));
    CEMux I__11085 (
            .O(N__46128),
            .I(N__46094));
    Span4Mux_h I__11084 (
            .O(N__46125),
            .I(N__46089));
    LocalMux I__11083 (
            .O(N__46122),
            .I(N__46089));
    InMux I__11082 (
            .O(N__46119),
            .I(N__46086));
    LocalMux I__11081 (
            .O(N__46116),
            .I(N__46083));
    Span4Mux_h I__11080 (
            .O(N__46113),
            .I(N__46080));
    InMux I__11079 (
            .O(N__46110),
            .I(N__46077));
    InMux I__11078 (
            .O(N__46107),
            .I(N__46074));
    CEMux I__11077 (
            .O(N__46106),
            .I(N__46071));
    LocalMux I__11076 (
            .O(N__46103),
            .I(N__46066));
    LocalMux I__11075 (
            .O(N__46100),
            .I(N__46066));
    LocalMux I__11074 (
            .O(N__46097),
            .I(N__46063));
    LocalMux I__11073 (
            .O(N__46094),
            .I(N__46058));
    Span4Mux_h I__11072 (
            .O(N__46089),
            .I(N__46058));
    LocalMux I__11071 (
            .O(N__46086),
            .I(N__46051));
    Span4Mux_s2_v I__11070 (
            .O(N__46083),
            .I(N__46051));
    Span4Mux_h I__11069 (
            .O(N__46080),
            .I(N__46051));
    LocalMux I__11068 (
            .O(N__46077),
            .I(N__46048));
    LocalMux I__11067 (
            .O(N__46074),
            .I(N__46041));
    LocalMux I__11066 (
            .O(N__46071),
            .I(N__46041));
    Span4Mux_h I__11065 (
            .O(N__46066),
            .I(N__46041));
    Span4Mux_h I__11064 (
            .O(N__46063),
            .I(N__46036));
    Span4Mux_h I__11063 (
            .O(N__46058),
            .I(N__46036));
    Span4Mux_h I__11062 (
            .O(N__46051),
            .I(N__46033));
    Odrv12 I__11061 (
            .O(N__46048),
            .I(n10055));
    Odrv4 I__11060 (
            .O(N__46041),
            .I(n10055));
    Odrv4 I__11059 (
            .O(N__46036),
            .I(n10055));
    Odrv4 I__11058 (
            .O(N__46033),
            .I(n10055));
    InMux I__11057 (
            .O(N__46024),
            .I(N__46021));
    LocalMux I__11056 (
            .O(N__46021),
            .I(N__46018));
    Span4Mux_s1_v I__11055 (
            .O(N__46018),
            .I(N__46014));
    CascadeMux I__11054 (
            .O(N__46017),
            .I(N__46011));
    Span4Mux_h I__11053 (
            .O(N__46014),
            .I(N__46008));
    InMux I__11052 (
            .O(N__46011),
            .I(N__46005));
    Odrv4 I__11051 (
            .O(N__46008),
            .I(rand_setpoint_10));
    LocalMux I__11050 (
            .O(N__46005),
            .I(rand_setpoint_10));
    CascadeMux I__11049 (
            .O(N__46000),
            .I(N__45983));
    CascadeMux I__11048 (
            .O(N__45999),
            .I(N__45979));
    InMux I__11047 (
            .O(N__45998),
            .I(N__45971));
    InMux I__11046 (
            .O(N__45997),
            .I(N__45971));
    InMux I__11045 (
            .O(N__45996),
            .I(N__45968));
    InMux I__11044 (
            .O(N__45995),
            .I(N__45957));
    InMux I__11043 (
            .O(N__45994),
            .I(N__45957));
    InMux I__11042 (
            .O(N__45993),
            .I(N__45957));
    InMux I__11041 (
            .O(N__45992),
            .I(N__45957));
    InMux I__11040 (
            .O(N__45991),
            .I(N__45957));
    CascadeMux I__11039 (
            .O(N__45990),
            .I(N__45948));
    CascadeMux I__11038 (
            .O(N__45989),
            .I(N__45944));
    CascadeMux I__11037 (
            .O(N__45988),
            .I(N__45940));
    CascadeMux I__11036 (
            .O(N__45987),
            .I(N__45937));
    InMux I__11035 (
            .O(N__45986),
            .I(N__45932));
    InMux I__11034 (
            .O(N__45983),
            .I(N__45925));
    CascadeMux I__11033 (
            .O(N__45982),
            .I(N__45921));
    InMux I__11032 (
            .O(N__45979),
            .I(N__45915));
    InMux I__11031 (
            .O(N__45978),
            .I(N__45915));
    InMux I__11030 (
            .O(N__45977),
            .I(N__45912));
    CascadeMux I__11029 (
            .O(N__45976),
            .I(N__45908));
    LocalMux I__11028 (
            .O(N__45971),
            .I(N__45898));
    LocalMux I__11027 (
            .O(N__45968),
            .I(N__45898));
    LocalMux I__11026 (
            .O(N__45957),
            .I(N__45898));
    InMux I__11025 (
            .O(N__45956),
            .I(N__45889));
    InMux I__11024 (
            .O(N__45955),
            .I(N__45889));
    InMux I__11023 (
            .O(N__45954),
            .I(N__45889));
    InMux I__11022 (
            .O(N__45953),
            .I(N__45889));
    CascadeMux I__11021 (
            .O(N__45952),
            .I(N__45886));
    CascadeMux I__11020 (
            .O(N__45951),
            .I(N__45883));
    InMux I__11019 (
            .O(N__45948),
            .I(N__45880));
    InMux I__11018 (
            .O(N__45947),
            .I(N__45876));
    InMux I__11017 (
            .O(N__45944),
            .I(N__45869));
    InMux I__11016 (
            .O(N__45943),
            .I(N__45869));
    InMux I__11015 (
            .O(N__45940),
            .I(N__45864));
    InMux I__11014 (
            .O(N__45937),
            .I(N__45864));
    InMux I__11013 (
            .O(N__45936),
            .I(N__45861));
    InMux I__11012 (
            .O(N__45935),
            .I(N__45858));
    LocalMux I__11011 (
            .O(N__45932),
            .I(N__45855));
    InMux I__11010 (
            .O(N__45931),
            .I(N__45852));
    InMux I__11009 (
            .O(N__45930),
            .I(N__45849));
    CascadeMux I__11008 (
            .O(N__45929),
            .I(N__45845));
    CascadeMux I__11007 (
            .O(N__45928),
            .I(N__45841));
    LocalMux I__11006 (
            .O(N__45925),
            .I(N__45838));
    InMux I__11005 (
            .O(N__45924),
            .I(N__45835));
    InMux I__11004 (
            .O(N__45921),
            .I(N__45830));
    InMux I__11003 (
            .O(N__45920),
            .I(N__45830));
    LocalMux I__11002 (
            .O(N__45915),
            .I(N__45825));
    LocalMux I__11001 (
            .O(N__45912),
            .I(N__45825));
    InMux I__11000 (
            .O(N__45911),
            .I(N__45820));
    InMux I__10999 (
            .O(N__45908),
            .I(N__45820));
    InMux I__10998 (
            .O(N__45907),
            .I(N__45817));
    InMux I__10997 (
            .O(N__45906),
            .I(N__45812));
    InMux I__10996 (
            .O(N__45905),
            .I(N__45812));
    Span4Mux_h I__10995 (
            .O(N__45898),
            .I(N__45807));
    LocalMux I__10994 (
            .O(N__45889),
            .I(N__45807));
    InMux I__10993 (
            .O(N__45886),
            .I(N__45804));
    InMux I__10992 (
            .O(N__45883),
            .I(N__45798));
    LocalMux I__10991 (
            .O(N__45880),
            .I(N__45795));
    InMux I__10990 (
            .O(N__45879),
            .I(N__45792));
    LocalMux I__10989 (
            .O(N__45876),
            .I(N__45789));
    InMux I__10988 (
            .O(N__45875),
            .I(N__45786));
    InMux I__10987 (
            .O(N__45874),
            .I(N__45778));
    LocalMux I__10986 (
            .O(N__45869),
            .I(N__45771));
    LocalMux I__10985 (
            .O(N__45864),
            .I(N__45771));
    LocalMux I__10984 (
            .O(N__45861),
            .I(N__45771));
    LocalMux I__10983 (
            .O(N__45858),
            .I(N__45762));
    Span4Mux_h I__10982 (
            .O(N__45855),
            .I(N__45762));
    LocalMux I__10981 (
            .O(N__45852),
            .I(N__45762));
    LocalMux I__10980 (
            .O(N__45849),
            .I(N__45762));
    CascadeMux I__10979 (
            .O(N__45848),
            .I(N__45757));
    InMux I__10978 (
            .O(N__45845),
            .I(N__45754));
    InMux I__10977 (
            .O(N__45844),
            .I(N__45751));
    InMux I__10976 (
            .O(N__45841),
            .I(N__45748));
    Span4Mux_v I__10975 (
            .O(N__45838),
            .I(N__45745));
    LocalMux I__10974 (
            .O(N__45835),
            .I(N__45742));
    LocalMux I__10973 (
            .O(N__45830),
            .I(N__45739));
    Span4Mux_v I__10972 (
            .O(N__45825),
            .I(N__45734));
    LocalMux I__10971 (
            .O(N__45820),
            .I(N__45734));
    LocalMux I__10970 (
            .O(N__45817),
            .I(N__45725));
    LocalMux I__10969 (
            .O(N__45812),
            .I(N__45725));
    Span4Mux_h I__10968 (
            .O(N__45807),
            .I(N__45725));
    LocalMux I__10967 (
            .O(N__45804),
            .I(N__45725));
    InMux I__10966 (
            .O(N__45803),
            .I(N__45718));
    InMux I__10965 (
            .O(N__45802),
            .I(N__45718));
    InMux I__10964 (
            .O(N__45801),
            .I(N__45718));
    LocalMux I__10963 (
            .O(N__45798),
            .I(N__45713));
    Span4Mux_v I__10962 (
            .O(N__45795),
            .I(N__45713));
    LocalMux I__10961 (
            .O(N__45792),
            .I(N__45706));
    Span4Mux_s1_v I__10960 (
            .O(N__45789),
            .I(N__45706));
    LocalMux I__10959 (
            .O(N__45786),
            .I(N__45706));
    InMux I__10958 (
            .O(N__45785),
            .I(N__45695));
    InMux I__10957 (
            .O(N__45784),
            .I(N__45695));
    InMux I__10956 (
            .O(N__45783),
            .I(N__45695));
    InMux I__10955 (
            .O(N__45782),
            .I(N__45695));
    InMux I__10954 (
            .O(N__45781),
            .I(N__45695));
    LocalMux I__10953 (
            .O(N__45778),
            .I(N__45688));
    Span4Mux_v I__10952 (
            .O(N__45771),
            .I(N__45688));
    Span4Mux_v I__10951 (
            .O(N__45762),
            .I(N__45688));
    InMux I__10950 (
            .O(N__45761),
            .I(N__45683));
    InMux I__10949 (
            .O(N__45760),
            .I(N__45683));
    InMux I__10948 (
            .O(N__45757),
            .I(N__45680));
    LocalMux I__10947 (
            .O(N__45754),
            .I(N__45667));
    LocalMux I__10946 (
            .O(N__45751),
            .I(N__45667));
    LocalMux I__10945 (
            .O(N__45748),
            .I(N__45667));
    Span4Mux_h I__10944 (
            .O(N__45745),
            .I(N__45667));
    Span4Mux_v I__10943 (
            .O(N__45742),
            .I(N__45667));
    Span4Mux_v I__10942 (
            .O(N__45739),
            .I(N__45667));
    Span4Mux_h I__10941 (
            .O(N__45734),
            .I(N__45662));
    Span4Mux_h I__10940 (
            .O(N__45725),
            .I(N__45662));
    LocalMux I__10939 (
            .O(N__45718),
            .I(N__45651));
    Sp12to4 I__10938 (
            .O(N__45713),
            .I(N__45651));
    Sp12to4 I__10937 (
            .O(N__45706),
            .I(N__45651));
    LocalMux I__10936 (
            .O(N__45695),
            .I(N__45651));
    Sp12to4 I__10935 (
            .O(N__45688),
            .I(N__45651));
    LocalMux I__10934 (
            .O(N__45683),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__10933 (
            .O(N__45680),
            .I(UART_TRANSMITTER_state_0));
    Odrv4 I__10932 (
            .O(N__45667),
            .I(UART_TRANSMITTER_state_0));
    Odrv4 I__10931 (
            .O(N__45662),
            .I(UART_TRANSMITTER_state_0));
    Odrv12 I__10930 (
            .O(N__45651),
            .I(UART_TRANSMITTER_state_0));
    CascadeMux I__10929 (
            .O(N__45640),
            .I(N__45637));
    InMux I__10928 (
            .O(N__45637),
            .I(N__45634));
    LocalMux I__10927 (
            .O(N__45634),
            .I(N__45631));
    Odrv12 I__10926 (
            .O(N__45631),
            .I(\c0.n17450 ));
    InMux I__10925 (
            .O(N__45628),
            .I(N__45625));
    LocalMux I__10924 (
            .O(N__45625),
            .I(N__45621));
    CascadeMux I__10923 (
            .O(N__45624),
            .I(N__45618));
    Span4Mux_v I__10922 (
            .O(N__45621),
            .I(N__45613));
    InMux I__10921 (
            .O(N__45618),
            .I(N__45606));
    InMux I__10920 (
            .O(N__45617),
            .I(N__45606));
    InMux I__10919 (
            .O(N__45616),
            .I(N__45606));
    Odrv4 I__10918 (
            .O(N__45613),
            .I(data_out_frame2_7_5));
    LocalMux I__10917 (
            .O(N__45606),
            .I(data_out_frame2_7_5));
    CascadeMux I__10916 (
            .O(N__45601),
            .I(N__45598));
    InMux I__10915 (
            .O(N__45598),
            .I(N__45593));
    InMux I__10914 (
            .O(N__45597),
            .I(N__45590));
    InMux I__10913 (
            .O(N__45596),
            .I(N__45587));
    LocalMux I__10912 (
            .O(N__45593),
            .I(N__45582));
    LocalMux I__10911 (
            .O(N__45590),
            .I(N__45582));
    LocalMux I__10910 (
            .O(N__45587),
            .I(\c0.n9678 ));
    Odrv12 I__10909 (
            .O(N__45582),
            .I(\c0.n9678 ));
    InMux I__10908 (
            .O(N__45577),
            .I(N__45574));
    LocalMux I__10907 (
            .O(N__45574),
            .I(\c0.n18092 ));
    InMux I__10906 (
            .O(N__45571),
            .I(N__45568));
    LocalMux I__10905 (
            .O(N__45568),
            .I(\c0.n22_adj_2352 ));
    InMux I__10904 (
            .O(N__45565),
            .I(N__45562));
    LocalMux I__10903 (
            .O(N__45562),
            .I(N__45559));
    Span4Mux_v I__10902 (
            .O(N__45559),
            .I(N__45556));
    Span4Mux_h I__10901 (
            .O(N__45556),
            .I(N__45553));
    Odrv4 I__10900 (
            .O(N__45553),
            .I(\c0.tx2.r_Tx_Data_7 ));
    SRMux I__10899 (
            .O(N__45550),
            .I(N__45541));
    CascadeMux I__10898 (
            .O(N__45549),
            .I(N__45538));
    InMux I__10897 (
            .O(N__45548),
            .I(N__45533));
    InMux I__10896 (
            .O(N__45547),
            .I(N__45526));
    InMux I__10895 (
            .O(N__45546),
            .I(N__45526));
    InMux I__10894 (
            .O(N__45545),
            .I(N__45526));
    InMux I__10893 (
            .O(N__45544),
            .I(N__45523));
    LocalMux I__10892 (
            .O(N__45541),
            .I(N__45520));
    InMux I__10891 (
            .O(N__45538),
            .I(N__45517));
    CascadeMux I__10890 (
            .O(N__45537),
            .I(N__45511));
    InMux I__10889 (
            .O(N__45536),
            .I(N__45507));
    LocalMux I__10888 (
            .O(N__45533),
            .I(N__45504));
    LocalMux I__10887 (
            .O(N__45526),
            .I(N__45499));
    LocalMux I__10886 (
            .O(N__45523),
            .I(N__45499));
    Span4Mux_s2_v I__10885 (
            .O(N__45520),
            .I(N__45496));
    LocalMux I__10884 (
            .O(N__45517),
            .I(N__45493));
    InMux I__10883 (
            .O(N__45516),
            .I(N__45488));
    InMux I__10882 (
            .O(N__45515),
            .I(N__45483));
    InMux I__10881 (
            .O(N__45514),
            .I(N__45480));
    InMux I__10880 (
            .O(N__45511),
            .I(N__45477));
    InMux I__10879 (
            .O(N__45510),
            .I(N__45474));
    LocalMux I__10878 (
            .O(N__45507),
            .I(N__45471));
    Span4Mux_s2_v I__10877 (
            .O(N__45504),
            .I(N__45462));
    Span4Mux_v I__10876 (
            .O(N__45499),
            .I(N__45462));
    Span4Mux_h I__10875 (
            .O(N__45496),
            .I(N__45462));
    Span4Mux_s2_v I__10874 (
            .O(N__45493),
            .I(N__45462));
    InMux I__10873 (
            .O(N__45492),
            .I(N__45457));
    InMux I__10872 (
            .O(N__45491),
            .I(N__45457));
    LocalMux I__10871 (
            .O(N__45488),
            .I(N__45451));
    InMux I__10870 (
            .O(N__45487),
            .I(N__45446));
    InMux I__10869 (
            .O(N__45486),
            .I(N__45446));
    LocalMux I__10868 (
            .O(N__45483),
            .I(N__45443));
    LocalMux I__10867 (
            .O(N__45480),
            .I(N__45436));
    LocalMux I__10866 (
            .O(N__45477),
            .I(N__45436));
    LocalMux I__10865 (
            .O(N__45474),
            .I(N__45436));
    Span4Mux_s2_v I__10864 (
            .O(N__45471),
            .I(N__45428));
    Span4Mux_h I__10863 (
            .O(N__45462),
            .I(N__45428));
    LocalMux I__10862 (
            .O(N__45457),
            .I(N__45428));
    InMux I__10861 (
            .O(N__45456),
            .I(N__45425));
    InMux I__10860 (
            .O(N__45455),
            .I(N__45422));
    InMux I__10859 (
            .O(N__45454),
            .I(N__45419));
    Span4Mux_v I__10858 (
            .O(N__45451),
            .I(N__45416));
    LocalMux I__10857 (
            .O(N__45446),
            .I(N__45411));
    Span12Mux_s3_v I__10856 (
            .O(N__45443),
            .I(N__45411));
    Span4Mux_v I__10855 (
            .O(N__45436),
            .I(N__45408));
    InMux I__10854 (
            .O(N__45435),
            .I(N__45405));
    Span4Mux_h I__10853 (
            .O(N__45428),
            .I(N__45402));
    LocalMux I__10852 (
            .O(N__45425),
            .I(N__45399));
    LocalMux I__10851 (
            .O(N__45422),
            .I(n4445));
    LocalMux I__10850 (
            .O(N__45419),
            .I(n4445));
    Odrv4 I__10849 (
            .O(N__45416),
            .I(n4445));
    Odrv12 I__10848 (
            .O(N__45411),
            .I(n4445));
    Odrv4 I__10847 (
            .O(N__45408),
            .I(n4445));
    LocalMux I__10846 (
            .O(N__45405),
            .I(n4445));
    Odrv4 I__10845 (
            .O(N__45402),
            .I(n4445));
    Odrv4 I__10844 (
            .O(N__45399),
            .I(n4445));
    CascadeMux I__10843 (
            .O(N__45382),
            .I(N__45379));
    InMux I__10842 (
            .O(N__45379),
            .I(N__45375));
    InMux I__10841 (
            .O(N__45378),
            .I(N__45372));
    LocalMux I__10840 (
            .O(N__45375),
            .I(data_out_0_0));
    LocalMux I__10839 (
            .O(N__45372),
            .I(data_out_0_0));
    InMux I__10838 (
            .O(N__45367),
            .I(N__45364));
    LocalMux I__10837 (
            .O(N__45364),
            .I(N__45358));
    InMux I__10836 (
            .O(N__45363),
            .I(N__45355));
    InMux I__10835 (
            .O(N__45362),
            .I(N__45352));
    CascadeMux I__10834 (
            .O(N__45361),
            .I(N__45349));
    Span4Mux_h I__10833 (
            .O(N__45358),
            .I(N__45343));
    LocalMux I__10832 (
            .O(N__45355),
            .I(N__45343));
    LocalMux I__10831 (
            .O(N__45352),
            .I(N__45340));
    InMux I__10830 (
            .O(N__45349),
            .I(N__45337));
    InMux I__10829 (
            .O(N__45348),
            .I(N__45333));
    Span4Mux_h I__10828 (
            .O(N__45343),
            .I(N__45330));
    Span4Mux_h I__10827 (
            .O(N__45340),
            .I(N__45327));
    LocalMux I__10826 (
            .O(N__45337),
            .I(N__45324));
    InMux I__10825 (
            .O(N__45336),
            .I(N__45321));
    LocalMux I__10824 (
            .O(N__45333),
            .I(N__45318));
    Span4Mux_v I__10823 (
            .O(N__45330),
            .I(N__45315));
    Span4Mux_v I__10822 (
            .O(N__45327),
            .I(N__45310));
    Span4Mux_v I__10821 (
            .O(N__45324),
            .I(N__45310));
    LocalMux I__10820 (
            .O(N__45321),
            .I(data_out_frame2_12_3));
    Odrv4 I__10819 (
            .O(N__45318),
            .I(data_out_frame2_12_3));
    Odrv4 I__10818 (
            .O(N__45315),
            .I(data_out_frame2_12_3));
    Odrv4 I__10817 (
            .O(N__45310),
            .I(data_out_frame2_12_3));
    InMux I__10816 (
            .O(N__45301),
            .I(N__45297));
    InMux I__10815 (
            .O(N__45300),
            .I(N__45294));
    LocalMux I__10814 (
            .O(N__45297),
            .I(N__45289));
    LocalMux I__10813 (
            .O(N__45294),
            .I(N__45286));
    InMux I__10812 (
            .O(N__45293),
            .I(N__45283));
    InMux I__10811 (
            .O(N__45292),
            .I(N__45280));
    Span4Mux_v I__10810 (
            .O(N__45289),
            .I(N__45272));
    Span4Mux_v I__10809 (
            .O(N__45286),
            .I(N__45272));
    LocalMux I__10808 (
            .O(N__45283),
            .I(N__45272));
    LocalMux I__10807 (
            .O(N__45280),
            .I(N__45269));
    InMux I__10806 (
            .O(N__45279),
            .I(N__45266));
    Span4Mux_h I__10805 (
            .O(N__45272),
            .I(N__45261));
    Span4Mux_s2_v I__10804 (
            .O(N__45269),
            .I(N__45261));
    LocalMux I__10803 (
            .O(N__45266),
            .I(rand_data_29));
    Odrv4 I__10802 (
            .O(N__45261),
            .I(rand_data_29));
    CascadeMux I__10801 (
            .O(N__45256),
            .I(N__45253));
    InMux I__10800 (
            .O(N__45253),
            .I(N__45249));
    InMux I__10799 (
            .O(N__45252),
            .I(N__45245));
    LocalMux I__10798 (
            .O(N__45249),
            .I(N__45242));
    InMux I__10797 (
            .O(N__45248),
            .I(N__45239));
    LocalMux I__10796 (
            .O(N__45245),
            .I(N__45235));
    Span4Mux_v I__10795 (
            .O(N__45242),
            .I(N__45230));
    LocalMux I__10794 (
            .O(N__45239),
            .I(N__45230));
    InMux I__10793 (
            .O(N__45238),
            .I(N__45227));
    Span4Mux_h I__10792 (
            .O(N__45235),
            .I(N__45224));
    Span4Mux_h I__10791 (
            .O(N__45230),
            .I(N__45221));
    LocalMux I__10790 (
            .O(N__45227),
            .I(data_out_frame2_13_5));
    Odrv4 I__10789 (
            .O(N__45224),
            .I(data_out_frame2_13_5));
    Odrv4 I__10788 (
            .O(N__45221),
            .I(data_out_frame2_13_5));
    CascadeMux I__10787 (
            .O(N__45214),
            .I(N__45210));
    InMux I__10786 (
            .O(N__45213),
            .I(N__45207));
    InMux I__10785 (
            .O(N__45210),
            .I(N__45202));
    LocalMux I__10784 (
            .O(N__45207),
            .I(N__45198));
    InMux I__10783 (
            .O(N__45206),
            .I(N__45195));
    InMux I__10782 (
            .O(N__45205),
            .I(N__45192));
    LocalMux I__10781 (
            .O(N__45202),
            .I(N__45188));
    InMux I__10780 (
            .O(N__45201),
            .I(N__45185));
    Span4Mux_v I__10779 (
            .O(N__45198),
            .I(N__45182));
    LocalMux I__10778 (
            .O(N__45195),
            .I(N__45177));
    LocalMux I__10777 (
            .O(N__45192),
            .I(N__45177));
    InMux I__10776 (
            .O(N__45191),
            .I(N__45174));
    Span4Mux_s3_v I__10775 (
            .O(N__45188),
            .I(N__45169));
    LocalMux I__10774 (
            .O(N__45185),
            .I(N__45169));
    Span4Mux_h I__10773 (
            .O(N__45182),
            .I(N__45166));
    Span4Mux_h I__10772 (
            .O(N__45177),
            .I(N__45161));
    LocalMux I__10771 (
            .O(N__45174),
            .I(N__45161));
    Span4Mux_h I__10770 (
            .O(N__45169),
            .I(N__45158));
    Odrv4 I__10769 (
            .O(N__45166),
            .I(\c0.data_out_5_1 ));
    Odrv4 I__10768 (
            .O(N__45161),
            .I(\c0.data_out_5_1 ));
    Odrv4 I__10767 (
            .O(N__45158),
            .I(\c0.data_out_5_1 ));
    InMux I__10766 (
            .O(N__45151),
            .I(N__45148));
    LocalMux I__10765 (
            .O(N__45148),
            .I(N__45145));
    Span4Mux_h I__10764 (
            .O(N__45145),
            .I(N__45141));
    InMux I__10763 (
            .O(N__45144),
            .I(N__45138));
    Odrv4 I__10762 (
            .O(N__45141),
            .I(\c0.n17043 ));
    LocalMux I__10761 (
            .O(N__45138),
            .I(\c0.n17043 ));
    CascadeMux I__10760 (
            .O(N__45133),
            .I(N__45130));
    InMux I__10759 (
            .O(N__45130),
            .I(N__45127));
    LocalMux I__10758 (
            .O(N__45127),
            .I(N__45124));
    Span4Mux_v I__10757 (
            .O(N__45124),
            .I(N__45121));
    Odrv4 I__10756 (
            .O(N__45121),
            .I(\c0.n16949 ));
    InMux I__10755 (
            .O(N__45118),
            .I(N__45115));
    LocalMux I__10754 (
            .O(N__45115),
            .I(N__45111));
    InMux I__10753 (
            .O(N__45114),
            .I(N__45108));
    Span4Mux_v I__10752 (
            .O(N__45111),
            .I(N__45103));
    LocalMux I__10751 (
            .O(N__45108),
            .I(N__45100));
    InMux I__10750 (
            .O(N__45107),
            .I(N__45094));
    InMux I__10749 (
            .O(N__45106),
            .I(N__45094));
    Span4Mux_h I__10748 (
            .O(N__45103),
            .I(N__45089));
    Span4Mux_h I__10747 (
            .O(N__45100),
            .I(N__45089));
    InMux I__10746 (
            .O(N__45099),
            .I(N__45086));
    LocalMux I__10745 (
            .O(N__45094),
            .I(data_out_8_7));
    Odrv4 I__10744 (
            .O(N__45089),
            .I(data_out_8_7));
    LocalMux I__10743 (
            .O(N__45086),
            .I(data_out_8_7));
    InMux I__10742 (
            .O(N__45079),
            .I(N__45076));
    LocalMux I__10741 (
            .O(N__45076),
            .I(N__45071));
    InMux I__10740 (
            .O(N__45075),
            .I(N__45064));
    InMux I__10739 (
            .O(N__45074),
            .I(N__45064));
    Span4Mux_h I__10738 (
            .O(N__45071),
            .I(N__45061));
    InMux I__10737 (
            .O(N__45070),
            .I(N__45058));
    InMux I__10736 (
            .O(N__45069),
            .I(N__45054));
    LocalMux I__10735 (
            .O(N__45064),
            .I(N__45051));
    Span4Mux_h I__10734 (
            .O(N__45061),
            .I(N__45046));
    LocalMux I__10733 (
            .O(N__45058),
            .I(N__45046));
    InMux I__10732 (
            .O(N__45057),
            .I(N__45043));
    LocalMux I__10731 (
            .O(N__45054),
            .I(\c0.data_out_7__3__N_441 ));
    Odrv4 I__10730 (
            .O(N__45051),
            .I(\c0.data_out_7__3__N_441 ));
    Odrv4 I__10729 (
            .O(N__45046),
            .I(\c0.data_out_7__3__N_441 ));
    LocalMux I__10728 (
            .O(N__45043),
            .I(\c0.data_out_7__3__N_441 ));
    InMux I__10727 (
            .O(N__45034),
            .I(N__45031));
    LocalMux I__10726 (
            .O(N__45031),
            .I(N__45028));
    Span4Mux_h I__10725 (
            .O(N__45028),
            .I(N__45025));
    Odrv4 I__10724 (
            .O(N__45025),
            .I(\c0.n10_adj_2276 ));
    InMux I__10723 (
            .O(N__45022),
            .I(N__45017));
    InMux I__10722 (
            .O(N__45021),
            .I(N__45012));
    InMux I__10721 (
            .O(N__45020),
            .I(N__45012));
    LocalMux I__10720 (
            .O(N__45017),
            .I(N__45009));
    LocalMux I__10719 (
            .O(N__45012),
            .I(\c0.data_out_9_3 ));
    Odrv4 I__10718 (
            .O(N__45009),
            .I(\c0.data_out_9_3 ));
    InMux I__10717 (
            .O(N__45004),
            .I(N__45001));
    LocalMux I__10716 (
            .O(N__45001),
            .I(N__44997));
    InMux I__10715 (
            .O(N__45000),
            .I(N__44994));
    Span4Mux_v I__10714 (
            .O(N__44997),
            .I(N__44991));
    LocalMux I__10713 (
            .O(N__44994),
            .I(N__44988));
    Span4Mux_h I__10712 (
            .O(N__44991),
            .I(N__44985));
    Span4Mux_v I__10711 (
            .O(N__44988),
            .I(N__44982));
    Odrv4 I__10710 (
            .O(N__44985),
            .I(\c0.n16981 ));
    Odrv4 I__10709 (
            .O(N__44982),
            .I(\c0.n16981 ));
    InMux I__10708 (
            .O(N__44977),
            .I(N__44974));
    LocalMux I__10707 (
            .O(N__44974),
            .I(N__44970));
    CascadeMux I__10706 (
            .O(N__44973),
            .I(N__44967));
    Span4Mux_v I__10705 (
            .O(N__44970),
            .I(N__44964));
    InMux I__10704 (
            .O(N__44967),
            .I(N__44961));
    Span4Mux_h I__10703 (
            .O(N__44964),
            .I(N__44958));
    LocalMux I__10702 (
            .O(N__44961),
            .I(N__44955));
    Odrv4 I__10701 (
            .O(N__44958),
            .I(\c0.n16969 ));
    Odrv4 I__10700 (
            .O(N__44955),
            .I(\c0.n16969 ));
    InMux I__10699 (
            .O(N__44950),
            .I(N__44947));
    LocalMux I__10698 (
            .O(N__44947),
            .I(N__44940));
    InMux I__10697 (
            .O(N__44946),
            .I(N__44937));
    InMux I__10696 (
            .O(N__44945),
            .I(N__44934));
    InMux I__10695 (
            .O(N__44944),
            .I(N__44931));
    CascadeMux I__10694 (
            .O(N__44943),
            .I(N__44928));
    Span4Mux_v I__10693 (
            .O(N__44940),
            .I(N__44925));
    LocalMux I__10692 (
            .O(N__44937),
            .I(N__44922));
    LocalMux I__10691 (
            .O(N__44934),
            .I(N__44919));
    LocalMux I__10690 (
            .O(N__44931),
            .I(N__44915));
    InMux I__10689 (
            .O(N__44928),
            .I(N__44912));
    Span4Mux_h I__10688 (
            .O(N__44925),
            .I(N__44907));
    Span4Mux_h I__10687 (
            .O(N__44922),
            .I(N__44907));
    Span4Mux_h I__10686 (
            .O(N__44919),
            .I(N__44904));
    InMux I__10685 (
            .O(N__44918),
            .I(N__44901));
    Span12Mux_h I__10684 (
            .O(N__44915),
            .I(N__44896));
    LocalMux I__10683 (
            .O(N__44912),
            .I(N__44896));
    Odrv4 I__10682 (
            .O(N__44907),
            .I(rand_data_15));
    Odrv4 I__10681 (
            .O(N__44904),
            .I(rand_data_15));
    LocalMux I__10680 (
            .O(N__44901),
            .I(rand_data_15));
    Odrv12 I__10679 (
            .O(N__44896),
            .I(rand_data_15));
    InMux I__10678 (
            .O(N__44887),
            .I(N__44883));
    InMux I__10677 (
            .O(N__44886),
            .I(N__44879));
    LocalMux I__10676 (
            .O(N__44883),
            .I(N__44874));
    InMux I__10675 (
            .O(N__44882),
            .I(N__44871));
    LocalMux I__10674 (
            .O(N__44879),
            .I(N__44868));
    InMux I__10673 (
            .O(N__44878),
            .I(N__44863));
    InMux I__10672 (
            .O(N__44877),
            .I(N__44863));
    Odrv12 I__10671 (
            .O(N__44874),
            .I(data_out_frame2_9_7));
    LocalMux I__10670 (
            .O(N__44871),
            .I(data_out_frame2_9_7));
    Odrv4 I__10669 (
            .O(N__44868),
            .I(data_out_frame2_9_7));
    LocalMux I__10668 (
            .O(N__44863),
            .I(data_out_frame2_9_7));
    InMux I__10667 (
            .O(N__44854),
            .I(N__44849));
    InMux I__10666 (
            .O(N__44853),
            .I(N__44846));
    CascadeMux I__10665 (
            .O(N__44852),
            .I(N__44843));
    LocalMux I__10664 (
            .O(N__44849),
            .I(N__44838));
    LocalMux I__10663 (
            .O(N__44846),
            .I(N__44835));
    InMux I__10662 (
            .O(N__44843),
            .I(N__44832));
    InMux I__10661 (
            .O(N__44842),
            .I(N__44829));
    InMux I__10660 (
            .O(N__44841),
            .I(N__44826));
    Span4Mux_h I__10659 (
            .O(N__44838),
            .I(N__44823));
    Span4Mux_h I__10658 (
            .O(N__44835),
            .I(N__44820));
    LocalMux I__10657 (
            .O(N__44832),
            .I(N__44817));
    LocalMux I__10656 (
            .O(N__44829),
            .I(data_out_frame2_9_5));
    LocalMux I__10655 (
            .O(N__44826),
            .I(data_out_frame2_9_5));
    Odrv4 I__10654 (
            .O(N__44823),
            .I(data_out_frame2_9_5));
    Odrv4 I__10653 (
            .O(N__44820),
            .I(data_out_frame2_9_5));
    Odrv4 I__10652 (
            .O(N__44817),
            .I(data_out_frame2_9_5));
    CascadeMux I__10651 (
            .O(N__44806),
            .I(N__44803));
    InMux I__10650 (
            .O(N__44803),
            .I(N__44800));
    LocalMux I__10649 (
            .O(N__44800),
            .I(N__44797));
    Span4Mux_h I__10648 (
            .O(N__44797),
            .I(N__44794));
    Span4Mux_h I__10647 (
            .O(N__44794),
            .I(N__44791));
    Odrv4 I__10646 (
            .O(N__44791),
            .I(\c0.n16926 ));
    InMux I__10645 (
            .O(N__44788),
            .I(N__44785));
    LocalMux I__10644 (
            .O(N__44785),
            .I(N__44779));
    InMux I__10643 (
            .O(N__44784),
            .I(N__44776));
    InMux I__10642 (
            .O(N__44783),
            .I(N__44773));
    InMux I__10641 (
            .O(N__44782),
            .I(N__44770));
    Span4Mux_h I__10640 (
            .O(N__44779),
            .I(N__44765));
    LocalMux I__10639 (
            .O(N__44776),
            .I(N__44765));
    LocalMux I__10638 (
            .O(N__44773),
            .I(N__44762));
    LocalMux I__10637 (
            .O(N__44770),
            .I(N__44758));
    Span4Mux_h I__10636 (
            .O(N__44765),
            .I(N__44755));
    Span4Mux_h I__10635 (
            .O(N__44762),
            .I(N__44752));
    InMux I__10634 (
            .O(N__44761),
            .I(N__44749));
    Span4Mux_s2_v I__10633 (
            .O(N__44758),
            .I(N__44746));
    Odrv4 I__10632 (
            .O(N__44755),
            .I(rand_data_24));
    Odrv4 I__10631 (
            .O(N__44752),
            .I(rand_data_24));
    LocalMux I__10630 (
            .O(N__44749),
            .I(rand_data_24));
    Odrv4 I__10629 (
            .O(N__44746),
            .I(rand_data_24));
    InMux I__10628 (
            .O(N__44737),
            .I(N__44731));
    CascadeMux I__10627 (
            .O(N__44736),
            .I(N__44728));
    InMux I__10626 (
            .O(N__44735),
            .I(N__44723));
    InMux I__10625 (
            .O(N__44734),
            .I(N__44723));
    LocalMux I__10624 (
            .O(N__44731),
            .I(N__44720));
    InMux I__10623 (
            .O(N__44728),
            .I(N__44717));
    LocalMux I__10622 (
            .O(N__44723),
            .I(N__44713));
    Span4Mux_v I__10621 (
            .O(N__44720),
            .I(N__44708));
    LocalMux I__10620 (
            .O(N__44717),
            .I(N__44708));
    InMux I__10619 (
            .O(N__44716),
            .I(N__44705));
    Span4Mux_v I__10618 (
            .O(N__44713),
            .I(N__44700));
    Span4Mux_h I__10617 (
            .O(N__44708),
            .I(N__44700));
    LocalMux I__10616 (
            .O(N__44705),
            .I(data_out_frame2_5_0));
    Odrv4 I__10615 (
            .O(N__44700),
            .I(data_out_frame2_5_0));
    InMux I__10614 (
            .O(N__44695),
            .I(N__44691));
    CascadeMux I__10613 (
            .O(N__44694),
            .I(N__44688));
    LocalMux I__10612 (
            .O(N__44691),
            .I(N__44683));
    InMux I__10611 (
            .O(N__44688),
            .I(N__44680));
    InMux I__10610 (
            .O(N__44687),
            .I(N__44677));
    InMux I__10609 (
            .O(N__44686),
            .I(N__44674));
    Span4Mux_h I__10608 (
            .O(N__44683),
            .I(N__44667));
    LocalMux I__10607 (
            .O(N__44680),
            .I(N__44667));
    LocalMux I__10606 (
            .O(N__44677),
            .I(N__44667));
    LocalMux I__10605 (
            .O(N__44674),
            .I(N__44663));
    Span4Mux_h I__10604 (
            .O(N__44667),
            .I(N__44660));
    InMux I__10603 (
            .O(N__44666),
            .I(N__44657));
    Span4Mux_s2_v I__10602 (
            .O(N__44663),
            .I(N__44654));
    Odrv4 I__10601 (
            .O(N__44660),
            .I(rand_data_25));
    LocalMux I__10600 (
            .O(N__44657),
            .I(rand_data_25));
    Odrv4 I__10599 (
            .O(N__44654),
            .I(rand_data_25));
    InMux I__10598 (
            .O(N__44647),
            .I(N__44643));
    InMux I__10597 (
            .O(N__44646),
            .I(N__44639));
    LocalMux I__10596 (
            .O(N__44643),
            .I(N__44636));
    CascadeMux I__10595 (
            .O(N__44642),
            .I(N__44633));
    LocalMux I__10594 (
            .O(N__44639),
            .I(N__44629));
    Span4Mux_v I__10593 (
            .O(N__44636),
            .I(N__44626));
    InMux I__10592 (
            .O(N__44633),
            .I(N__44621));
    InMux I__10591 (
            .O(N__44632),
            .I(N__44621));
    Odrv12 I__10590 (
            .O(N__44629),
            .I(data_out_frame2_6_5));
    Odrv4 I__10589 (
            .O(N__44626),
            .I(data_out_frame2_6_5));
    LocalMux I__10588 (
            .O(N__44621),
            .I(data_out_frame2_6_5));
    CascadeMux I__10587 (
            .O(N__44614),
            .I(N__44611));
    InMux I__10586 (
            .O(N__44611),
            .I(N__44607));
    InMux I__10585 (
            .O(N__44610),
            .I(N__44602));
    LocalMux I__10584 (
            .O(N__44607),
            .I(N__44599));
    InMux I__10583 (
            .O(N__44606),
            .I(N__44596));
    InMux I__10582 (
            .O(N__44605),
            .I(N__44593));
    LocalMux I__10581 (
            .O(N__44602),
            .I(data_out_frame2_5_5));
    Odrv4 I__10580 (
            .O(N__44599),
            .I(data_out_frame2_5_5));
    LocalMux I__10579 (
            .O(N__44596),
            .I(data_out_frame2_5_5));
    LocalMux I__10578 (
            .O(N__44593),
            .I(data_out_frame2_5_5));
    CascadeMux I__10577 (
            .O(N__44584),
            .I(\c0.n5_adj_2349_cascade_ ));
    InMux I__10576 (
            .O(N__44581),
            .I(N__44578));
    LocalMux I__10575 (
            .O(N__44578),
            .I(N__44575));
    Span4Mux_h I__10574 (
            .O(N__44575),
            .I(N__44572));
    Odrv4 I__10573 (
            .O(N__44572),
            .I(\c0.n6_adj_2280 ));
    InMux I__10572 (
            .O(N__44569),
            .I(N__44563));
    InMux I__10571 (
            .O(N__44568),
            .I(N__44558));
    InMux I__10570 (
            .O(N__44567),
            .I(N__44558));
    CascadeMux I__10569 (
            .O(N__44566),
            .I(N__44554));
    LocalMux I__10568 (
            .O(N__44563),
            .I(N__44551));
    LocalMux I__10567 (
            .O(N__44558),
            .I(N__44548));
    InMux I__10566 (
            .O(N__44557),
            .I(N__44544));
    InMux I__10565 (
            .O(N__44554),
            .I(N__44541));
    Span4Mux_h I__10564 (
            .O(N__44551),
            .I(N__44538));
    Span4Mux_v I__10563 (
            .O(N__44548),
            .I(N__44535));
    InMux I__10562 (
            .O(N__44547),
            .I(N__44532));
    LocalMux I__10561 (
            .O(N__44544),
            .I(N__44527));
    LocalMux I__10560 (
            .O(N__44541),
            .I(N__44527));
    Odrv4 I__10559 (
            .O(N__44538),
            .I(rand_data_13));
    Odrv4 I__10558 (
            .O(N__44535),
            .I(rand_data_13));
    LocalMux I__10557 (
            .O(N__44532),
            .I(rand_data_13));
    Odrv12 I__10556 (
            .O(N__44527),
            .I(rand_data_13));
    InMux I__10555 (
            .O(N__44518),
            .I(N__44515));
    LocalMux I__10554 (
            .O(N__44515),
            .I(N__44512));
    Odrv12 I__10553 (
            .O(N__44512),
            .I(\c0.n6_adj_2278 ));
    InMux I__10552 (
            .O(N__44509),
            .I(N__44506));
    LocalMux I__10551 (
            .O(N__44506),
            .I(N__44503));
    Odrv4 I__10550 (
            .O(N__44503),
            .I(\c0.n18089 ));
    CascadeMux I__10549 (
            .O(N__44500),
            .I(N__44497));
    InMux I__10548 (
            .O(N__44497),
            .I(N__44494));
    LocalMux I__10547 (
            .O(N__44494),
            .I(N__44491));
    Odrv12 I__10546 (
            .O(N__44491),
            .I(\c0.n17561 ));
    InMux I__10545 (
            .O(N__44488),
            .I(N__44484));
    InMux I__10544 (
            .O(N__44487),
            .I(N__44481));
    LocalMux I__10543 (
            .O(N__44484),
            .I(N__44477));
    LocalMux I__10542 (
            .O(N__44481),
            .I(N__44474));
    InMux I__10541 (
            .O(N__44480),
            .I(N__44471));
    Span4Mux_v I__10540 (
            .O(N__44477),
            .I(N__44463));
    Span4Mux_v I__10539 (
            .O(N__44474),
            .I(N__44463));
    LocalMux I__10538 (
            .O(N__44471),
            .I(N__44463));
    InMux I__10537 (
            .O(N__44470),
            .I(N__44459));
    Span4Mux_h I__10536 (
            .O(N__44463),
            .I(N__44456));
    InMux I__10535 (
            .O(N__44462),
            .I(N__44453));
    LocalMux I__10534 (
            .O(N__44459),
            .I(N__44450));
    Odrv4 I__10533 (
            .O(N__44456),
            .I(rand_data_18));
    LocalMux I__10532 (
            .O(N__44453),
            .I(rand_data_18));
    Odrv12 I__10531 (
            .O(N__44450),
            .I(rand_data_18));
    CascadeMux I__10530 (
            .O(N__44443),
            .I(N__44438));
    InMux I__10529 (
            .O(N__44442),
            .I(N__44435));
    InMux I__10528 (
            .O(N__44441),
            .I(N__44431));
    InMux I__10527 (
            .O(N__44438),
            .I(N__44428));
    LocalMux I__10526 (
            .O(N__44435),
            .I(N__44425));
    InMux I__10525 (
            .O(N__44434),
            .I(N__44422));
    LocalMux I__10524 (
            .O(N__44431),
            .I(N__44418));
    LocalMux I__10523 (
            .O(N__44428),
            .I(N__44411));
    Span4Mux_v I__10522 (
            .O(N__44425),
            .I(N__44411));
    LocalMux I__10521 (
            .O(N__44422),
            .I(N__44411));
    InMux I__10520 (
            .O(N__44421),
            .I(N__44408));
    Span4Mux_v I__10519 (
            .O(N__44418),
            .I(N__44405));
    Span4Mux_h I__10518 (
            .O(N__44411),
            .I(N__44402));
    LocalMux I__10517 (
            .O(N__44408),
            .I(data_out_frame2_6_2));
    Odrv4 I__10516 (
            .O(N__44405),
            .I(data_out_frame2_6_2));
    Odrv4 I__10515 (
            .O(N__44402),
            .I(data_out_frame2_6_2));
    InMux I__10514 (
            .O(N__44395),
            .I(N__44390));
    InMux I__10513 (
            .O(N__44394),
            .I(N__44385));
    InMux I__10512 (
            .O(N__44393),
            .I(N__44385));
    LocalMux I__10511 (
            .O(N__44390),
            .I(N__44382));
    LocalMux I__10510 (
            .O(N__44385),
            .I(N__44379));
    Span4Mux_h I__10509 (
            .O(N__44382),
            .I(N__44375));
    Span4Mux_h I__10508 (
            .O(N__44379),
            .I(N__44372));
    InMux I__10507 (
            .O(N__44378),
            .I(N__44369));
    Span4Mux_h I__10506 (
            .O(N__44375),
            .I(N__44366));
    Span4Mux_h I__10505 (
            .O(N__44372),
            .I(N__44363));
    LocalMux I__10504 (
            .O(N__44369),
            .I(data_out_frame2_15_6));
    Odrv4 I__10503 (
            .O(N__44366),
            .I(data_out_frame2_15_6));
    Odrv4 I__10502 (
            .O(N__44363),
            .I(data_out_frame2_15_6));
    InMux I__10501 (
            .O(N__44356),
            .I(N__44351));
    InMux I__10500 (
            .O(N__44355),
            .I(N__44348));
    InMux I__10499 (
            .O(N__44354),
            .I(N__44342));
    LocalMux I__10498 (
            .O(N__44351),
            .I(N__44339));
    LocalMux I__10497 (
            .O(N__44348),
            .I(N__44336));
    InMux I__10496 (
            .O(N__44347),
            .I(N__44333));
    InMux I__10495 (
            .O(N__44346),
            .I(N__44328));
    InMux I__10494 (
            .O(N__44345),
            .I(N__44328));
    LocalMux I__10493 (
            .O(N__44342),
            .I(N__44323));
    Span4Mux_v I__10492 (
            .O(N__44339),
            .I(N__44323));
    Span4Mux_h I__10491 (
            .O(N__44336),
            .I(N__44320));
    LocalMux I__10490 (
            .O(N__44333),
            .I(N__44315));
    LocalMux I__10489 (
            .O(N__44328),
            .I(N__44315));
    Odrv4 I__10488 (
            .O(N__44323),
            .I(data_out_frame2_7_6));
    Odrv4 I__10487 (
            .O(N__44320),
            .I(data_out_frame2_7_6));
    Odrv12 I__10486 (
            .O(N__44315),
            .I(data_out_frame2_7_6));
    InMux I__10485 (
            .O(N__44308),
            .I(N__44304));
    InMux I__10484 (
            .O(N__44307),
            .I(N__44301));
    LocalMux I__10483 (
            .O(N__44304),
            .I(N__44298));
    LocalMux I__10482 (
            .O(N__44301),
            .I(N__44295));
    Sp12to4 I__10481 (
            .O(N__44298),
            .I(N__44292));
    Span4Mux_h I__10480 (
            .O(N__44295),
            .I(N__44289));
    Odrv12 I__10479 (
            .O(N__44292),
            .I(\c0.n17127 ));
    Odrv4 I__10478 (
            .O(N__44289),
            .I(\c0.n17127 ));
    InMux I__10477 (
            .O(N__44284),
            .I(N__44279));
    CascadeMux I__10476 (
            .O(N__44283),
            .I(N__44276));
    InMux I__10475 (
            .O(N__44282),
            .I(N__44273));
    LocalMux I__10474 (
            .O(N__44279),
            .I(N__44269));
    InMux I__10473 (
            .O(N__44276),
            .I(N__44266));
    LocalMux I__10472 (
            .O(N__44273),
            .I(N__44263));
    InMux I__10471 (
            .O(N__44272),
            .I(N__44260));
    Span4Mux_h I__10470 (
            .O(N__44269),
            .I(N__44257));
    LocalMux I__10469 (
            .O(N__44266),
            .I(N__44254));
    Span4Mux_h I__10468 (
            .O(N__44263),
            .I(N__44251));
    LocalMux I__10467 (
            .O(N__44260),
            .I(data_out_frame2_8_7));
    Odrv4 I__10466 (
            .O(N__44257),
            .I(data_out_frame2_8_7));
    Odrv4 I__10465 (
            .O(N__44254),
            .I(data_out_frame2_8_7));
    Odrv4 I__10464 (
            .O(N__44251),
            .I(data_out_frame2_8_7));
    InMux I__10463 (
            .O(N__44242),
            .I(N__44238));
    InMux I__10462 (
            .O(N__44241),
            .I(N__44235));
    LocalMux I__10461 (
            .O(N__44238),
            .I(N__44232));
    LocalMux I__10460 (
            .O(N__44235),
            .I(N__44225));
    Span4Mux_v I__10459 (
            .O(N__44232),
            .I(N__44225));
    InMux I__10458 (
            .O(N__44231),
            .I(N__44222));
    InMux I__10457 (
            .O(N__44230),
            .I(N__44218));
    Span4Mux_v I__10456 (
            .O(N__44225),
            .I(N__44215));
    LocalMux I__10455 (
            .O(N__44222),
            .I(N__44212));
    InMux I__10454 (
            .O(N__44221),
            .I(N__44209));
    LocalMux I__10453 (
            .O(N__44218),
            .I(data_out_frame2_11_6));
    Odrv4 I__10452 (
            .O(N__44215),
            .I(data_out_frame2_11_6));
    Odrv12 I__10451 (
            .O(N__44212),
            .I(data_out_frame2_11_6));
    LocalMux I__10450 (
            .O(N__44209),
            .I(data_out_frame2_11_6));
    InMux I__10449 (
            .O(N__44200),
            .I(N__44197));
    LocalMux I__10448 (
            .O(N__44197),
            .I(N__44192));
    InMux I__10447 (
            .O(N__44196),
            .I(N__44189));
    InMux I__10446 (
            .O(N__44195),
            .I(N__44186));
    Span4Mux_v I__10445 (
            .O(N__44192),
            .I(N__44183));
    LocalMux I__10444 (
            .O(N__44189),
            .I(N__44180));
    LocalMux I__10443 (
            .O(N__44186),
            .I(data_out_frame2_14_7));
    Odrv4 I__10442 (
            .O(N__44183),
            .I(data_out_frame2_14_7));
    Odrv4 I__10441 (
            .O(N__44180),
            .I(data_out_frame2_14_7));
    CascadeMux I__10440 (
            .O(N__44173),
            .I(N__44169));
    InMux I__10439 (
            .O(N__44172),
            .I(N__44166));
    InMux I__10438 (
            .O(N__44169),
            .I(N__44161));
    LocalMux I__10437 (
            .O(N__44166),
            .I(N__44157));
    InMux I__10436 (
            .O(N__44165),
            .I(N__44154));
    CascadeMux I__10435 (
            .O(N__44164),
            .I(N__44151));
    LocalMux I__10434 (
            .O(N__44161),
            .I(N__44148));
    InMux I__10433 (
            .O(N__44160),
            .I(N__44145));
    Span4Mux_v I__10432 (
            .O(N__44157),
            .I(N__44140));
    LocalMux I__10431 (
            .O(N__44154),
            .I(N__44140));
    InMux I__10430 (
            .O(N__44151),
            .I(N__44136));
    Span4Mux_h I__10429 (
            .O(N__44148),
            .I(N__44133));
    LocalMux I__10428 (
            .O(N__44145),
            .I(N__44130));
    Span4Mux_h I__10427 (
            .O(N__44140),
            .I(N__44127));
    InMux I__10426 (
            .O(N__44139),
            .I(N__44124));
    LocalMux I__10425 (
            .O(N__44136),
            .I(N__44121));
    Odrv4 I__10424 (
            .O(N__44133),
            .I(rand_data_12));
    Odrv4 I__10423 (
            .O(N__44130),
            .I(rand_data_12));
    Odrv4 I__10422 (
            .O(N__44127),
            .I(rand_data_12));
    LocalMux I__10421 (
            .O(N__44124),
            .I(rand_data_12));
    Odrv12 I__10420 (
            .O(N__44121),
            .I(rand_data_12));
    CascadeMux I__10419 (
            .O(N__44110),
            .I(N__44107));
    InMux I__10418 (
            .O(N__44107),
            .I(N__44103));
    InMux I__10417 (
            .O(N__44106),
            .I(N__44100));
    LocalMux I__10416 (
            .O(N__44103),
            .I(N__44097));
    LocalMux I__10415 (
            .O(N__44100),
            .I(data_out_frame2_17_4));
    Odrv4 I__10414 (
            .O(N__44097),
            .I(data_out_frame2_17_4));
    InMux I__10413 (
            .O(N__44092),
            .I(N__44087));
    InMux I__10412 (
            .O(N__44091),
            .I(N__44082));
    InMux I__10411 (
            .O(N__44090),
            .I(N__44082));
    LocalMux I__10410 (
            .O(N__44087),
            .I(N__44078));
    LocalMux I__10409 (
            .O(N__44082),
            .I(N__44075));
    InMux I__10408 (
            .O(N__44081),
            .I(N__44072));
    Span4Mux_h I__10407 (
            .O(N__44078),
            .I(N__44069));
    Span4Mux_v I__10406 (
            .O(N__44075),
            .I(N__44065));
    LocalMux I__10405 (
            .O(N__44072),
            .I(N__44062));
    Span4Mux_v I__10404 (
            .O(N__44069),
            .I(N__44059));
    InMux I__10403 (
            .O(N__44068),
            .I(N__44056));
    Span4Mux_h I__10402 (
            .O(N__44065),
            .I(N__44051));
    Span4Mux_s2_v I__10401 (
            .O(N__44062),
            .I(N__44051));
    Odrv4 I__10400 (
            .O(N__44059),
            .I(rand_data_23));
    LocalMux I__10399 (
            .O(N__44056),
            .I(rand_data_23));
    Odrv4 I__10398 (
            .O(N__44051),
            .I(rand_data_23));
    InMux I__10397 (
            .O(N__44044),
            .I(N__44041));
    LocalMux I__10396 (
            .O(N__44041),
            .I(N__44035));
    InMux I__10395 (
            .O(N__44040),
            .I(N__44032));
    InMux I__10394 (
            .O(N__44039),
            .I(N__44029));
    InMux I__10393 (
            .O(N__44038),
            .I(N__44026));
    Span4Mux_h I__10392 (
            .O(N__44035),
            .I(N__44019));
    LocalMux I__10391 (
            .O(N__44032),
            .I(N__44019));
    LocalMux I__10390 (
            .O(N__44029),
            .I(N__44019));
    LocalMux I__10389 (
            .O(N__44026),
            .I(data_out_frame2_6_7));
    Odrv4 I__10388 (
            .O(N__44019),
            .I(data_out_frame2_6_7));
    InMux I__10387 (
            .O(N__44014),
            .I(N__44009));
    InMux I__10386 (
            .O(N__44013),
            .I(N__44006));
    InMux I__10385 (
            .O(N__44012),
            .I(N__44003));
    LocalMux I__10384 (
            .O(N__44009),
            .I(N__43997));
    LocalMux I__10383 (
            .O(N__44006),
            .I(N__43997));
    LocalMux I__10382 (
            .O(N__44003),
            .I(N__43994));
    InMux I__10381 (
            .O(N__44002),
            .I(N__43991));
    Span4Mux_h I__10380 (
            .O(N__43997),
            .I(N__43987));
    Span4Mux_v I__10379 (
            .O(N__43994),
            .I(N__43984));
    LocalMux I__10378 (
            .O(N__43991),
            .I(N__43981));
    InMux I__10377 (
            .O(N__43990),
            .I(N__43978));
    Span4Mux_v I__10376 (
            .O(N__43987),
            .I(N__43973));
    Span4Mux_v I__10375 (
            .O(N__43984),
            .I(N__43973));
    Span4Mux_s2_v I__10374 (
            .O(N__43981),
            .I(N__43970));
    LocalMux I__10373 (
            .O(N__43978),
            .I(rand_data_31));
    Odrv4 I__10372 (
            .O(N__43973),
            .I(rand_data_31));
    Odrv4 I__10371 (
            .O(N__43970),
            .I(rand_data_31));
    InMux I__10370 (
            .O(N__43963),
            .I(N__43960));
    LocalMux I__10369 (
            .O(N__43960),
            .I(N__43955));
    InMux I__10368 (
            .O(N__43959),
            .I(N__43952));
    CascadeMux I__10367 (
            .O(N__43958),
            .I(N__43949));
    Span4Mux_v I__10366 (
            .O(N__43955),
            .I(N__43944));
    LocalMux I__10365 (
            .O(N__43952),
            .I(N__43941));
    InMux I__10364 (
            .O(N__43949),
            .I(N__43938));
    InMux I__10363 (
            .O(N__43948),
            .I(N__43935));
    InMux I__10362 (
            .O(N__43947),
            .I(N__43932));
    Span4Mux_h I__10361 (
            .O(N__43944),
            .I(N__43929));
    Span4Mux_h I__10360 (
            .O(N__43941),
            .I(N__43924));
    LocalMux I__10359 (
            .O(N__43938),
            .I(N__43924));
    LocalMux I__10358 (
            .O(N__43935),
            .I(data_out_frame2_5_7));
    LocalMux I__10357 (
            .O(N__43932),
            .I(data_out_frame2_5_7));
    Odrv4 I__10356 (
            .O(N__43929),
            .I(data_out_frame2_5_7));
    Odrv4 I__10355 (
            .O(N__43924),
            .I(data_out_frame2_5_7));
    InMux I__10354 (
            .O(N__43915),
            .I(N__43912));
    LocalMux I__10353 (
            .O(N__43912),
            .I(\c0.n24_adj_2272 ));
    CascadeMux I__10352 (
            .O(N__43909),
            .I(N__43903));
    CascadeMux I__10351 (
            .O(N__43908),
            .I(N__43899));
    InMux I__10350 (
            .O(N__43907),
            .I(N__43896));
    InMux I__10349 (
            .O(N__43906),
            .I(N__43891));
    InMux I__10348 (
            .O(N__43903),
            .I(N__43891));
    InMux I__10347 (
            .O(N__43902),
            .I(N__43888));
    InMux I__10346 (
            .O(N__43899),
            .I(N__43885));
    LocalMux I__10345 (
            .O(N__43896),
            .I(N__43881));
    LocalMux I__10344 (
            .O(N__43891),
            .I(N__43878));
    LocalMux I__10343 (
            .O(N__43888),
            .I(N__43873));
    LocalMux I__10342 (
            .O(N__43885),
            .I(N__43873));
    InMux I__10341 (
            .O(N__43884),
            .I(N__43870));
    Span4Mux_v I__10340 (
            .O(N__43881),
            .I(N__43867));
    Span4Mux_v I__10339 (
            .O(N__43878),
            .I(N__43864));
    Span4Mux_v I__10338 (
            .O(N__43873),
            .I(N__43861));
    LocalMux I__10337 (
            .O(N__43870),
            .I(N__43852));
    Span4Mux_h I__10336 (
            .O(N__43867),
            .I(N__43852));
    Span4Mux_h I__10335 (
            .O(N__43864),
            .I(N__43852));
    Span4Mux_v I__10334 (
            .O(N__43861),
            .I(N__43852));
    Odrv4 I__10333 (
            .O(N__43852),
            .I(data_out_frame2_9_2));
    InMux I__10332 (
            .O(N__43849),
            .I(N__43844));
    InMux I__10331 (
            .O(N__43848),
            .I(N__43841));
    InMux I__10330 (
            .O(N__43847),
            .I(N__43838));
    LocalMux I__10329 (
            .O(N__43844),
            .I(N__43833));
    LocalMux I__10328 (
            .O(N__43841),
            .I(N__43833));
    LocalMux I__10327 (
            .O(N__43838),
            .I(N__43828));
    Sp12to4 I__10326 (
            .O(N__43833),
            .I(N__43825));
    InMux I__10325 (
            .O(N__43832),
            .I(N__43822));
    InMux I__10324 (
            .O(N__43831),
            .I(N__43819));
    Span4Mux_h I__10323 (
            .O(N__43828),
            .I(N__43816));
    Span12Mux_v I__10322 (
            .O(N__43825),
            .I(N__43811));
    LocalMux I__10321 (
            .O(N__43822),
            .I(N__43811));
    LocalMux I__10320 (
            .O(N__43819),
            .I(data_out_frame2_16_0));
    Odrv4 I__10319 (
            .O(N__43816),
            .I(data_out_frame2_16_0));
    Odrv12 I__10318 (
            .O(N__43811),
            .I(data_out_frame2_16_0));
    InMux I__10317 (
            .O(N__43804),
            .I(N__43801));
    LocalMux I__10316 (
            .O(N__43801),
            .I(N__43798));
    Odrv4 I__10315 (
            .O(N__43798),
            .I(\c0.n9892 ));
    CascadeMux I__10314 (
            .O(N__43795),
            .I(N__43792));
    InMux I__10313 (
            .O(N__43792),
            .I(N__43789));
    LocalMux I__10312 (
            .O(N__43789),
            .I(N__43786));
    Odrv4 I__10311 (
            .O(N__43786),
            .I(\c0.n20_adj_2205 ));
    InMux I__10310 (
            .O(N__43783),
            .I(N__43780));
    LocalMux I__10309 (
            .O(N__43780),
            .I(N__43777));
    Odrv12 I__10308 (
            .O(N__43777),
            .I(\c0.n18071 ));
    CascadeMux I__10307 (
            .O(N__43774),
            .I(\c0.n18074_cascade_ ));
    InMux I__10306 (
            .O(N__43771),
            .I(N__43768));
    LocalMux I__10305 (
            .O(N__43768),
            .I(N__43763));
    InMux I__10304 (
            .O(N__43767),
            .I(N__43760));
    InMux I__10303 (
            .O(N__43766),
            .I(N__43757));
    Span4Mux_v I__10302 (
            .O(N__43763),
            .I(N__43753));
    LocalMux I__10301 (
            .O(N__43760),
            .I(N__43750));
    LocalMux I__10300 (
            .O(N__43757),
            .I(N__43747));
    InMux I__10299 (
            .O(N__43756),
            .I(N__43744));
    Span4Mux_h I__10298 (
            .O(N__43753),
            .I(N__43739));
    Span4Mux_v I__10297 (
            .O(N__43750),
            .I(N__43739));
    Odrv12 I__10296 (
            .O(N__43747),
            .I(data_out_frame2_12_7));
    LocalMux I__10295 (
            .O(N__43744),
            .I(data_out_frame2_12_7));
    Odrv4 I__10294 (
            .O(N__43739),
            .I(data_out_frame2_12_7));
    InMux I__10293 (
            .O(N__43732),
            .I(N__43729));
    LocalMux I__10292 (
            .O(N__43729),
            .I(N__43725));
    CascadeMux I__10291 (
            .O(N__43728),
            .I(N__43721));
    Span4Mux_v I__10290 (
            .O(N__43725),
            .I(N__43718));
    InMux I__10289 (
            .O(N__43724),
            .I(N__43715));
    InMux I__10288 (
            .O(N__43721),
            .I(N__43712));
    Span4Mux_h I__10287 (
            .O(N__43718),
            .I(N__43709));
    LocalMux I__10286 (
            .O(N__43715),
            .I(N__43704));
    LocalMux I__10285 (
            .O(N__43712),
            .I(N__43704));
    Odrv4 I__10284 (
            .O(N__43709),
            .I(data_out_frame2_13_7));
    Odrv4 I__10283 (
            .O(N__43704),
            .I(data_out_frame2_13_7));
    CascadeMux I__10282 (
            .O(N__43699),
            .I(\c0.n18065_cascade_ ));
    InMux I__10281 (
            .O(N__43696),
            .I(N__43693));
    LocalMux I__10280 (
            .O(N__43693),
            .I(\c0.n18068 ));
    InMux I__10279 (
            .O(N__43690),
            .I(N__43687));
    LocalMux I__10278 (
            .O(N__43687),
            .I(N__43683));
    InMux I__10277 (
            .O(N__43686),
            .I(N__43679));
    Span4Mux_h I__10276 (
            .O(N__43683),
            .I(N__43675));
    InMux I__10275 (
            .O(N__43682),
            .I(N__43672));
    LocalMux I__10274 (
            .O(N__43679),
            .I(N__43669));
    InMux I__10273 (
            .O(N__43678),
            .I(N__43666));
    Sp12to4 I__10272 (
            .O(N__43675),
            .I(N__43663));
    LocalMux I__10271 (
            .O(N__43672),
            .I(N__43658));
    Span4Mux_h I__10270 (
            .O(N__43669),
            .I(N__43658));
    LocalMux I__10269 (
            .O(N__43666),
            .I(data_out_frame2_14_6));
    Odrv12 I__10268 (
            .O(N__43663),
            .I(data_out_frame2_14_6));
    Odrv4 I__10267 (
            .O(N__43658),
            .I(data_out_frame2_14_6));
    InMux I__10266 (
            .O(N__43651),
            .I(N__43648));
    LocalMux I__10265 (
            .O(N__43648),
            .I(N__43643));
    InMux I__10264 (
            .O(N__43647),
            .I(N__43640));
    InMux I__10263 (
            .O(N__43646),
            .I(N__43637));
    Span4Mux_h I__10262 (
            .O(N__43643),
            .I(N__43633));
    LocalMux I__10261 (
            .O(N__43640),
            .I(N__43630));
    LocalMux I__10260 (
            .O(N__43637),
            .I(N__43627));
    InMux I__10259 (
            .O(N__43636),
            .I(N__43623));
    Span4Mux_v I__10258 (
            .O(N__43633),
            .I(N__43620));
    Span4Mux_h I__10257 (
            .O(N__43630),
            .I(N__43617));
    Span4Mux_h I__10256 (
            .O(N__43627),
            .I(N__43614));
    InMux I__10255 (
            .O(N__43626),
            .I(N__43611));
    LocalMux I__10254 (
            .O(N__43623),
            .I(data_out_frame2_12_6));
    Odrv4 I__10253 (
            .O(N__43620),
            .I(data_out_frame2_12_6));
    Odrv4 I__10252 (
            .O(N__43617),
            .I(data_out_frame2_12_6));
    Odrv4 I__10251 (
            .O(N__43614),
            .I(data_out_frame2_12_6));
    LocalMux I__10250 (
            .O(N__43611),
            .I(data_out_frame2_12_6));
    CascadeMux I__10249 (
            .O(N__43600),
            .I(\c0.n18005_cascade_ ));
    CascadeMux I__10248 (
            .O(N__43597),
            .I(N__43594));
    InMux I__10247 (
            .O(N__43594),
            .I(N__43591));
    LocalMux I__10246 (
            .O(N__43591),
            .I(N__43588));
    Odrv4 I__10245 (
            .O(N__43588),
            .I(\c0.n18008 ));
    InMux I__10244 (
            .O(N__43585),
            .I(N__43581));
    InMux I__10243 (
            .O(N__43584),
            .I(N__43578));
    LocalMux I__10242 (
            .O(N__43581),
            .I(N__43575));
    LocalMux I__10241 (
            .O(N__43578),
            .I(N__43569));
    Span4Mux_v I__10240 (
            .O(N__43575),
            .I(N__43566));
    InMux I__10239 (
            .O(N__43574),
            .I(N__43563));
    InMux I__10238 (
            .O(N__43573),
            .I(N__43560));
    InMux I__10237 (
            .O(N__43572),
            .I(N__43557));
    Span4Mux_v I__10236 (
            .O(N__43569),
            .I(N__43554));
    Span4Mux_h I__10235 (
            .O(N__43566),
            .I(N__43549));
    LocalMux I__10234 (
            .O(N__43563),
            .I(N__43549));
    LocalMux I__10233 (
            .O(N__43560),
            .I(N__43546));
    LocalMux I__10232 (
            .O(N__43557),
            .I(data_out_frame2_10_0));
    Odrv4 I__10231 (
            .O(N__43554),
            .I(data_out_frame2_10_0));
    Odrv4 I__10230 (
            .O(N__43549),
            .I(data_out_frame2_10_0));
    Odrv4 I__10229 (
            .O(N__43546),
            .I(data_out_frame2_10_0));
    InMux I__10228 (
            .O(N__43537),
            .I(N__43534));
    LocalMux I__10227 (
            .O(N__43534),
            .I(N__43531));
    Span4Mux_v I__10226 (
            .O(N__43531),
            .I(N__43528));
    Odrv4 I__10225 (
            .O(N__43528),
            .I(\c0.n17347 ));
    InMux I__10224 (
            .O(N__43525),
            .I(N__43520));
    InMux I__10223 (
            .O(N__43524),
            .I(N__43516));
    InMux I__10222 (
            .O(N__43523),
            .I(N__43513));
    LocalMux I__10221 (
            .O(N__43520),
            .I(N__43510));
    InMux I__10220 (
            .O(N__43519),
            .I(N__43507));
    LocalMux I__10219 (
            .O(N__43516),
            .I(N__43504));
    LocalMux I__10218 (
            .O(N__43513),
            .I(N__43501));
    Span4Mux_h I__10217 (
            .O(N__43510),
            .I(N__43498));
    LocalMux I__10216 (
            .O(N__43507),
            .I(data_out_frame2_5_4));
    Odrv4 I__10215 (
            .O(N__43504),
            .I(data_out_frame2_5_4));
    Odrv12 I__10214 (
            .O(N__43501),
            .I(data_out_frame2_5_4));
    Odrv4 I__10213 (
            .O(N__43498),
            .I(data_out_frame2_5_4));
    InMux I__10212 (
            .O(N__43489),
            .I(N__43486));
    LocalMux I__10211 (
            .O(N__43486),
            .I(N__43483));
    Span4Mux_v I__10210 (
            .O(N__43483),
            .I(N__43480));
    Odrv4 I__10209 (
            .O(N__43480),
            .I(\c0.n17495 ));
    InMux I__10208 (
            .O(N__43477),
            .I(N__43474));
    LocalMux I__10207 (
            .O(N__43474),
            .I(N__43469));
    InMux I__10206 (
            .O(N__43473),
            .I(N__43466));
    InMux I__10205 (
            .O(N__43472),
            .I(N__43460));
    Span4Mux_v I__10204 (
            .O(N__43469),
            .I(N__43457));
    LocalMux I__10203 (
            .O(N__43466),
            .I(N__43454));
    InMux I__10202 (
            .O(N__43465),
            .I(N__43451));
    InMux I__10201 (
            .O(N__43464),
            .I(N__43448));
    InMux I__10200 (
            .O(N__43463),
            .I(N__43445));
    LocalMux I__10199 (
            .O(N__43460),
            .I(N__43438));
    Span4Mux_h I__10198 (
            .O(N__43457),
            .I(N__43438));
    Span4Mux_v I__10197 (
            .O(N__43454),
            .I(N__43438));
    LocalMux I__10196 (
            .O(N__43451),
            .I(N__43433));
    LocalMux I__10195 (
            .O(N__43448),
            .I(N__43433));
    LocalMux I__10194 (
            .O(N__43445),
            .I(N__43430));
    Sp12to4 I__10193 (
            .O(N__43438),
            .I(N__43427));
    Span4Mux_h I__10192 (
            .O(N__43433),
            .I(N__43424));
    Odrv12 I__10191 (
            .O(N__43430),
            .I(data_out_frame2_9_6));
    Odrv12 I__10190 (
            .O(N__43427),
            .I(data_out_frame2_9_6));
    Odrv4 I__10189 (
            .O(N__43424),
            .I(data_out_frame2_9_6));
    InMux I__10188 (
            .O(N__43417),
            .I(N__43414));
    LocalMux I__10187 (
            .O(N__43414),
            .I(\c0.n18047 ));
    InMux I__10186 (
            .O(N__43411),
            .I(N__43407));
    InMux I__10185 (
            .O(N__43410),
            .I(N__43404));
    LocalMux I__10184 (
            .O(N__43407),
            .I(N__43401));
    LocalMux I__10183 (
            .O(N__43404),
            .I(N__43398));
    Span4Mux_h I__10182 (
            .O(N__43401),
            .I(N__43395));
    Span4Mux_v I__10181 (
            .O(N__43398),
            .I(N__43392));
    Odrv4 I__10180 (
            .O(N__43395),
            .I(\c0.n9859 ));
    Odrv4 I__10179 (
            .O(N__43392),
            .I(\c0.n9859 ));
    CascadeMux I__10178 (
            .O(N__43387),
            .I(N__43384));
    InMux I__10177 (
            .O(N__43384),
            .I(N__43381));
    LocalMux I__10176 (
            .O(N__43381),
            .I(N__43377));
    InMux I__10175 (
            .O(N__43380),
            .I(N__43374));
    Span4Mux_v I__10174 (
            .O(N__43377),
            .I(N__43369));
    LocalMux I__10173 (
            .O(N__43374),
            .I(N__43366));
    InMux I__10172 (
            .O(N__43373),
            .I(N__43363));
    InMux I__10171 (
            .O(N__43372),
            .I(N__43360));
    Span4Mux_v I__10170 (
            .O(N__43369),
            .I(N__43357));
    Span4Mux_v I__10169 (
            .O(N__43366),
            .I(N__43354));
    LocalMux I__10168 (
            .O(N__43363),
            .I(N__43351));
    LocalMux I__10167 (
            .O(N__43360),
            .I(N__43346));
    Span4Mux_h I__10166 (
            .O(N__43357),
            .I(N__43346));
    Span4Mux_h I__10165 (
            .O(N__43354),
            .I(N__43341));
    Span4Mux_v I__10164 (
            .O(N__43351),
            .I(N__43341));
    Odrv4 I__10163 (
            .O(N__43346),
            .I(data_out_frame2_13_2));
    Odrv4 I__10162 (
            .O(N__43341),
            .I(data_out_frame2_13_2));
    InMux I__10161 (
            .O(N__43336),
            .I(N__43332));
    InMux I__10160 (
            .O(N__43335),
            .I(N__43329));
    LocalMux I__10159 (
            .O(N__43332),
            .I(N__43324));
    LocalMux I__10158 (
            .O(N__43329),
            .I(N__43324));
    Span4Mux_h I__10157 (
            .O(N__43324),
            .I(N__43321));
    Odrv4 I__10156 (
            .O(N__43321),
            .I(\c0.n17133 ));
    InMux I__10155 (
            .O(N__43318),
            .I(N__43315));
    LocalMux I__10154 (
            .O(N__43315),
            .I(N__43312));
    Odrv4 I__10153 (
            .O(N__43312),
            .I(\c0.n27_adj_2277 ));
    InMux I__10152 (
            .O(N__43309),
            .I(N__43306));
    LocalMux I__10151 (
            .O(N__43306),
            .I(N__43301));
    CascadeMux I__10150 (
            .O(N__43305),
            .I(N__43297));
    InMux I__10149 (
            .O(N__43304),
            .I(N__43294));
    Span4Mux_v I__10148 (
            .O(N__43301),
            .I(N__43291));
    InMux I__10147 (
            .O(N__43300),
            .I(N__43286));
    InMux I__10146 (
            .O(N__43297),
            .I(N__43286));
    LocalMux I__10145 (
            .O(N__43294),
            .I(data_out_frame2_8_6));
    Odrv4 I__10144 (
            .O(N__43291),
            .I(data_out_frame2_8_6));
    LocalMux I__10143 (
            .O(N__43286),
            .I(data_out_frame2_8_6));
    InMux I__10142 (
            .O(N__43279),
            .I(N__43274));
    InMux I__10141 (
            .O(N__43278),
            .I(N__43271));
    InMux I__10140 (
            .O(N__43277),
            .I(N__43268));
    LocalMux I__10139 (
            .O(N__43274),
            .I(N__43263));
    LocalMux I__10138 (
            .O(N__43271),
            .I(N__43258));
    LocalMux I__10137 (
            .O(N__43268),
            .I(N__43258));
    CascadeMux I__10136 (
            .O(N__43267),
            .I(N__43255));
    InMux I__10135 (
            .O(N__43266),
            .I(N__43252));
    Span4Mux_h I__10134 (
            .O(N__43263),
            .I(N__43247));
    Span4Mux_h I__10133 (
            .O(N__43258),
            .I(N__43247));
    InMux I__10132 (
            .O(N__43255),
            .I(N__43244));
    LocalMux I__10131 (
            .O(N__43252),
            .I(data_out_frame2_6_6));
    Odrv4 I__10130 (
            .O(N__43247),
            .I(data_out_frame2_6_6));
    LocalMux I__10129 (
            .O(N__43244),
            .I(data_out_frame2_6_6));
    InMux I__10128 (
            .O(N__43237),
            .I(N__43234));
    LocalMux I__10127 (
            .O(N__43234),
            .I(\c0.n18050 ));
    InMux I__10126 (
            .O(N__43231),
            .I(N__43228));
    LocalMux I__10125 (
            .O(N__43228),
            .I(N__43224));
    InMux I__10124 (
            .O(N__43227),
            .I(N__43221));
    Odrv4 I__10123 (
            .O(N__43224),
            .I(\c0.n9671 ));
    LocalMux I__10122 (
            .O(N__43221),
            .I(\c0.n9671 ));
    InMux I__10121 (
            .O(N__43216),
            .I(N__43212));
    InMux I__10120 (
            .O(N__43215),
            .I(N__43209));
    LocalMux I__10119 (
            .O(N__43212),
            .I(\c0.n17016 ));
    LocalMux I__10118 (
            .O(N__43209),
            .I(\c0.n17016 ));
    InMux I__10117 (
            .O(N__43204),
            .I(N__43201));
    LocalMux I__10116 (
            .O(N__43201),
            .I(N__43198));
    Span4Mux_h I__10115 (
            .O(N__43198),
            .I(N__43195));
    Span4Mux_h I__10114 (
            .O(N__43195),
            .I(N__43192));
    Odrv4 I__10113 (
            .O(N__43192),
            .I(\c0.n6_adj_2293 ));
    InMux I__10112 (
            .O(N__43189),
            .I(N__43186));
    LocalMux I__10111 (
            .O(N__43186),
            .I(N__43183));
    Span4Mux_h I__10110 (
            .O(N__43183),
            .I(N__43179));
    InMux I__10109 (
            .O(N__43182),
            .I(N__43176));
    Odrv4 I__10108 (
            .O(N__43179),
            .I(\c0.n16960 ));
    LocalMux I__10107 (
            .O(N__43176),
            .I(\c0.n16960 ));
    CascadeMux I__10106 (
            .O(N__43171),
            .I(\c0.n18017_cascade_ ));
    InMux I__10105 (
            .O(N__43168),
            .I(N__43165));
    LocalMux I__10104 (
            .O(N__43165),
            .I(\c0.n17593 ));
    InMux I__10103 (
            .O(N__43162),
            .I(N__43159));
    LocalMux I__10102 (
            .O(N__43159),
            .I(\c0.n10_adj_2154 ));
    CascadeMux I__10101 (
            .O(N__43156),
            .I(\c0.n18020_cascade_ ));
    InMux I__10100 (
            .O(N__43153),
            .I(N__43143));
    InMux I__10099 (
            .O(N__43152),
            .I(N__43140));
    InMux I__10098 (
            .O(N__43151),
            .I(N__43136));
    InMux I__10097 (
            .O(N__43150),
            .I(N__43133));
    InMux I__10096 (
            .O(N__43149),
            .I(N__43130));
    InMux I__10095 (
            .O(N__43148),
            .I(N__43127));
    InMux I__10094 (
            .O(N__43147),
            .I(N__43124));
    InMux I__10093 (
            .O(N__43146),
            .I(N__43121));
    LocalMux I__10092 (
            .O(N__43143),
            .I(N__43116));
    LocalMux I__10091 (
            .O(N__43140),
            .I(N__43113));
    CascadeMux I__10090 (
            .O(N__43139),
            .I(N__43109));
    LocalMux I__10089 (
            .O(N__43136),
            .I(N__43106));
    LocalMux I__10088 (
            .O(N__43133),
            .I(N__43103));
    LocalMux I__10087 (
            .O(N__43130),
            .I(N__43096));
    LocalMux I__10086 (
            .O(N__43127),
            .I(N__43096));
    LocalMux I__10085 (
            .O(N__43124),
            .I(N__43096));
    LocalMux I__10084 (
            .O(N__43121),
            .I(N__43093));
    InMux I__10083 (
            .O(N__43120),
            .I(N__43090));
    InMux I__10082 (
            .O(N__43119),
            .I(N__43087));
    Span4Mux_v I__10081 (
            .O(N__43116),
            .I(N__43082));
    Span4Mux_v I__10080 (
            .O(N__43113),
            .I(N__43082));
    InMux I__10079 (
            .O(N__43112),
            .I(N__43079));
    InMux I__10078 (
            .O(N__43109),
            .I(N__43075));
    Span4Mux_s1_v I__10077 (
            .O(N__43106),
            .I(N__43072));
    Span4Mux_h I__10076 (
            .O(N__43103),
            .I(N__43069));
    Span4Mux_v I__10075 (
            .O(N__43096),
            .I(N__43064));
    Span4Mux_s1_v I__10074 (
            .O(N__43093),
            .I(N__43064));
    LocalMux I__10073 (
            .O(N__43090),
            .I(N__43055));
    LocalMux I__10072 (
            .O(N__43087),
            .I(N__43055));
    Sp12to4 I__10071 (
            .O(N__43082),
            .I(N__43055));
    LocalMux I__10070 (
            .O(N__43079),
            .I(N__43055));
    InMux I__10069 (
            .O(N__43078),
            .I(N__43052));
    LocalMux I__10068 (
            .O(N__43075),
            .I(byte_transmit_counter_3));
    Odrv4 I__10067 (
            .O(N__43072),
            .I(byte_transmit_counter_3));
    Odrv4 I__10066 (
            .O(N__43069),
            .I(byte_transmit_counter_3));
    Odrv4 I__10065 (
            .O(N__43064),
            .I(byte_transmit_counter_3));
    Odrv12 I__10064 (
            .O(N__43055),
            .I(byte_transmit_counter_3));
    LocalMux I__10063 (
            .O(N__43052),
            .I(byte_transmit_counter_3));
    InMux I__10062 (
            .O(N__43039),
            .I(N__43036));
    LocalMux I__10061 (
            .O(N__43036),
            .I(N__43033));
    Odrv12 I__10060 (
            .O(N__43033),
            .I(\c0.n10_adj_2155 ));
    InMux I__10059 (
            .O(N__43030),
            .I(N__43027));
    LocalMux I__10058 (
            .O(N__43027),
            .I(N__43024));
    Odrv4 I__10057 (
            .O(N__43024),
            .I(\c0.n10_adj_2268 ));
    InMux I__10056 (
            .O(N__43021),
            .I(N__43017));
    InMux I__10055 (
            .O(N__43020),
            .I(N__43014));
    LocalMux I__10054 (
            .O(N__43017),
            .I(N__43008));
    LocalMux I__10053 (
            .O(N__43014),
            .I(N__43005));
    InMux I__10052 (
            .O(N__43013),
            .I(N__43002));
    InMux I__10051 (
            .O(N__43012),
            .I(N__42999));
    InMux I__10050 (
            .O(N__43011),
            .I(N__42996));
    Span4Mux_s3_v I__10049 (
            .O(N__43008),
            .I(N__42989));
    Span4Mux_v I__10048 (
            .O(N__43005),
            .I(N__42989));
    LocalMux I__10047 (
            .O(N__43002),
            .I(N__42989));
    LocalMux I__10046 (
            .O(N__42999),
            .I(\c0.data_out_8_3 ));
    LocalMux I__10045 (
            .O(N__42996),
            .I(\c0.data_out_8_3 ));
    Odrv4 I__10044 (
            .O(N__42989),
            .I(\c0.data_out_8_3 ));
    CascadeMux I__10043 (
            .O(N__42982),
            .I(N__42978));
    InMux I__10042 (
            .O(N__42981),
            .I(N__42975));
    InMux I__10041 (
            .O(N__42978),
            .I(N__42972));
    LocalMux I__10040 (
            .O(N__42975),
            .I(N__42969));
    LocalMux I__10039 (
            .O(N__42972),
            .I(N__42965));
    Span4Mux_s3_v I__10038 (
            .O(N__42969),
            .I(N__42962));
    InMux I__10037 (
            .O(N__42968),
            .I(N__42959));
    Span4Mux_h I__10036 (
            .O(N__42965),
            .I(N__42954));
    Span4Mux_h I__10035 (
            .O(N__42962),
            .I(N__42949));
    LocalMux I__10034 (
            .O(N__42959),
            .I(N__42949));
    InMux I__10033 (
            .O(N__42958),
            .I(N__42944));
    InMux I__10032 (
            .O(N__42957),
            .I(N__42944));
    Odrv4 I__10031 (
            .O(N__42954),
            .I(data_out_8_4));
    Odrv4 I__10030 (
            .O(N__42949),
            .I(data_out_8_4));
    LocalMux I__10029 (
            .O(N__42944),
            .I(data_out_8_4));
    InMux I__10028 (
            .O(N__42937),
            .I(N__42933));
    InMux I__10027 (
            .O(N__42936),
            .I(N__42930));
    LocalMux I__10026 (
            .O(N__42933),
            .I(N__42927));
    LocalMux I__10025 (
            .O(N__42930),
            .I(N__42922));
    Span4Mux_s2_v I__10024 (
            .O(N__42927),
            .I(N__42922));
    Span4Mux_h I__10023 (
            .O(N__42922),
            .I(N__42918));
    InMux I__10022 (
            .O(N__42921),
            .I(N__42915));
    Odrv4 I__10021 (
            .O(N__42918),
            .I(\c0.data_out_9_1 ));
    LocalMux I__10020 (
            .O(N__42915),
            .I(\c0.data_out_9_1 ));
    InMux I__10019 (
            .O(N__42910),
            .I(N__42906));
    InMux I__10018 (
            .O(N__42909),
            .I(N__42903));
    LocalMux I__10017 (
            .O(N__42906),
            .I(data_out_3_4));
    LocalMux I__10016 (
            .O(N__42903),
            .I(data_out_3_4));
    InMux I__10015 (
            .O(N__42898),
            .I(N__42895));
    LocalMux I__10014 (
            .O(N__42895),
            .I(N__42892));
    Span4Mux_s2_v I__10013 (
            .O(N__42892),
            .I(N__42889));
    Span4Mux_h I__10012 (
            .O(N__42889),
            .I(N__42886));
    Odrv4 I__10011 (
            .O(N__42886),
            .I(\c0.n17591 ));
    InMux I__10010 (
            .O(N__42883),
            .I(N__42879));
    CascadeMux I__10009 (
            .O(N__42882),
            .I(N__42876));
    LocalMux I__10008 (
            .O(N__42879),
            .I(N__42873));
    InMux I__10007 (
            .O(N__42876),
            .I(N__42870));
    Odrv4 I__10006 (
            .O(N__42873),
            .I(rand_setpoint_16));
    LocalMux I__10005 (
            .O(N__42870),
            .I(rand_setpoint_16));
    InMux I__10004 (
            .O(N__42865),
            .I(N__42855));
    InMux I__10003 (
            .O(N__42864),
            .I(N__42855));
    InMux I__10002 (
            .O(N__42863),
            .I(N__42852));
    CascadeMux I__10001 (
            .O(N__42862),
            .I(N__42848));
    CascadeMux I__10000 (
            .O(N__42861),
            .I(N__42844));
    CascadeMux I__9999 (
            .O(N__42860),
            .I(N__42839));
    LocalMux I__9998 (
            .O(N__42855),
            .I(N__42835));
    LocalMux I__9997 (
            .O(N__42852),
            .I(N__42832));
    InMux I__9996 (
            .O(N__42851),
            .I(N__42829));
    InMux I__9995 (
            .O(N__42848),
            .I(N__42826));
    InMux I__9994 (
            .O(N__42847),
            .I(N__42823));
    InMux I__9993 (
            .O(N__42844),
            .I(N__42817));
    InMux I__9992 (
            .O(N__42843),
            .I(N__42817));
    InMux I__9991 (
            .O(N__42842),
            .I(N__42812));
    InMux I__9990 (
            .O(N__42839),
            .I(N__42812));
    InMux I__9989 (
            .O(N__42838),
            .I(N__42809));
    Span4Mux_s3_v I__9988 (
            .O(N__42835),
            .I(N__42804));
    Span4Mux_s3_v I__9987 (
            .O(N__42832),
            .I(N__42804));
    LocalMux I__9986 (
            .O(N__42829),
            .I(N__42799));
    LocalMux I__9985 (
            .O(N__42826),
            .I(N__42799));
    LocalMux I__9984 (
            .O(N__42823),
            .I(N__42795));
    InMux I__9983 (
            .O(N__42822),
            .I(N__42792));
    LocalMux I__9982 (
            .O(N__42817),
            .I(N__42781));
    LocalMux I__9981 (
            .O(N__42812),
            .I(N__42781));
    LocalMux I__9980 (
            .O(N__42809),
            .I(N__42781));
    Span4Mux_v I__9979 (
            .O(N__42804),
            .I(N__42781));
    Span4Mux_s3_v I__9978 (
            .O(N__42799),
            .I(N__42781));
    InMux I__9977 (
            .O(N__42798),
            .I(N__42778));
    Span4Mux_v I__9976 (
            .O(N__42795),
            .I(N__42775));
    LocalMux I__9975 (
            .O(N__42792),
            .I(N__42770));
    Span4Mux_h I__9974 (
            .O(N__42781),
            .I(N__42770));
    LocalMux I__9973 (
            .O(N__42778),
            .I(n2547));
    Odrv4 I__9972 (
            .O(N__42775),
            .I(n2547));
    Odrv4 I__9971 (
            .O(N__42770),
            .I(n2547));
    CascadeMux I__9970 (
            .O(N__42763),
            .I(N__42755));
    CascadeMux I__9969 (
            .O(N__42762),
            .I(N__42746));
    CascadeMux I__9968 (
            .O(N__42761),
            .I(N__42742));
    InMux I__9967 (
            .O(N__42760),
            .I(N__42739));
    InMux I__9966 (
            .O(N__42759),
            .I(N__42736));
    InMux I__9965 (
            .O(N__42758),
            .I(N__42733));
    InMux I__9964 (
            .O(N__42755),
            .I(N__42728));
    InMux I__9963 (
            .O(N__42754),
            .I(N__42728));
    InMux I__9962 (
            .O(N__42753),
            .I(N__42722));
    InMux I__9961 (
            .O(N__42752),
            .I(N__42719));
    CascadeMux I__9960 (
            .O(N__42751),
            .I(N__42716));
    CascadeMux I__9959 (
            .O(N__42750),
            .I(N__42713));
    CascadeMux I__9958 (
            .O(N__42749),
            .I(N__42705));
    InMux I__9957 (
            .O(N__42746),
            .I(N__42702));
    InMux I__9956 (
            .O(N__42745),
            .I(N__42698));
    InMux I__9955 (
            .O(N__42742),
            .I(N__42695));
    LocalMux I__9954 (
            .O(N__42739),
            .I(N__42692));
    LocalMux I__9953 (
            .O(N__42736),
            .I(N__42687));
    LocalMux I__9952 (
            .O(N__42733),
            .I(N__42687));
    LocalMux I__9951 (
            .O(N__42728),
            .I(N__42684));
    InMux I__9950 (
            .O(N__42727),
            .I(N__42681));
    InMux I__9949 (
            .O(N__42726),
            .I(N__42675));
    InMux I__9948 (
            .O(N__42725),
            .I(N__42675));
    LocalMux I__9947 (
            .O(N__42722),
            .I(N__42670));
    LocalMux I__9946 (
            .O(N__42719),
            .I(N__42670));
    InMux I__9945 (
            .O(N__42716),
            .I(N__42661));
    InMux I__9944 (
            .O(N__42713),
            .I(N__42661));
    InMux I__9943 (
            .O(N__42712),
            .I(N__42661));
    InMux I__9942 (
            .O(N__42711),
            .I(N__42661));
    InMux I__9941 (
            .O(N__42710),
            .I(N__42657));
    InMux I__9940 (
            .O(N__42709),
            .I(N__42654));
    CascadeMux I__9939 (
            .O(N__42708),
            .I(N__42649));
    InMux I__9938 (
            .O(N__42705),
            .I(N__42641));
    LocalMux I__9937 (
            .O(N__42702),
            .I(N__42638));
    InMux I__9936 (
            .O(N__42701),
            .I(N__42635));
    LocalMux I__9935 (
            .O(N__42698),
            .I(N__42624));
    LocalMux I__9934 (
            .O(N__42695),
            .I(N__42624));
    Span4Mux_s3_v I__9933 (
            .O(N__42692),
            .I(N__42624));
    Span4Mux_s3_v I__9932 (
            .O(N__42687),
            .I(N__42624));
    Span4Mux_v I__9931 (
            .O(N__42684),
            .I(N__42624));
    LocalMux I__9930 (
            .O(N__42681),
            .I(N__42619));
    InMux I__9929 (
            .O(N__42680),
            .I(N__42616));
    LocalMux I__9928 (
            .O(N__42675),
            .I(N__42611));
    Span4Mux_v I__9927 (
            .O(N__42670),
            .I(N__42611));
    LocalMux I__9926 (
            .O(N__42661),
            .I(N__42608));
    CascadeMux I__9925 (
            .O(N__42660),
            .I(N__42604));
    LocalMux I__9924 (
            .O(N__42657),
            .I(N__42598));
    LocalMux I__9923 (
            .O(N__42654),
            .I(N__42598));
    InMux I__9922 (
            .O(N__42653),
            .I(N__42593));
    InMux I__9921 (
            .O(N__42652),
            .I(N__42593));
    InMux I__9920 (
            .O(N__42649),
            .I(N__42589));
    InMux I__9919 (
            .O(N__42648),
            .I(N__42584));
    InMux I__9918 (
            .O(N__42647),
            .I(N__42584));
    InMux I__9917 (
            .O(N__42646),
            .I(N__42581));
    CascadeMux I__9916 (
            .O(N__42645),
            .I(N__42577));
    InMux I__9915 (
            .O(N__42644),
            .I(N__42571));
    LocalMux I__9914 (
            .O(N__42641),
            .I(N__42568));
    Span4Mux_h I__9913 (
            .O(N__42638),
            .I(N__42561));
    LocalMux I__9912 (
            .O(N__42635),
            .I(N__42561));
    Span4Mux_h I__9911 (
            .O(N__42624),
            .I(N__42561));
    CascadeMux I__9910 (
            .O(N__42623),
            .I(N__42558));
    CascadeMux I__9909 (
            .O(N__42622),
            .I(N__42555));
    Span4Mux_h I__9908 (
            .O(N__42619),
            .I(N__42546));
    LocalMux I__9907 (
            .O(N__42616),
            .I(N__42546));
    Span4Mux_s2_v I__9906 (
            .O(N__42611),
            .I(N__42546));
    Span4Mux_s2_v I__9905 (
            .O(N__42608),
            .I(N__42546));
    InMux I__9904 (
            .O(N__42607),
            .I(N__42543));
    InMux I__9903 (
            .O(N__42604),
            .I(N__42538));
    InMux I__9902 (
            .O(N__42603),
            .I(N__42538));
    Span4Mux_v I__9901 (
            .O(N__42598),
            .I(N__42533));
    LocalMux I__9900 (
            .O(N__42593),
            .I(N__42533));
    InMux I__9899 (
            .O(N__42592),
            .I(N__42530));
    LocalMux I__9898 (
            .O(N__42589),
            .I(N__42525));
    LocalMux I__9897 (
            .O(N__42584),
            .I(N__42525));
    LocalMux I__9896 (
            .O(N__42581),
            .I(N__42522));
    InMux I__9895 (
            .O(N__42580),
            .I(N__42515));
    InMux I__9894 (
            .O(N__42577),
            .I(N__42515));
    InMux I__9893 (
            .O(N__42576),
            .I(N__42515));
    InMux I__9892 (
            .O(N__42575),
            .I(N__42510));
    InMux I__9891 (
            .O(N__42574),
            .I(N__42510));
    LocalMux I__9890 (
            .O(N__42571),
            .I(N__42503));
    Span4Mux_h I__9889 (
            .O(N__42568),
            .I(N__42503));
    Span4Mux_h I__9888 (
            .O(N__42561),
            .I(N__42503));
    InMux I__9887 (
            .O(N__42558),
            .I(N__42498));
    InMux I__9886 (
            .O(N__42555),
            .I(N__42498));
    Span4Mux_h I__9885 (
            .O(N__42546),
            .I(N__42495));
    LocalMux I__9884 (
            .O(N__42543),
            .I(N__42484));
    LocalMux I__9883 (
            .O(N__42538),
            .I(N__42484));
    Sp12to4 I__9882 (
            .O(N__42533),
            .I(N__42484));
    LocalMux I__9881 (
            .O(N__42530),
            .I(N__42484));
    Span12Mux_v I__9880 (
            .O(N__42525),
            .I(N__42484));
    Odrv4 I__9879 (
            .O(N__42522),
            .I(UART_TRANSMITTER_state_2));
    LocalMux I__9878 (
            .O(N__42515),
            .I(UART_TRANSMITTER_state_2));
    LocalMux I__9877 (
            .O(N__42510),
            .I(UART_TRANSMITTER_state_2));
    Odrv4 I__9876 (
            .O(N__42503),
            .I(UART_TRANSMITTER_state_2));
    LocalMux I__9875 (
            .O(N__42498),
            .I(UART_TRANSMITTER_state_2));
    Odrv4 I__9874 (
            .O(N__42495),
            .I(UART_TRANSMITTER_state_2));
    Odrv12 I__9873 (
            .O(N__42484),
            .I(UART_TRANSMITTER_state_2));
    InMux I__9872 (
            .O(N__42469),
            .I(N__42461));
    InMux I__9871 (
            .O(N__42468),
            .I(N__42458));
    InMux I__9870 (
            .O(N__42467),
            .I(N__42455));
    InMux I__9869 (
            .O(N__42466),
            .I(N__42452));
    InMux I__9868 (
            .O(N__42465),
            .I(N__42449));
    InMux I__9867 (
            .O(N__42464),
            .I(N__42446));
    LocalMux I__9866 (
            .O(N__42461),
            .I(N__42443));
    LocalMux I__9865 (
            .O(N__42458),
            .I(N__42440));
    LocalMux I__9864 (
            .O(N__42455),
            .I(N__42436));
    LocalMux I__9863 (
            .O(N__42452),
            .I(N__42431));
    LocalMux I__9862 (
            .O(N__42449),
            .I(N__42431));
    LocalMux I__9861 (
            .O(N__42446),
            .I(N__42428));
    Span4Mux_v I__9860 (
            .O(N__42443),
            .I(N__42425));
    Span4Mux_h I__9859 (
            .O(N__42440),
            .I(N__42422));
    InMux I__9858 (
            .O(N__42439),
            .I(N__42419));
    Span4Mux_h I__9857 (
            .O(N__42436),
            .I(N__42414));
    Span4Mux_h I__9856 (
            .O(N__42431),
            .I(N__42414));
    Odrv12 I__9855 (
            .O(N__42428),
            .I(\c0.data_out_5_3 ));
    Odrv4 I__9854 (
            .O(N__42425),
            .I(\c0.data_out_5_3 ));
    Odrv4 I__9853 (
            .O(N__42422),
            .I(\c0.data_out_5_3 ));
    LocalMux I__9852 (
            .O(N__42419),
            .I(\c0.data_out_5_3 ));
    Odrv4 I__9851 (
            .O(N__42414),
            .I(\c0.data_out_5_3 ));
    InMux I__9850 (
            .O(N__42403),
            .I(N__42397));
    InMux I__9849 (
            .O(N__42402),
            .I(N__42393));
    InMux I__9848 (
            .O(N__42401),
            .I(N__42390));
    InMux I__9847 (
            .O(N__42400),
            .I(N__42387));
    LocalMux I__9846 (
            .O(N__42397),
            .I(N__42384));
    InMux I__9845 (
            .O(N__42396),
            .I(N__42380));
    LocalMux I__9844 (
            .O(N__42393),
            .I(N__42375));
    LocalMux I__9843 (
            .O(N__42390),
            .I(N__42375));
    LocalMux I__9842 (
            .O(N__42387),
            .I(N__42372));
    Span4Mux_v I__9841 (
            .O(N__42384),
            .I(N__42368));
    InMux I__9840 (
            .O(N__42383),
            .I(N__42365));
    LocalMux I__9839 (
            .O(N__42380),
            .I(N__42362));
    Span4Mux_v I__9838 (
            .O(N__42375),
            .I(N__42357));
    Span4Mux_v I__9837 (
            .O(N__42372),
            .I(N__42357));
    InMux I__9836 (
            .O(N__42371),
            .I(N__42354));
    Sp12to4 I__9835 (
            .O(N__42368),
            .I(N__42349));
    LocalMux I__9834 (
            .O(N__42365),
            .I(N__42349));
    Odrv12 I__9833 (
            .O(N__42362),
            .I(\c0.data_out_5_4 ));
    Odrv4 I__9832 (
            .O(N__42357),
            .I(\c0.data_out_5_4 ));
    LocalMux I__9831 (
            .O(N__42354),
            .I(\c0.data_out_5_4 ));
    Odrv12 I__9830 (
            .O(N__42349),
            .I(\c0.data_out_5_4 ));
    InMux I__9829 (
            .O(N__42340),
            .I(N__42337));
    LocalMux I__9828 (
            .O(N__42337),
            .I(N__42334));
    Odrv12 I__9827 (
            .O(N__42334),
            .I(\c0.n9783 ));
    InMux I__9826 (
            .O(N__42331),
            .I(N__42328));
    LocalMux I__9825 (
            .O(N__42328),
            .I(N__42323));
    InMux I__9824 (
            .O(N__42327),
            .I(N__42320));
    InMux I__9823 (
            .O(N__42326),
            .I(N__42317));
    Span4Mux_h I__9822 (
            .O(N__42323),
            .I(N__42310));
    LocalMux I__9821 (
            .O(N__42320),
            .I(N__42310));
    LocalMux I__9820 (
            .O(N__42317),
            .I(N__42307));
    InMux I__9819 (
            .O(N__42316),
            .I(N__42302));
    InMux I__9818 (
            .O(N__42315),
            .I(N__42302));
    Span4Mux_v I__9817 (
            .O(N__42310),
            .I(N__42299));
    Span4Mux_h I__9816 (
            .O(N__42307),
            .I(N__42296));
    LocalMux I__9815 (
            .O(N__42302),
            .I(data_out_frame2_10_6));
    Odrv4 I__9814 (
            .O(N__42299),
            .I(data_out_frame2_10_6));
    Odrv4 I__9813 (
            .O(N__42296),
            .I(data_out_frame2_10_6));
    InMux I__9812 (
            .O(N__42289),
            .I(N__42285));
    InMux I__9811 (
            .O(N__42288),
            .I(N__42281));
    LocalMux I__9810 (
            .O(N__42285),
            .I(N__42278));
    InMux I__9809 (
            .O(N__42284),
            .I(N__42275));
    LocalMux I__9808 (
            .O(N__42281),
            .I(N__42270));
    Span4Mux_h I__9807 (
            .O(N__42278),
            .I(N__42270));
    LocalMux I__9806 (
            .O(N__42275),
            .I(N__42267));
    Span4Mux_h I__9805 (
            .O(N__42270),
            .I(N__42264));
    Odrv4 I__9804 (
            .O(N__42267),
            .I(\c0.data_out_7_3 ));
    Odrv4 I__9803 (
            .O(N__42264),
            .I(\c0.data_out_7_3 ));
    InMux I__9802 (
            .O(N__42259),
            .I(N__42256));
    LocalMux I__9801 (
            .O(N__42256),
            .I(\c0.n8_adj_2153 ));
    InMux I__9800 (
            .O(N__42253),
            .I(N__42250));
    LocalMux I__9799 (
            .O(N__42250),
            .I(N__42246));
    InMux I__9798 (
            .O(N__42249),
            .I(N__42243));
    Odrv4 I__9797 (
            .O(N__42246),
            .I(\c0.n17070 ));
    LocalMux I__9796 (
            .O(N__42243),
            .I(\c0.n17070 ));
    CascadeMux I__9795 (
            .O(N__42238),
            .I(N__42235));
    InMux I__9794 (
            .O(N__42235),
            .I(N__42232));
    LocalMux I__9793 (
            .O(N__42232),
            .I(N__42229));
    Span4Mux_h I__9792 (
            .O(N__42229),
            .I(N__42225));
    InMux I__9791 (
            .O(N__42228),
            .I(N__42222));
    Odrv4 I__9790 (
            .O(N__42225),
            .I(\c0.n9737 ));
    LocalMux I__9789 (
            .O(N__42222),
            .I(\c0.n9737 ));
    CascadeMux I__9788 (
            .O(N__42217),
            .I(N__42214));
    InMux I__9787 (
            .O(N__42214),
            .I(N__42211));
    LocalMux I__9786 (
            .O(N__42211),
            .I(N__42208));
    Odrv4 I__9785 (
            .O(N__42208),
            .I(\c0.n12_adj_2285 ));
    InMux I__9784 (
            .O(N__42205),
            .I(N__42199));
    InMux I__9783 (
            .O(N__42204),
            .I(N__42194));
    InMux I__9782 (
            .O(N__42203),
            .I(N__42194));
    InMux I__9781 (
            .O(N__42202),
            .I(N__42191));
    LocalMux I__9780 (
            .O(N__42199),
            .I(N__42188));
    LocalMux I__9779 (
            .O(N__42194),
            .I(N__42185));
    LocalMux I__9778 (
            .O(N__42191),
            .I(N__42180));
    Span4Mux_v I__9777 (
            .O(N__42188),
            .I(N__42180));
    Span4Mux_h I__9776 (
            .O(N__42185),
            .I(N__42177));
    Odrv4 I__9775 (
            .O(N__42180),
            .I(\c0.data_out_6_3 ));
    Odrv4 I__9774 (
            .O(N__42177),
            .I(\c0.data_out_6_3 ));
    InMux I__9773 (
            .O(N__42172),
            .I(N__42166));
    InMux I__9772 (
            .O(N__42171),
            .I(N__42166));
    LocalMux I__9771 (
            .O(N__42166),
            .I(\c0.data_out_2_3 ));
    CascadeMux I__9770 (
            .O(N__42163),
            .I(N__42160));
    InMux I__9769 (
            .O(N__42160),
            .I(N__42157));
    LocalMux I__9768 (
            .O(N__42157),
            .I(N__42152));
    InMux I__9767 (
            .O(N__42156),
            .I(N__42149));
    CascadeMux I__9766 (
            .O(N__42155),
            .I(N__42146));
    Span4Mux_v I__9765 (
            .O(N__42152),
            .I(N__42141));
    LocalMux I__9764 (
            .O(N__42149),
            .I(N__42141));
    InMux I__9763 (
            .O(N__42146),
            .I(N__42138));
    Span4Mux_h I__9762 (
            .O(N__42141),
            .I(N__42135));
    LocalMux I__9761 (
            .O(N__42138),
            .I(N__42132));
    Span4Mux_v I__9760 (
            .O(N__42135),
            .I(N__42126));
    Span4Mux_v I__9759 (
            .O(N__42132),
            .I(N__42126));
    InMux I__9758 (
            .O(N__42131),
            .I(N__42123));
    Odrv4 I__9757 (
            .O(N__42126),
            .I(n2652));
    LocalMux I__9756 (
            .O(N__42123),
            .I(n2652));
    InMux I__9755 (
            .O(N__42118),
            .I(N__42115));
    LocalMux I__9754 (
            .O(N__42115),
            .I(\c0.n5_adj_2350 ));
    CascadeMux I__9753 (
            .O(N__42112),
            .I(\c0.n17546_cascade_ ));
    InMux I__9752 (
            .O(N__42109),
            .I(N__42106));
    LocalMux I__9751 (
            .O(N__42106),
            .I(N__42103));
    Span4Mux_v I__9750 (
            .O(N__42103),
            .I(N__42100));
    Span4Mux_h I__9749 (
            .O(N__42100),
            .I(N__42097));
    Odrv4 I__9748 (
            .O(N__42097),
            .I(\c0.n17592 ));
    CascadeMux I__9747 (
            .O(N__42094),
            .I(\c0.n18059_cascade_ ));
    InMux I__9746 (
            .O(N__42091),
            .I(N__42088));
    LocalMux I__9745 (
            .O(N__42088),
            .I(N__42085));
    Span4Mux_v I__9744 (
            .O(N__42085),
            .I(N__42082));
    Span4Mux_h I__9743 (
            .O(N__42082),
            .I(N__42079));
    Odrv4 I__9742 (
            .O(N__42079),
            .I(\c0.data_out_frame2_20_7 ));
    CascadeMux I__9741 (
            .O(N__42076),
            .I(\c0.n18062_cascade_ ));
    InMux I__9740 (
            .O(N__42073),
            .I(N__42069));
    InMux I__9739 (
            .O(N__42072),
            .I(N__42063));
    LocalMux I__9738 (
            .O(N__42069),
            .I(N__42060));
    InMux I__9737 (
            .O(N__42068),
            .I(N__42057));
    InMux I__9736 (
            .O(N__42067),
            .I(N__42054));
    InMux I__9735 (
            .O(N__42066),
            .I(N__42051));
    LocalMux I__9734 (
            .O(N__42063),
            .I(N__42048));
    Span4Mux_h I__9733 (
            .O(N__42060),
            .I(N__42043));
    LocalMux I__9732 (
            .O(N__42057),
            .I(N__42043));
    LocalMux I__9731 (
            .O(N__42054),
            .I(data_out_frame2_11_4));
    LocalMux I__9730 (
            .O(N__42051),
            .I(data_out_frame2_11_4));
    Odrv12 I__9729 (
            .O(N__42048),
            .I(data_out_frame2_11_4));
    Odrv4 I__9728 (
            .O(N__42043),
            .I(data_out_frame2_11_4));
    InMux I__9727 (
            .O(N__42034),
            .I(N__42028));
    InMux I__9726 (
            .O(N__42033),
            .I(N__42028));
    LocalMux I__9725 (
            .O(N__42028),
            .I(data_out_frame2_17_7));
    InMux I__9724 (
            .O(N__42025),
            .I(N__42020));
    InMux I__9723 (
            .O(N__42024),
            .I(N__42015));
    InMux I__9722 (
            .O(N__42023),
            .I(N__42015));
    LocalMux I__9721 (
            .O(N__42020),
            .I(data_out_frame2_14_0));
    LocalMux I__9720 (
            .O(N__42015),
            .I(data_out_frame2_14_0));
    CascadeMux I__9719 (
            .O(N__42010),
            .I(N__42007));
    InMux I__9718 (
            .O(N__42007),
            .I(N__42004));
    LocalMux I__9717 (
            .O(N__42004),
            .I(N__42001));
    Span12Mux_v I__9716 (
            .O(N__42001),
            .I(N__41998));
    Odrv12 I__9715 (
            .O(N__41998),
            .I(\c0.n9853 ));
    CascadeMux I__9714 (
            .O(N__41995),
            .I(N__41991));
    InMux I__9713 (
            .O(N__41994),
            .I(N__41988));
    InMux I__9712 (
            .O(N__41991),
            .I(N__41985));
    LocalMux I__9711 (
            .O(N__41988),
            .I(N__41982));
    LocalMux I__9710 (
            .O(N__41985),
            .I(N__41979));
    Span4Mux_v I__9709 (
            .O(N__41982),
            .I(N__41974));
    Span4Mux_v I__9708 (
            .O(N__41979),
            .I(N__41974));
    Odrv4 I__9707 (
            .O(N__41974),
            .I(\c0.n9589 ));
    CascadeMux I__9706 (
            .O(N__41971),
            .I(\c0.n9853_cascade_ ));
    CascadeMux I__9705 (
            .O(N__41968),
            .I(N__41965));
    InMux I__9704 (
            .O(N__41965),
            .I(N__41962));
    LocalMux I__9703 (
            .O(N__41962),
            .I(N__41959));
    Span12Mux_v I__9702 (
            .O(N__41959),
            .I(N__41953));
    InMux I__9701 (
            .O(N__41958),
            .I(N__41950));
    InMux I__9700 (
            .O(N__41957),
            .I(N__41945));
    InMux I__9699 (
            .O(N__41956),
            .I(N__41945));
    Odrv12 I__9698 (
            .O(N__41953),
            .I(data_out_frame2_13_0));
    LocalMux I__9697 (
            .O(N__41950),
            .I(data_out_frame2_13_0));
    LocalMux I__9696 (
            .O(N__41945),
            .I(data_out_frame2_13_0));
    InMux I__9695 (
            .O(N__41938),
            .I(N__41935));
    LocalMux I__9694 (
            .O(N__41935),
            .I(N__41931));
    InMux I__9693 (
            .O(N__41934),
            .I(N__41928));
    Span4Mux_v I__9692 (
            .O(N__41931),
            .I(N__41923));
    LocalMux I__9691 (
            .O(N__41928),
            .I(N__41923));
    Span4Mux_h I__9690 (
            .O(N__41923),
            .I(N__41920));
    Span4Mux_v I__9689 (
            .O(N__41920),
            .I(N__41917));
    Span4Mux_h I__9688 (
            .O(N__41917),
            .I(N__41914));
    Odrv4 I__9687 (
            .O(N__41914),
            .I(\c0.n17046 ));
    InMux I__9686 (
            .O(N__41911),
            .I(N__41908));
    LocalMux I__9685 (
            .O(N__41908),
            .I(N__41905));
    Span4Mux_h I__9684 (
            .O(N__41905),
            .I(N__41902));
    Span4Mux_h I__9683 (
            .O(N__41902),
            .I(N__41899));
    Odrv4 I__9682 (
            .O(N__41899),
            .I(\c0.n17581 ));
    SRMux I__9681 (
            .O(N__41896),
            .I(N__41893));
    LocalMux I__9680 (
            .O(N__41893),
            .I(N__41890));
    Span4Mux_h I__9679 (
            .O(N__41890),
            .I(N__41886));
    SRMux I__9678 (
            .O(N__41889),
            .I(N__41883));
    Span4Mux_s0_v I__9677 (
            .O(N__41886),
            .I(N__41878));
    LocalMux I__9676 (
            .O(N__41883),
            .I(N__41878));
    Span4Mux_v I__9675 (
            .O(N__41878),
            .I(N__41875));
    Odrv4 I__9674 (
            .O(N__41875),
            .I(\c0.n10259 ));
    InMux I__9673 (
            .O(N__41872),
            .I(N__41869));
    LocalMux I__9672 (
            .O(N__41869),
            .I(N__41863));
    InMux I__9671 (
            .O(N__41868),
            .I(N__41860));
    InMux I__9670 (
            .O(N__41867),
            .I(N__41856));
    InMux I__9669 (
            .O(N__41866),
            .I(N__41853));
    Span4Mux_h I__9668 (
            .O(N__41863),
            .I(N__41850));
    LocalMux I__9667 (
            .O(N__41860),
            .I(N__41847));
    InMux I__9666 (
            .O(N__41859),
            .I(N__41844));
    LocalMux I__9665 (
            .O(N__41856),
            .I(data_out_frame2_8_5));
    LocalMux I__9664 (
            .O(N__41853),
            .I(data_out_frame2_8_5));
    Odrv4 I__9663 (
            .O(N__41850),
            .I(data_out_frame2_8_5));
    Odrv12 I__9662 (
            .O(N__41847),
            .I(data_out_frame2_8_5));
    LocalMux I__9661 (
            .O(N__41844),
            .I(data_out_frame2_8_5));
    InMux I__9660 (
            .O(N__41833),
            .I(N__41828));
    InMux I__9659 (
            .O(N__41832),
            .I(N__41825));
    InMux I__9658 (
            .O(N__41831),
            .I(N__41822));
    LocalMux I__9657 (
            .O(N__41828),
            .I(N__41819));
    LocalMux I__9656 (
            .O(N__41825),
            .I(N__41816));
    LocalMux I__9655 (
            .O(N__41822),
            .I(N__41812));
    Span4Mux_v I__9654 (
            .O(N__41819),
            .I(N__41809));
    Span4Mux_h I__9653 (
            .O(N__41816),
            .I(N__41806));
    InMux I__9652 (
            .O(N__41815),
            .I(N__41803));
    Span4Mux_h I__9651 (
            .O(N__41812),
            .I(N__41800));
    Span4Mux_h I__9650 (
            .O(N__41809),
            .I(N__41795));
    Span4Mux_v I__9649 (
            .O(N__41806),
            .I(N__41795));
    LocalMux I__9648 (
            .O(N__41803),
            .I(data_out_frame2_10_3));
    Odrv4 I__9647 (
            .O(N__41800),
            .I(data_out_frame2_10_3));
    Odrv4 I__9646 (
            .O(N__41795),
            .I(data_out_frame2_10_3));
    InMux I__9645 (
            .O(N__41788),
            .I(N__41785));
    LocalMux I__9644 (
            .O(N__41785),
            .I(N__41782));
    Span4Mux_h I__9643 (
            .O(N__41782),
            .I(N__41779));
    Span4Mux_v I__9642 (
            .O(N__41779),
            .I(N__41776));
    Odrv4 I__9641 (
            .O(N__41776),
            .I(\c0.n20_adj_2252 ));
    InMux I__9640 (
            .O(N__41773),
            .I(N__41770));
    LocalMux I__9639 (
            .O(N__41770),
            .I(\c0.n17322 ));
    CascadeMux I__9638 (
            .O(N__41767),
            .I(\c0.n17323_cascade_ ));
    CascadeMux I__9637 (
            .O(N__41764),
            .I(N__41761));
    InMux I__9636 (
            .O(N__41761),
            .I(N__41758));
    LocalMux I__9635 (
            .O(N__41758),
            .I(\c0.n18053 ));
    InMux I__9634 (
            .O(N__41755),
            .I(N__41749));
    InMux I__9633 (
            .O(N__41754),
            .I(N__41746));
    InMux I__9632 (
            .O(N__41753),
            .I(N__41743));
    InMux I__9631 (
            .O(N__41752),
            .I(N__41740));
    LocalMux I__9630 (
            .O(N__41749),
            .I(N__41737));
    LocalMux I__9629 (
            .O(N__41746),
            .I(N__41734));
    LocalMux I__9628 (
            .O(N__41743),
            .I(N__41730));
    LocalMux I__9627 (
            .O(N__41740),
            .I(N__41727));
    Span4Mux_v I__9626 (
            .O(N__41737),
            .I(N__41724));
    Span4Mux_v I__9625 (
            .O(N__41734),
            .I(N__41721));
    InMux I__9624 (
            .O(N__41733),
            .I(N__41718));
    Span4Mux_v I__9623 (
            .O(N__41730),
            .I(N__41713));
    Span4Mux_s3_v I__9622 (
            .O(N__41727),
            .I(N__41713));
    Odrv4 I__9621 (
            .O(N__41724),
            .I(rand_data_16));
    Odrv4 I__9620 (
            .O(N__41721),
            .I(rand_data_16));
    LocalMux I__9619 (
            .O(N__41718),
            .I(rand_data_16));
    Odrv4 I__9618 (
            .O(N__41713),
            .I(rand_data_16));
    InMux I__9617 (
            .O(N__41704),
            .I(N__41700));
    InMux I__9616 (
            .O(N__41703),
            .I(N__41697));
    LocalMux I__9615 (
            .O(N__41700),
            .I(N__41691));
    LocalMux I__9614 (
            .O(N__41697),
            .I(N__41691));
    InMux I__9613 (
            .O(N__41696),
            .I(N__41686));
    Span12Mux_h I__9612 (
            .O(N__41691),
            .I(N__41683));
    InMux I__9611 (
            .O(N__41690),
            .I(N__41680));
    InMux I__9610 (
            .O(N__41689),
            .I(N__41677));
    LocalMux I__9609 (
            .O(N__41686),
            .I(data_out_frame2_9_1));
    Odrv12 I__9608 (
            .O(N__41683),
            .I(data_out_frame2_9_1));
    LocalMux I__9607 (
            .O(N__41680),
            .I(data_out_frame2_9_1));
    LocalMux I__9606 (
            .O(N__41677),
            .I(data_out_frame2_9_1));
    InMux I__9605 (
            .O(N__41668),
            .I(N__41665));
    LocalMux I__9604 (
            .O(N__41665),
            .I(\c0.n17921 ));
    InMux I__9603 (
            .O(N__41662),
            .I(N__41659));
    LocalMux I__9602 (
            .O(N__41659),
            .I(N__41656));
    Span4Mux_h I__9601 (
            .O(N__41656),
            .I(N__41653));
    Span4Mux_h I__9600 (
            .O(N__41653),
            .I(N__41650));
    Odrv4 I__9599 (
            .O(N__41650),
            .I(\c0.n17924 ));
    InMux I__9598 (
            .O(N__41647),
            .I(N__41641));
    InMux I__9597 (
            .O(N__41646),
            .I(N__41641));
    LocalMux I__9596 (
            .O(N__41641),
            .I(data_out_frame2_18_7));
    CascadeMux I__9595 (
            .O(N__41638),
            .I(N__41635));
    InMux I__9594 (
            .O(N__41635),
            .I(N__41632));
    LocalMux I__9593 (
            .O(N__41632),
            .I(N__41629));
    Span4Mux_v I__9592 (
            .O(N__41629),
            .I(N__41626));
    Odrv4 I__9591 (
            .O(N__41626),
            .I(\c0.data_out_frame2_19_7 ));
    CascadeMux I__9590 (
            .O(N__41623),
            .I(N__41620));
    InMux I__9589 (
            .O(N__41620),
            .I(N__41617));
    LocalMux I__9588 (
            .O(N__41617),
            .I(N__41614));
    Odrv4 I__9587 (
            .O(N__41614),
            .I(\c0.n17034 ));
    CascadeMux I__9586 (
            .O(N__41611),
            .I(\c0.n17034_cascade_ ));
    InMux I__9585 (
            .O(N__41608),
            .I(N__41605));
    LocalMux I__9584 (
            .O(N__41605),
            .I(N__41602));
    Span4Mux_h I__9583 (
            .O(N__41602),
            .I(N__41599));
    Odrv4 I__9582 (
            .O(N__41599),
            .I(\c0.n9688 ));
    InMux I__9581 (
            .O(N__41596),
            .I(N__41591));
    InMux I__9580 (
            .O(N__41595),
            .I(N__41588));
    InMux I__9579 (
            .O(N__41594),
            .I(N__41585));
    LocalMux I__9578 (
            .O(N__41591),
            .I(N__41582));
    LocalMux I__9577 (
            .O(N__41588),
            .I(N__41579));
    LocalMux I__9576 (
            .O(N__41585),
            .I(N__41576));
    Span4Mux_v I__9575 (
            .O(N__41582),
            .I(N__41571));
    Span4Mux_v I__9574 (
            .O(N__41579),
            .I(N__41571));
    Span4Mux_v I__9573 (
            .O(N__41576),
            .I(N__41566));
    Span4Mux_h I__9572 (
            .O(N__41571),
            .I(N__41563));
    InMux I__9571 (
            .O(N__41570),
            .I(N__41558));
    InMux I__9570 (
            .O(N__41569),
            .I(N__41558));
    Odrv4 I__9569 (
            .O(N__41566),
            .I(data_out_frame2_12_1));
    Odrv4 I__9568 (
            .O(N__41563),
            .I(data_out_frame2_12_1));
    LocalMux I__9567 (
            .O(N__41558),
            .I(data_out_frame2_12_1));
    CascadeMux I__9566 (
            .O(N__41551),
            .I(\c0.n9688_cascade_ ));
    InMux I__9565 (
            .O(N__41548),
            .I(N__41545));
    LocalMux I__9564 (
            .O(N__41545),
            .I(\c0.n6_adj_2325 ));
    InMux I__9563 (
            .O(N__41542),
            .I(N__41539));
    LocalMux I__9562 (
            .O(N__41539),
            .I(N__41536));
    Span4Mux_h I__9561 (
            .O(N__41536),
            .I(N__41531));
    InMux I__9560 (
            .O(N__41535),
            .I(N__41526));
    InMux I__9559 (
            .O(N__41534),
            .I(N__41526));
    Odrv4 I__9558 (
            .O(N__41531),
            .I(data_out_frame2_11_1));
    LocalMux I__9557 (
            .O(N__41526),
            .I(data_out_frame2_11_1));
    InMux I__9556 (
            .O(N__41521),
            .I(N__41518));
    LocalMux I__9555 (
            .O(N__41518),
            .I(N__41515));
    Span4Mux_h I__9554 (
            .O(N__41515),
            .I(N__41510));
    InMux I__9553 (
            .O(N__41514),
            .I(N__41506));
    InMux I__9552 (
            .O(N__41513),
            .I(N__41503));
    Span4Mux_h I__9551 (
            .O(N__41510),
            .I(N__41500));
    InMux I__9550 (
            .O(N__41509),
            .I(N__41497));
    LocalMux I__9549 (
            .O(N__41506),
            .I(data_out_frame2_6_1));
    LocalMux I__9548 (
            .O(N__41503),
            .I(data_out_frame2_6_1));
    Odrv4 I__9547 (
            .O(N__41500),
            .I(data_out_frame2_6_1));
    LocalMux I__9546 (
            .O(N__41497),
            .I(data_out_frame2_6_1));
    InMux I__9545 (
            .O(N__41488),
            .I(N__41484));
    InMux I__9544 (
            .O(N__41487),
            .I(N__41481));
    LocalMux I__9543 (
            .O(N__41484),
            .I(N__41476));
    LocalMux I__9542 (
            .O(N__41481),
            .I(N__41476));
    Sp12to4 I__9541 (
            .O(N__41476),
            .I(N__41473));
    Odrv12 I__9540 (
            .O(N__41473),
            .I(\c0.n17115 ));
    InMux I__9539 (
            .O(N__41470),
            .I(N__41466));
    InMux I__9538 (
            .O(N__41469),
            .I(N__41461));
    LocalMux I__9537 (
            .O(N__41466),
            .I(N__41458));
    InMux I__9536 (
            .O(N__41465),
            .I(N__41455));
    InMux I__9535 (
            .O(N__41464),
            .I(N__41451));
    LocalMux I__9534 (
            .O(N__41461),
            .I(N__41448));
    Span4Mux_h I__9533 (
            .O(N__41458),
            .I(N__41445));
    LocalMux I__9532 (
            .O(N__41455),
            .I(N__41441));
    InMux I__9531 (
            .O(N__41454),
            .I(N__41438));
    LocalMux I__9530 (
            .O(N__41451),
            .I(N__41433));
    Span12Mux_v I__9529 (
            .O(N__41448),
            .I(N__41433));
    Span4Mux_v I__9528 (
            .O(N__41445),
            .I(N__41430));
    InMux I__9527 (
            .O(N__41444),
            .I(N__41427));
    Span4Mux_v I__9526 (
            .O(N__41441),
            .I(N__41424));
    LocalMux I__9525 (
            .O(N__41438),
            .I(rand_data_5));
    Odrv12 I__9524 (
            .O(N__41433),
            .I(rand_data_5));
    Odrv4 I__9523 (
            .O(N__41430),
            .I(rand_data_5));
    LocalMux I__9522 (
            .O(N__41427),
            .I(rand_data_5));
    Odrv4 I__9521 (
            .O(N__41424),
            .I(rand_data_5));
    CascadeMux I__9520 (
            .O(N__41413),
            .I(N__41410));
    InMux I__9519 (
            .O(N__41410),
            .I(N__41407));
    LocalMux I__9518 (
            .O(N__41407),
            .I(N__41403));
    InMux I__9517 (
            .O(N__41406),
            .I(N__41400));
    Span4Mux_h I__9516 (
            .O(N__41403),
            .I(N__41395));
    LocalMux I__9515 (
            .O(N__41400),
            .I(N__41392));
    InMux I__9514 (
            .O(N__41399),
            .I(N__41387));
    InMux I__9513 (
            .O(N__41398),
            .I(N__41387));
    Odrv4 I__9512 (
            .O(N__41395),
            .I(data_out_frame2_16_5));
    Odrv12 I__9511 (
            .O(N__41392),
            .I(data_out_frame2_16_5));
    LocalMux I__9510 (
            .O(N__41387),
            .I(data_out_frame2_16_5));
    InMux I__9509 (
            .O(N__41380),
            .I(N__41376));
    InMux I__9508 (
            .O(N__41379),
            .I(N__41373));
    LocalMux I__9507 (
            .O(N__41376),
            .I(N__41370));
    LocalMux I__9506 (
            .O(N__41373),
            .I(N__41367));
    Span4Mux_v I__9505 (
            .O(N__41370),
            .I(N__41364));
    Odrv12 I__9504 (
            .O(N__41367),
            .I(\c0.n17040 ));
    Odrv4 I__9503 (
            .O(N__41364),
            .I(\c0.n17040 ));
    InMux I__9502 (
            .O(N__41359),
            .I(N__41356));
    LocalMux I__9501 (
            .O(N__41356),
            .I(\c0.n16972 ));
    InMux I__9500 (
            .O(N__41353),
            .I(N__41350));
    LocalMux I__9499 (
            .O(N__41350),
            .I(\c0.n30_adj_2295 ));
    InMux I__9498 (
            .O(N__41347),
            .I(N__41340));
    InMux I__9497 (
            .O(N__41346),
            .I(N__41337));
    InMux I__9496 (
            .O(N__41345),
            .I(N__41334));
    InMux I__9495 (
            .O(N__41344),
            .I(N__41331));
    InMux I__9494 (
            .O(N__41343),
            .I(N__41328));
    LocalMux I__9493 (
            .O(N__41340),
            .I(N__41325));
    LocalMux I__9492 (
            .O(N__41337),
            .I(N__41322));
    LocalMux I__9491 (
            .O(N__41334),
            .I(N__41319));
    LocalMux I__9490 (
            .O(N__41331),
            .I(N__41313));
    LocalMux I__9489 (
            .O(N__41328),
            .I(N__41313));
    Span4Mux_v I__9488 (
            .O(N__41325),
            .I(N__41308));
    Span4Mux_v I__9487 (
            .O(N__41322),
            .I(N__41308));
    Span4Mux_v I__9486 (
            .O(N__41319),
            .I(N__41305));
    InMux I__9485 (
            .O(N__41318),
            .I(N__41302));
    Span4Mux_v I__9484 (
            .O(N__41313),
            .I(N__41297));
    Span4Mux_h I__9483 (
            .O(N__41308),
            .I(N__41297));
    Span4Mux_h I__9482 (
            .O(N__41305),
            .I(N__41294));
    LocalMux I__9481 (
            .O(N__41302),
            .I(data_out_frame2_7_7));
    Odrv4 I__9480 (
            .O(N__41297),
            .I(data_out_frame2_7_7));
    Odrv4 I__9479 (
            .O(N__41294),
            .I(data_out_frame2_7_7));
    CascadeMux I__9478 (
            .O(N__41287),
            .I(N__41284));
    InMux I__9477 (
            .O(N__41284),
            .I(N__41281));
    LocalMux I__9476 (
            .O(N__41281),
            .I(N__41278));
    Span4Mux_h I__9475 (
            .O(N__41278),
            .I(N__41275));
    Span4Mux_h I__9474 (
            .O(N__41275),
            .I(N__41272));
    Odrv4 I__9473 (
            .O(N__41272),
            .I(\c0.n5_adj_2351 ));
    CascadeMux I__9472 (
            .O(N__41269),
            .I(N__41265));
    InMux I__9471 (
            .O(N__41268),
            .I(N__41260));
    InMux I__9470 (
            .O(N__41265),
            .I(N__41255));
    InMux I__9469 (
            .O(N__41264),
            .I(N__41255));
    InMux I__9468 (
            .O(N__41263),
            .I(N__41252));
    LocalMux I__9467 (
            .O(N__41260),
            .I(N__41249));
    LocalMux I__9466 (
            .O(N__41255),
            .I(data_out_frame2_11_3));
    LocalMux I__9465 (
            .O(N__41252),
            .I(data_out_frame2_11_3));
    Odrv4 I__9464 (
            .O(N__41249),
            .I(data_out_frame2_11_3));
    InMux I__9463 (
            .O(N__41242),
            .I(N__41239));
    LocalMux I__9462 (
            .O(N__41239),
            .I(N__41235));
    InMux I__9461 (
            .O(N__41238),
            .I(N__41232));
    Span4Mux_h I__9460 (
            .O(N__41235),
            .I(N__41229));
    LocalMux I__9459 (
            .O(N__41232),
            .I(N__41226));
    Odrv4 I__9458 (
            .O(N__41229),
            .I(\c0.n9695 ));
    Odrv12 I__9457 (
            .O(N__41226),
            .I(\c0.n9695 ));
    CascadeMux I__9456 (
            .O(N__41221),
            .I(\c0.n9695_cascade_ ));
    InMux I__9455 (
            .O(N__41218),
            .I(N__41214));
    CascadeMux I__9454 (
            .O(N__41217),
            .I(N__41211));
    LocalMux I__9453 (
            .O(N__41214),
            .I(N__41208));
    InMux I__9452 (
            .O(N__41211),
            .I(N__41205));
    Span4Mux_h I__9451 (
            .O(N__41208),
            .I(N__41198));
    LocalMux I__9450 (
            .O(N__41205),
            .I(N__41198));
    InMux I__9449 (
            .O(N__41204),
            .I(N__41195));
    InMux I__9448 (
            .O(N__41203),
            .I(N__41192));
    Span4Mux_h I__9447 (
            .O(N__41198),
            .I(N__41189));
    LocalMux I__9446 (
            .O(N__41195),
            .I(N__41186));
    LocalMux I__9445 (
            .O(N__41192),
            .I(N__41182));
    Span4Mux_v I__9444 (
            .O(N__41189),
            .I(N__41179));
    Span4Mux_v I__9443 (
            .O(N__41186),
            .I(N__41176));
    InMux I__9442 (
            .O(N__41185),
            .I(N__41173));
    Span4Mux_s2_v I__9441 (
            .O(N__41182),
            .I(N__41170));
    Odrv4 I__9440 (
            .O(N__41179),
            .I(rand_data_22));
    Odrv4 I__9439 (
            .O(N__41176),
            .I(rand_data_22));
    LocalMux I__9438 (
            .O(N__41173),
            .I(rand_data_22));
    Odrv4 I__9437 (
            .O(N__41170),
            .I(rand_data_22));
    InMux I__9436 (
            .O(N__41161),
            .I(N__41155));
    InMux I__9435 (
            .O(N__41160),
            .I(N__41150));
    InMux I__9434 (
            .O(N__41159),
            .I(N__41150));
    InMux I__9433 (
            .O(N__41158),
            .I(N__41147));
    LocalMux I__9432 (
            .O(N__41155),
            .I(data_out_frame2_11_7));
    LocalMux I__9431 (
            .O(N__41150),
            .I(data_out_frame2_11_7));
    LocalMux I__9430 (
            .O(N__41147),
            .I(data_out_frame2_11_7));
    InMux I__9429 (
            .O(N__41140),
            .I(N__41137));
    LocalMux I__9428 (
            .O(N__41137),
            .I(N__41132));
    InMux I__9427 (
            .O(N__41136),
            .I(N__41128));
    InMux I__9426 (
            .O(N__41135),
            .I(N__41125));
    Span4Mux_h I__9425 (
            .O(N__41132),
            .I(N__41122));
    InMux I__9424 (
            .O(N__41131),
            .I(N__41119));
    LocalMux I__9423 (
            .O(N__41128),
            .I(data_out_frame2_11_5));
    LocalMux I__9422 (
            .O(N__41125),
            .I(data_out_frame2_11_5));
    Odrv4 I__9421 (
            .O(N__41122),
            .I(data_out_frame2_11_5));
    LocalMux I__9420 (
            .O(N__41119),
            .I(data_out_frame2_11_5));
    InMux I__9419 (
            .O(N__41110),
            .I(N__41106));
    InMux I__9418 (
            .O(N__41109),
            .I(N__41103));
    LocalMux I__9417 (
            .O(N__41106),
            .I(N__41100));
    LocalMux I__9416 (
            .O(N__41103),
            .I(N__41097));
    Span4Mux_v I__9415 (
            .O(N__41100),
            .I(N__41094));
    Span12Mux_s11_v I__9414 (
            .O(N__41097),
            .I(N__41091));
    Odrv4 I__9413 (
            .O(N__41094),
            .I(\c0.n9919 ));
    Odrv12 I__9412 (
            .O(N__41091),
            .I(\c0.n9919 ));
    InMux I__9411 (
            .O(N__41086),
            .I(N__41083));
    LocalMux I__9410 (
            .O(N__41083),
            .I(N__41080));
    Span4Mux_h I__9409 (
            .O(N__41080),
            .I(N__41077));
    Odrv4 I__9408 (
            .O(N__41077),
            .I(\c0.n9901 ));
    InMux I__9407 (
            .O(N__41074),
            .I(N__41071));
    LocalMux I__9406 (
            .O(N__41071),
            .I(\c0.n10_adj_2292 ));
    InMux I__9405 (
            .O(N__41068),
            .I(N__41064));
    CascadeMux I__9404 (
            .O(N__41067),
            .I(N__41061));
    LocalMux I__9403 (
            .O(N__41064),
            .I(N__41058));
    InMux I__9402 (
            .O(N__41061),
            .I(N__41055));
    Span4Mux_v I__9401 (
            .O(N__41058),
            .I(N__41050));
    LocalMux I__9400 (
            .O(N__41055),
            .I(N__41050));
    Span4Mux_v I__9399 (
            .O(N__41050),
            .I(N__41046));
    InMux I__9398 (
            .O(N__41049),
            .I(N__41043));
    Span4Mux_h I__9397 (
            .O(N__41046),
            .I(N__41037));
    LocalMux I__9396 (
            .O(N__41043),
            .I(N__41034));
    InMux I__9395 (
            .O(N__41042),
            .I(N__41031));
    InMux I__9394 (
            .O(N__41041),
            .I(N__41026));
    InMux I__9393 (
            .O(N__41040),
            .I(N__41026));
    Odrv4 I__9392 (
            .O(N__41037),
            .I(data_out_frame2_7_4));
    Odrv4 I__9391 (
            .O(N__41034),
            .I(data_out_frame2_7_4));
    LocalMux I__9390 (
            .O(N__41031),
            .I(data_out_frame2_7_4));
    LocalMux I__9389 (
            .O(N__41026),
            .I(data_out_frame2_7_4));
    InMux I__9388 (
            .O(N__41017),
            .I(N__41014));
    LocalMux I__9387 (
            .O(N__41014),
            .I(N__41011));
    Span4Mux_h I__9386 (
            .O(N__41011),
            .I(N__41008));
    Odrv4 I__9385 (
            .O(N__41008),
            .I(\c0.n9913 ));
    InMux I__9384 (
            .O(N__41005),
            .I(N__41002));
    LocalMux I__9383 (
            .O(N__41002),
            .I(\c0.n29_adj_2296 ));
    InMux I__9382 (
            .O(N__40999),
            .I(N__40996));
    LocalMux I__9381 (
            .O(N__40996),
            .I(N__40993));
    Span4Mux_v I__9380 (
            .O(N__40993),
            .I(N__40990));
    Odrv4 I__9379 (
            .O(N__40990),
            .I(\c0.n16933 ));
    CascadeMux I__9378 (
            .O(N__40987),
            .I(\c0.n16915_cascade_ ));
    InMux I__9377 (
            .O(N__40984),
            .I(N__40980));
    InMux I__9376 (
            .O(N__40983),
            .I(N__40974));
    LocalMux I__9375 (
            .O(N__40980),
            .I(N__40971));
    InMux I__9374 (
            .O(N__40979),
            .I(N__40968));
    InMux I__9373 (
            .O(N__40978),
            .I(N__40965));
    InMux I__9372 (
            .O(N__40977),
            .I(N__40962));
    LocalMux I__9371 (
            .O(N__40974),
            .I(N__40957));
    Span4Mux_h I__9370 (
            .O(N__40971),
            .I(N__40957));
    LocalMux I__9369 (
            .O(N__40968),
            .I(N__40954));
    LocalMux I__9368 (
            .O(N__40965),
            .I(N__40949));
    LocalMux I__9367 (
            .O(N__40962),
            .I(N__40949));
    Odrv4 I__9366 (
            .O(N__40957),
            .I(data_out_frame2_7_2));
    Odrv4 I__9365 (
            .O(N__40954),
            .I(data_out_frame2_7_2));
    Odrv12 I__9364 (
            .O(N__40949),
            .I(data_out_frame2_7_2));
    InMux I__9363 (
            .O(N__40942),
            .I(N__40939));
    LocalMux I__9362 (
            .O(N__40939),
            .I(\c0.n19_adj_2303 ));
    CascadeMux I__9361 (
            .O(N__40936),
            .I(\c0.n20_adj_2302_cascade_ ));
    InMux I__9360 (
            .O(N__40933),
            .I(N__40930));
    LocalMux I__9359 (
            .O(N__40930),
            .I(N__40927));
    Odrv4 I__9358 (
            .O(N__40927),
            .I(\c0.n21_adj_2304 ));
    CascadeMux I__9357 (
            .O(N__40924),
            .I(N__40921));
    InMux I__9356 (
            .O(N__40921),
            .I(N__40918));
    LocalMux I__9355 (
            .O(N__40918),
            .I(N__40915));
    Odrv4 I__9354 (
            .O(N__40915),
            .I(\c0.data_out_frame2_19_6 ));
    InMux I__9353 (
            .O(N__40912),
            .I(N__40909));
    LocalMux I__9352 (
            .O(N__40909),
            .I(N__40906));
    Span4Mux_v I__9351 (
            .O(N__40906),
            .I(N__40901));
    InMux I__9350 (
            .O(N__40905),
            .I(N__40895));
    InMux I__9349 (
            .O(N__40904),
            .I(N__40895));
    Span4Mux_h I__9348 (
            .O(N__40901),
            .I(N__40892));
    InMux I__9347 (
            .O(N__40900),
            .I(N__40889));
    LocalMux I__9346 (
            .O(N__40895),
            .I(N__40886));
    Odrv4 I__9345 (
            .O(N__40892),
            .I(\c0.data_out_frame2_0_0 ));
    LocalMux I__9344 (
            .O(N__40889),
            .I(\c0.data_out_frame2_0_0 ));
    Odrv12 I__9343 (
            .O(N__40886),
            .I(\c0.data_out_frame2_0_0 ));
    CascadeMux I__9342 (
            .O(N__40879),
            .I(\c0.n16972_cascade_ ));
    InMux I__9341 (
            .O(N__40876),
            .I(N__40872));
    InMux I__9340 (
            .O(N__40875),
            .I(N__40868));
    LocalMux I__9339 (
            .O(N__40872),
            .I(N__40865));
    InMux I__9338 (
            .O(N__40871),
            .I(N__40862));
    LocalMux I__9337 (
            .O(N__40868),
            .I(N__40857));
    Span4Mux_h I__9336 (
            .O(N__40865),
            .I(N__40852));
    LocalMux I__9335 (
            .O(N__40862),
            .I(N__40852));
    InMux I__9334 (
            .O(N__40861),
            .I(N__40849));
    InMux I__9333 (
            .O(N__40860),
            .I(N__40846));
    Span12Mux_v I__9332 (
            .O(N__40857),
            .I(N__40843));
    Span4Mux_h I__9331 (
            .O(N__40852),
            .I(N__40840));
    LocalMux I__9330 (
            .O(N__40849),
            .I(N__40835));
    LocalMux I__9329 (
            .O(N__40846),
            .I(N__40835));
    Odrv12 I__9328 (
            .O(N__40843),
            .I(data_out_frame2_11_2));
    Odrv4 I__9327 (
            .O(N__40840),
            .I(data_out_frame2_11_2));
    Odrv12 I__9326 (
            .O(N__40835),
            .I(data_out_frame2_11_2));
    InMux I__9325 (
            .O(N__40828),
            .I(N__40825));
    LocalMux I__9324 (
            .O(N__40825),
            .I(N__40822));
    Span4Mux_v I__9323 (
            .O(N__40822),
            .I(N__40819));
    Span4Mux_h I__9322 (
            .O(N__40819),
            .I(N__40816));
    Odrv4 I__9321 (
            .O(N__40816),
            .I(\c0.n10_adj_2281 ));
    InMux I__9320 (
            .O(N__40813),
            .I(N__40810));
    LocalMux I__9319 (
            .O(N__40810),
            .I(N__40807));
    Odrv12 I__9318 (
            .O(N__40807),
            .I(\c0.n17969 ));
    InMux I__9317 (
            .O(N__40804),
            .I(N__40800));
    InMux I__9316 (
            .O(N__40803),
            .I(N__40796));
    LocalMux I__9315 (
            .O(N__40800),
            .I(N__40793));
    InMux I__9314 (
            .O(N__40799),
            .I(N__40790));
    LocalMux I__9313 (
            .O(N__40796),
            .I(N__40783));
    Span4Mux_v I__9312 (
            .O(N__40793),
            .I(N__40783));
    LocalMux I__9311 (
            .O(N__40790),
            .I(N__40783));
    Span4Mux_h I__9310 (
            .O(N__40783),
            .I(N__40778));
    InMux I__9309 (
            .O(N__40782),
            .I(N__40775));
    InMux I__9308 (
            .O(N__40781),
            .I(N__40771));
    Span4Mux_v I__9307 (
            .O(N__40778),
            .I(N__40768));
    LocalMux I__9306 (
            .O(N__40775),
            .I(N__40765));
    InMux I__9305 (
            .O(N__40774),
            .I(N__40762));
    LocalMux I__9304 (
            .O(N__40771),
            .I(data_out_frame2_16_4));
    Odrv4 I__9303 (
            .O(N__40768),
            .I(data_out_frame2_16_4));
    Odrv4 I__9302 (
            .O(N__40765),
            .I(data_out_frame2_16_4));
    LocalMux I__9301 (
            .O(N__40762),
            .I(data_out_frame2_16_4));
    InMux I__9300 (
            .O(N__40753),
            .I(N__40750));
    LocalMux I__9299 (
            .O(N__40750),
            .I(\c0.data_out_frame2_20_4 ));
    CascadeMux I__9298 (
            .O(N__40747),
            .I(\c0.n17972_cascade_ ));
    CascadeMux I__9297 (
            .O(N__40744),
            .I(N__40741));
    InMux I__9296 (
            .O(N__40741),
            .I(N__40738));
    LocalMux I__9295 (
            .O(N__40738),
            .I(N__40735));
    Span4Mux_h I__9294 (
            .O(N__40735),
            .I(N__40732));
    Odrv4 I__9293 (
            .O(N__40732),
            .I(\c0.n17576 ));
    InMux I__9292 (
            .O(N__40729),
            .I(N__40726));
    LocalMux I__9291 (
            .O(N__40726),
            .I(N__40721));
    InMux I__9290 (
            .O(N__40725),
            .I(N__40718));
    InMux I__9289 (
            .O(N__40724),
            .I(N__40714));
    Span4Mux_h I__9288 (
            .O(N__40721),
            .I(N__40711));
    LocalMux I__9287 (
            .O(N__40718),
            .I(N__40708));
    InMux I__9286 (
            .O(N__40717),
            .I(N__40705));
    LocalMux I__9285 (
            .O(N__40714),
            .I(data_out_frame2_8_3));
    Odrv4 I__9284 (
            .O(N__40711),
            .I(data_out_frame2_8_3));
    Odrv4 I__9283 (
            .O(N__40708),
            .I(data_out_frame2_8_3));
    LocalMux I__9282 (
            .O(N__40705),
            .I(data_out_frame2_8_3));
    CascadeMux I__9281 (
            .O(N__40696),
            .I(N__40693));
    InMux I__9280 (
            .O(N__40693),
            .I(N__40689));
    CascadeMux I__9279 (
            .O(N__40692),
            .I(N__40686));
    LocalMux I__9278 (
            .O(N__40689),
            .I(N__40683));
    InMux I__9277 (
            .O(N__40686),
            .I(N__40680));
    Span4Mux_h I__9276 (
            .O(N__40683),
            .I(N__40677));
    LocalMux I__9275 (
            .O(N__40680),
            .I(N__40674));
    Odrv4 I__9274 (
            .O(N__40677),
            .I(\c0.n9839 ));
    Odrv4 I__9273 (
            .O(N__40674),
            .I(\c0.n9839 ));
    InMux I__9272 (
            .O(N__40669),
            .I(N__40665));
    InMux I__9271 (
            .O(N__40668),
            .I(N__40662));
    LocalMux I__9270 (
            .O(N__40665),
            .I(N__40659));
    LocalMux I__9269 (
            .O(N__40662),
            .I(data_out_frame2_18_6));
    Odrv4 I__9268 (
            .O(N__40659),
            .I(data_out_frame2_18_6));
    InMux I__9267 (
            .O(N__40654),
            .I(N__40651));
    LocalMux I__9266 (
            .O(N__40651),
            .I(N__40648));
    Odrv4 I__9265 (
            .O(N__40648),
            .I(\c0.n16994 ));
    InMux I__9264 (
            .O(N__40645),
            .I(N__40642));
    LocalMux I__9263 (
            .O(N__40642),
            .I(N__40638));
    InMux I__9262 (
            .O(N__40641),
            .I(N__40635));
    Span4Mux_v I__9261 (
            .O(N__40638),
            .I(N__40631));
    LocalMux I__9260 (
            .O(N__40635),
            .I(N__40628));
    InMux I__9259 (
            .O(N__40634),
            .I(N__40625));
    Span4Mux_h I__9258 (
            .O(N__40631),
            .I(N__40620));
    Span4Mux_h I__9257 (
            .O(N__40628),
            .I(N__40620));
    LocalMux I__9256 (
            .O(N__40625),
            .I(N__40615));
    Span4Mux_v I__9255 (
            .O(N__40620),
            .I(N__40612));
    InMux I__9254 (
            .O(N__40619),
            .I(N__40609));
    InMux I__9253 (
            .O(N__40618),
            .I(N__40606));
    Span4Mux_s2_v I__9252 (
            .O(N__40615),
            .I(N__40603));
    Odrv4 I__9251 (
            .O(N__40612),
            .I(rand_data_21));
    LocalMux I__9250 (
            .O(N__40609),
            .I(rand_data_21));
    LocalMux I__9249 (
            .O(N__40606),
            .I(rand_data_21));
    Odrv4 I__9248 (
            .O(N__40603),
            .I(rand_data_21));
    InMux I__9247 (
            .O(N__40594),
            .I(N__40591));
    LocalMux I__9246 (
            .O(N__40591),
            .I(N__40588));
    Span4Mux_v I__9245 (
            .O(N__40588),
            .I(N__40585));
    Odrv4 I__9244 (
            .O(N__40585),
            .I(\c0.n28_adj_2294 ));
    CascadeMux I__9243 (
            .O(N__40582),
            .I(\c0.n32_cascade_ ));
    InMux I__9242 (
            .O(N__40579),
            .I(N__40576));
    LocalMux I__9241 (
            .O(N__40576),
            .I(\c0.n31 ));
    InMux I__9240 (
            .O(N__40573),
            .I(N__40570));
    LocalMux I__9239 (
            .O(N__40570),
            .I(N__40566));
    CascadeMux I__9238 (
            .O(N__40569),
            .I(N__40563));
    Span4Mux_h I__9237 (
            .O(N__40566),
            .I(N__40560));
    InMux I__9236 (
            .O(N__40563),
            .I(N__40557));
    Odrv4 I__9235 (
            .O(N__40560),
            .I(rand_setpoint_1));
    LocalMux I__9234 (
            .O(N__40557),
            .I(rand_setpoint_1));
    InMux I__9233 (
            .O(N__40552),
            .I(N__40547));
    InMux I__9232 (
            .O(N__40551),
            .I(N__40544));
    InMux I__9231 (
            .O(N__40550),
            .I(N__40541));
    LocalMux I__9230 (
            .O(N__40547),
            .I(N__40536));
    LocalMux I__9229 (
            .O(N__40544),
            .I(N__40536));
    LocalMux I__9228 (
            .O(N__40541),
            .I(N__40533));
    Span4Mux_v I__9227 (
            .O(N__40536),
            .I(N__40530));
    Odrv4 I__9226 (
            .O(N__40533),
            .I(\c0.data_out_7_1 ));
    Odrv4 I__9225 (
            .O(N__40530),
            .I(\c0.data_out_7_1 ));
    CascadeMux I__9224 (
            .O(N__40525),
            .I(N__40521));
    CascadeMux I__9223 (
            .O(N__40524),
            .I(N__40518));
    InMux I__9222 (
            .O(N__40521),
            .I(N__40515));
    InMux I__9221 (
            .O(N__40518),
            .I(N__40512));
    LocalMux I__9220 (
            .O(N__40515),
            .I(N__40509));
    LocalMux I__9219 (
            .O(N__40512),
            .I(N__40505));
    Span4Mux_v I__9218 (
            .O(N__40509),
            .I(N__40501));
    InMux I__9217 (
            .O(N__40508),
            .I(N__40498));
    Span4Mux_s3_v I__9216 (
            .O(N__40505),
            .I(N__40495));
    InMux I__9215 (
            .O(N__40504),
            .I(N__40492));
    Span4Mux_h I__9214 (
            .O(N__40501),
            .I(N__40487));
    LocalMux I__9213 (
            .O(N__40498),
            .I(N__40487));
    Odrv4 I__9212 (
            .O(N__40495),
            .I(\c0.data_out_9_0 ));
    LocalMux I__9211 (
            .O(N__40492),
            .I(\c0.data_out_9_0 ));
    Odrv4 I__9210 (
            .O(N__40487),
            .I(\c0.data_out_9_0 ));
    InMux I__9209 (
            .O(N__40480),
            .I(N__40475));
    InMux I__9208 (
            .O(N__40479),
            .I(N__40471));
    InMux I__9207 (
            .O(N__40478),
            .I(N__40468));
    LocalMux I__9206 (
            .O(N__40475),
            .I(N__40465));
    InMux I__9205 (
            .O(N__40474),
            .I(N__40462));
    LocalMux I__9204 (
            .O(N__40471),
            .I(N__40459));
    LocalMux I__9203 (
            .O(N__40468),
            .I(N__40456));
    Span4Mux_v I__9202 (
            .O(N__40465),
            .I(N__40449));
    LocalMux I__9201 (
            .O(N__40462),
            .I(N__40449));
    Span4Mux_v I__9200 (
            .O(N__40459),
            .I(N__40444));
    Span4Mux_h I__9199 (
            .O(N__40456),
            .I(N__40444));
    InMux I__9198 (
            .O(N__40455),
            .I(N__40439));
    InMux I__9197 (
            .O(N__40454),
            .I(N__40439));
    Span4Mux_v I__9196 (
            .O(N__40449),
            .I(N__40436));
    Odrv4 I__9195 (
            .O(N__40444),
            .I(\c0.data_out_5_2 ));
    LocalMux I__9194 (
            .O(N__40439),
            .I(\c0.data_out_5_2 ));
    Odrv4 I__9193 (
            .O(N__40436),
            .I(\c0.data_out_5_2 ));
    CascadeMux I__9192 (
            .O(N__40429),
            .I(N__40426));
    InMux I__9191 (
            .O(N__40426),
            .I(N__40420));
    InMux I__9190 (
            .O(N__40425),
            .I(N__40420));
    LocalMux I__9189 (
            .O(N__40420),
            .I(N__40417));
    Odrv4 I__9188 (
            .O(N__40417),
            .I(\c0.n9522 ));
    InMux I__9187 (
            .O(N__40414),
            .I(N__40409));
    CascadeMux I__9186 (
            .O(N__40413),
            .I(N__40405));
    InMux I__9185 (
            .O(N__40412),
            .I(N__40402));
    LocalMux I__9184 (
            .O(N__40409),
            .I(N__40399));
    InMux I__9183 (
            .O(N__40408),
            .I(N__40396));
    InMux I__9182 (
            .O(N__40405),
            .I(N__40393));
    LocalMux I__9181 (
            .O(N__40402),
            .I(N__40386));
    Span4Mux_v I__9180 (
            .O(N__40399),
            .I(N__40386));
    LocalMux I__9179 (
            .O(N__40396),
            .I(N__40386));
    LocalMux I__9178 (
            .O(N__40393),
            .I(N__40381));
    Span4Mux_h I__9177 (
            .O(N__40386),
            .I(N__40378));
    InMux I__9176 (
            .O(N__40385),
            .I(N__40373));
    InMux I__9175 (
            .O(N__40384),
            .I(N__40373));
    Odrv4 I__9174 (
            .O(N__40381),
            .I(data_out_8_1));
    Odrv4 I__9173 (
            .O(N__40378),
            .I(data_out_8_1));
    LocalMux I__9172 (
            .O(N__40373),
            .I(data_out_8_1));
    InMux I__9171 (
            .O(N__40366),
            .I(N__40363));
    LocalMux I__9170 (
            .O(N__40363),
            .I(N__40360));
    Span4Mux_s1_v I__9169 (
            .O(N__40360),
            .I(N__40357));
    Span4Mux_h I__9168 (
            .O(N__40357),
            .I(N__40354));
    Odrv4 I__9167 (
            .O(N__40354),
            .I(\c0.n18077 ));
    InMux I__9166 (
            .O(N__40351),
            .I(N__40348));
    LocalMux I__9165 (
            .O(N__40348),
            .I(N__40345));
    Span4Mux_h I__9164 (
            .O(N__40345),
            .I(N__40342));
    Span4Mux_v I__9163 (
            .O(N__40342),
            .I(N__40337));
    InMux I__9162 (
            .O(N__40341),
            .I(N__40332));
    InMux I__9161 (
            .O(N__40340),
            .I(N__40329));
    Span4Mux_v I__9160 (
            .O(N__40337),
            .I(N__40326));
    InMux I__9159 (
            .O(N__40336),
            .I(N__40323));
    InMux I__9158 (
            .O(N__40335),
            .I(N__40319));
    LocalMux I__9157 (
            .O(N__40332),
            .I(N__40316));
    LocalMux I__9156 (
            .O(N__40329),
            .I(N__40313));
    Span4Mux_v I__9155 (
            .O(N__40326),
            .I(N__40308));
    LocalMux I__9154 (
            .O(N__40323),
            .I(N__40308));
    InMux I__9153 (
            .O(N__40322),
            .I(N__40305));
    LocalMux I__9152 (
            .O(N__40319),
            .I(\c0.data_out_7__2__N_447 ));
    Odrv4 I__9151 (
            .O(N__40316),
            .I(\c0.data_out_7__2__N_447 ));
    Odrv4 I__9150 (
            .O(N__40313),
            .I(\c0.data_out_7__2__N_447 ));
    Odrv4 I__9149 (
            .O(N__40308),
            .I(\c0.data_out_7__2__N_447 ));
    LocalMux I__9148 (
            .O(N__40305),
            .I(\c0.data_out_7__2__N_447 ));
    InMux I__9147 (
            .O(N__40294),
            .I(N__40291));
    LocalMux I__9146 (
            .O(N__40291),
            .I(N__40287));
    CascadeMux I__9145 (
            .O(N__40290),
            .I(N__40284));
    Span4Mux_h I__9144 (
            .O(N__40287),
            .I(N__40281));
    InMux I__9143 (
            .O(N__40284),
            .I(N__40278));
    Odrv4 I__9142 (
            .O(N__40281),
            .I(rand_setpoint_23));
    LocalMux I__9141 (
            .O(N__40278),
            .I(rand_setpoint_23));
    CascadeMux I__9140 (
            .O(N__40273),
            .I(\c0.n17532_cascade_ ));
    InMux I__9139 (
            .O(N__40270),
            .I(N__40266));
    InMux I__9138 (
            .O(N__40269),
            .I(N__40263));
    LocalMux I__9137 (
            .O(N__40266),
            .I(N__40260));
    LocalMux I__9136 (
            .O(N__40263),
            .I(N__40254));
    Span4Mux_s2_v I__9135 (
            .O(N__40260),
            .I(N__40254));
    InMux I__9134 (
            .O(N__40259),
            .I(N__40251));
    Span4Mux_h I__9133 (
            .O(N__40254),
            .I(N__40248));
    LocalMux I__9132 (
            .O(N__40251),
            .I(\c0.data_out_6_7 ));
    Odrv4 I__9131 (
            .O(N__40248),
            .I(\c0.data_out_6_7 ));
    InMux I__9130 (
            .O(N__40243),
            .I(N__40238));
    InMux I__9129 (
            .O(N__40242),
            .I(N__40235));
    InMux I__9128 (
            .O(N__40241),
            .I(N__40232));
    LocalMux I__9127 (
            .O(N__40238),
            .I(N__40229));
    LocalMux I__9126 (
            .O(N__40235),
            .I(N__40223));
    LocalMux I__9125 (
            .O(N__40232),
            .I(N__40223));
    Span4Mux_v I__9124 (
            .O(N__40229),
            .I(N__40220));
    InMux I__9123 (
            .O(N__40228),
            .I(N__40216));
    Span4Mux_s2_v I__9122 (
            .O(N__40223),
            .I(N__40211));
    Span4Mux_h I__9121 (
            .O(N__40220),
            .I(N__40211));
    InMux I__9120 (
            .O(N__40219),
            .I(N__40208));
    LocalMux I__9119 (
            .O(N__40216),
            .I(N__40205));
    Span4Mux_h I__9118 (
            .O(N__40211),
            .I(N__40202));
    LocalMux I__9117 (
            .O(N__40208),
            .I(\c0.data_out_5_5 ));
    Odrv12 I__9116 (
            .O(N__40205),
            .I(\c0.data_out_5_5 ));
    Odrv4 I__9115 (
            .O(N__40202),
            .I(\c0.data_out_5_5 ));
    CascadeMux I__9114 (
            .O(N__40195),
            .I(N__40192));
    InMux I__9113 (
            .O(N__40192),
            .I(N__40189));
    LocalMux I__9112 (
            .O(N__40189),
            .I(N__40184));
    CascadeMux I__9111 (
            .O(N__40188),
            .I(N__40181));
    CascadeMux I__9110 (
            .O(N__40187),
            .I(N__40178));
    Span4Mux_s1_v I__9109 (
            .O(N__40184),
            .I(N__40175));
    InMux I__9108 (
            .O(N__40181),
            .I(N__40170));
    InMux I__9107 (
            .O(N__40178),
            .I(N__40170));
    Span4Mux_h I__9106 (
            .O(N__40175),
            .I(N__40167));
    LocalMux I__9105 (
            .O(N__40170),
            .I(\c0.n17025 ));
    Odrv4 I__9104 (
            .O(N__40167),
            .I(\c0.n17025 ));
    InMux I__9103 (
            .O(N__40162),
            .I(N__40159));
    LocalMux I__9102 (
            .O(N__40159),
            .I(N__40156));
    Odrv12 I__9101 (
            .O(N__40156),
            .I(\c0.n17534 ));
    InMux I__9100 (
            .O(N__40153),
            .I(N__40149));
    InMux I__9099 (
            .O(N__40152),
            .I(N__40143));
    LocalMux I__9098 (
            .O(N__40149),
            .I(N__40140));
    InMux I__9097 (
            .O(N__40148),
            .I(N__40137));
    InMux I__9096 (
            .O(N__40147),
            .I(N__40132));
    InMux I__9095 (
            .O(N__40146),
            .I(N__40132));
    LocalMux I__9094 (
            .O(N__40143),
            .I(N__40129));
    Span4Mux_h I__9093 (
            .O(N__40140),
            .I(N__40126));
    LocalMux I__9092 (
            .O(N__40137),
            .I(N__40121));
    LocalMux I__9091 (
            .O(N__40132),
            .I(N__40121));
    Span4Mux_h I__9090 (
            .O(N__40129),
            .I(N__40118));
    Span4Mux_v I__9089 (
            .O(N__40126),
            .I(N__40115));
    Span4Mux_h I__9088 (
            .O(N__40121),
            .I(N__40112));
    Odrv4 I__9087 (
            .O(N__40118),
            .I(\c0.data_out_frame2_0_3 ));
    Odrv4 I__9086 (
            .O(N__40115),
            .I(\c0.data_out_frame2_0_3 ));
    Odrv4 I__9085 (
            .O(N__40112),
            .I(\c0.data_out_frame2_0_3 ));
    InMux I__9084 (
            .O(N__40105),
            .I(N__40101));
    CascadeMux I__9083 (
            .O(N__40104),
            .I(N__40098));
    LocalMux I__9082 (
            .O(N__40101),
            .I(N__40095));
    InMux I__9081 (
            .O(N__40098),
            .I(N__40092));
    Odrv4 I__9080 (
            .O(N__40095),
            .I(rand_setpoint_5));
    LocalMux I__9079 (
            .O(N__40092),
            .I(rand_setpoint_5));
    InMux I__9078 (
            .O(N__40087),
            .I(N__40084));
    LocalMux I__9077 (
            .O(N__40084),
            .I(N__40081));
    Span4Mux_v I__9076 (
            .O(N__40081),
            .I(N__40074));
    InMux I__9075 (
            .O(N__40080),
            .I(N__40067));
    InMux I__9074 (
            .O(N__40079),
            .I(N__40067));
    InMux I__9073 (
            .O(N__40078),
            .I(N__40067));
    InMux I__9072 (
            .O(N__40077),
            .I(N__40064));
    Odrv4 I__9071 (
            .O(N__40074),
            .I(data_out_8_5));
    LocalMux I__9070 (
            .O(N__40067),
            .I(data_out_8_5));
    LocalMux I__9069 (
            .O(N__40064),
            .I(data_out_8_5));
    InMux I__9068 (
            .O(N__40057),
            .I(N__40053));
    InMux I__9067 (
            .O(N__40056),
            .I(N__40050));
    LocalMux I__9066 (
            .O(N__40053),
            .I(\c0.n28_adj_2287 ));
    LocalMux I__9065 (
            .O(N__40050),
            .I(\c0.n28_adj_2287 ));
    InMux I__9064 (
            .O(N__40045),
            .I(N__40041));
    CascadeMux I__9063 (
            .O(N__40044),
            .I(N__40038));
    LocalMux I__9062 (
            .O(N__40041),
            .I(N__40035));
    InMux I__9061 (
            .O(N__40038),
            .I(N__40032));
    Odrv12 I__9060 (
            .O(N__40035),
            .I(rand_setpoint_6));
    LocalMux I__9059 (
            .O(N__40032),
            .I(rand_setpoint_6));
    InMux I__9058 (
            .O(N__40027),
            .I(N__40018));
    InMux I__9057 (
            .O(N__40026),
            .I(N__40018));
    InMux I__9056 (
            .O(N__40025),
            .I(N__40013));
    InMux I__9055 (
            .O(N__40024),
            .I(N__40013));
    InMux I__9054 (
            .O(N__40023),
            .I(N__40010));
    LocalMux I__9053 (
            .O(N__40018),
            .I(N__40005));
    LocalMux I__9052 (
            .O(N__40013),
            .I(N__40005));
    LocalMux I__9051 (
            .O(N__40010),
            .I(data_out_8_6));
    Odrv4 I__9050 (
            .O(N__40005),
            .I(data_out_8_6));
    InMux I__9049 (
            .O(N__40000),
            .I(N__39997));
    LocalMux I__9048 (
            .O(N__39997),
            .I(N__39994));
    Span4Mux_h I__9047 (
            .O(N__39994),
            .I(N__39990));
    InMux I__9046 (
            .O(N__39993),
            .I(N__39987));
    Span4Mux_h I__9045 (
            .O(N__39990),
            .I(N__39984));
    LocalMux I__9044 (
            .O(N__39987),
            .I(N__39981));
    Odrv4 I__9043 (
            .O(N__39984),
            .I(\c0.data_out_10_7 ));
    Odrv4 I__9042 (
            .O(N__39981),
            .I(\c0.data_out_10_7 ));
    InMux I__9041 (
            .O(N__39976),
            .I(N__39973));
    LocalMux I__9040 (
            .O(N__39973),
            .I(\c0.n8_adj_2166 ));
    CascadeMux I__9039 (
            .O(N__39970),
            .I(N__39967));
    InMux I__9038 (
            .O(N__39967),
            .I(N__39964));
    LocalMux I__9037 (
            .O(N__39964),
            .I(N__39961));
    Odrv12 I__9036 (
            .O(N__39961),
            .I(n10_adj_2425));
    InMux I__9035 (
            .O(N__39958),
            .I(N__39954));
    InMux I__9034 (
            .O(N__39957),
            .I(N__39951));
    LocalMux I__9033 (
            .O(N__39954),
            .I(N__39948));
    LocalMux I__9032 (
            .O(N__39951),
            .I(N__39945));
    Span4Mux_s3_v I__9031 (
            .O(N__39948),
            .I(N__39942));
    Span4Mux_v I__9030 (
            .O(N__39945),
            .I(N__39939));
    Odrv4 I__9029 (
            .O(N__39942),
            .I(\c0.n17055 ));
    Odrv4 I__9028 (
            .O(N__39939),
            .I(\c0.n17055 ));
    InMux I__9027 (
            .O(N__39934),
            .I(N__39929));
    InMux I__9026 (
            .O(N__39933),
            .I(N__39924));
    InMux I__9025 (
            .O(N__39932),
            .I(N__39924));
    LocalMux I__9024 (
            .O(N__39929),
            .I(N__39919));
    LocalMux I__9023 (
            .O(N__39924),
            .I(N__39919));
    Odrv4 I__9022 (
            .O(N__39919),
            .I(\c0.data_out_9_5 ));
    CascadeMux I__9021 (
            .O(N__39916),
            .I(N__39912));
    InMux I__9020 (
            .O(N__39915),
            .I(N__39909));
    InMux I__9019 (
            .O(N__39912),
            .I(N__39906));
    LocalMux I__9018 (
            .O(N__39909),
            .I(N__39903));
    LocalMux I__9017 (
            .O(N__39906),
            .I(N__39900));
    Span4Mux_v I__9016 (
            .O(N__39903),
            .I(N__39895));
    Span4Mux_v I__9015 (
            .O(N__39900),
            .I(N__39892));
    InMux I__9014 (
            .O(N__39899),
            .I(N__39887));
    InMux I__9013 (
            .O(N__39898),
            .I(N__39887));
    Span4Mux_h I__9012 (
            .O(N__39895),
            .I(N__39884));
    Odrv4 I__9011 (
            .O(N__39892),
            .I(\c0.data_out_10_1 ));
    LocalMux I__9010 (
            .O(N__39887),
            .I(\c0.data_out_10_1 ));
    Odrv4 I__9009 (
            .O(N__39884),
            .I(\c0.data_out_10_1 ));
    InMux I__9008 (
            .O(N__39877),
            .I(N__39872));
    InMux I__9007 (
            .O(N__39876),
            .I(N__39868));
    InMux I__9006 (
            .O(N__39875),
            .I(N__39865));
    LocalMux I__9005 (
            .O(N__39872),
            .I(N__39862));
    InMux I__9004 (
            .O(N__39871),
            .I(N__39859));
    LocalMux I__9003 (
            .O(N__39868),
            .I(N__39851));
    LocalMux I__9002 (
            .O(N__39865),
            .I(N__39851));
    Span4Mux_v I__9001 (
            .O(N__39862),
            .I(N__39851));
    LocalMux I__9000 (
            .O(N__39859),
            .I(N__39848));
    InMux I__8999 (
            .O(N__39858),
            .I(N__39845));
    Odrv4 I__8998 (
            .O(N__39851),
            .I(\c0.data_out_8_2 ));
    Odrv4 I__8997 (
            .O(N__39848),
            .I(\c0.data_out_8_2 ));
    LocalMux I__8996 (
            .O(N__39845),
            .I(\c0.data_out_8_2 ));
    CascadeMux I__8995 (
            .O(N__39838),
            .I(N__39834));
    InMux I__8994 (
            .O(N__39837),
            .I(N__39827));
    InMux I__8993 (
            .O(N__39834),
            .I(N__39827));
    InMux I__8992 (
            .O(N__39833),
            .I(N__39822));
    InMux I__8991 (
            .O(N__39832),
            .I(N__39822));
    LocalMux I__8990 (
            .O(N__39827),
            .I(\c0.data_out_10_5 ));
    LocalMux I__8989 (
            .O(N__39822),
            .I(\c0.data_out_10_5 ));
    InMux I__8988 (
            .O(N__39817),
            .I(N__39814));
    LocalMux I__8987 (
            .O(N__39814),
            .I(N__39809));
    InMux I__8986 (
            .O(N__39813),
            .I(N__39806));
    InMux I__8985 (
            .O(N__39812),
            .I(N__39803));
    Span4Mux_s3_v I__8984 (
            .O(N__39809),
            .I(N__39800));
    LocalMux I__8983 (
            .O(N__39806),
            .I(N__39795));
    LocalMux I__8982 (
            .O(N__39803),
            .I(N__39795));
    Span4Mux_h I__8981 (
            .O(N__39800),
            .I(N__39792));
    Odrv4 I__8980 (
            .O(N__39795),
            .I(\c0.data_out_6_4 ));
    Odrv4 I__8979 (
            .O(N__39792),
            .I(\c0.data_out_6_4 ));
    CascadeMux I__8978 (
            .O(N__39787),
            .I(N__39783));
    InMux I__8977 (
            .O(N__39786),
            .I(N__39779));
    InMux I__8976 (
            .O(N__39783),
            .I(N__39776));
    CascadeMux I__8975 (
            .O(N__39782),
            .I(N__39773));
    LocalMux I__8974 (
            .O(N__39779),
            .I(N__39768));
    LocalMux I__8973 (
            .O(N__39776),
            .I(N__39768));
    InMux I__8972 (
            .O(N__39773),
            .I(N__39765));
    Odrv12 I__8971 (
            .O(N__39768),
            .I(\c0.data_out_10_0 ));
    LocalMux I__8970 (
            .O(N__39765),
            .I(\c0.data_out_10_0 ));
    InMux I__8969 (
            .O(N__39760),
            .I(N__39757));
    LocalMux I__8968 (
            .O(N__39757),
            .I(N__39754));
    Span4Mux_v I__8967 (
            .O(N__39754),
            .I(N__39751));
    Span4Mux_h I__8966 (
            .O(N__39751),
            .I(N__39748));
    Odrv4 I__8965 (
            .O(N__39748),
            .I(\c0.n16966 ));
    CascadeMux I__8964 (
            .O(N__39745),
            .I(\c0.n16966_cascade_ ));
    InMux I__8963 (
            .O(N__39742),
            .I(N__39739));
    LocalMux I__8962 (
            .O(N__39739),
            .I(N__39736));
    Odrv4 I__8961 (
            .O(N__39736),
            .I(\c0.n16918 ));
    CascadeMux I__8960 (
            .O(N__39733),
            .I(\c0.n10_adj_2288_cascade_ ));
    InMux I__8959 (
            .O(N__39730),
            .I(N__39724));
    InMux I__8958 (
            .O(N__39729),
            .I(N__39724));
    LocalMux I__8957 (
            .O(N__39724),
            .I(\c0.n17109 ));
    InMux I__8956 (
            .O(N__39721),
            .I(N__39717));
    InMux I__8955 (
            .O(N__39720),
            .I(N__39714));
    LocalMux I__8954 (
            .O(N__39717),
            .I(N__39709));
    LocalMux I__8953 (
            .O(N__39714),
            .I(N__39709));
    Odrv12 I__8952 (
            .O(N__39709),
            .I(\c0.n16990 ));
    CascadeMux I__8951 (
            .O(N__39706),
            .I(N__39701));
    InMux I__8950 (
            .O(N__39705),
            .I(N__39698));
    InMux I__8949 (
            .O(N__39704),
            .I(N__39695));
    InMux I__8948 (
            .O(N__39701),
            .I(N__39692));
    LocalMux I__8947 (
            .O(N__39698),
            .I(N__39689));
    LocalMux I__8946 (
            .O(N__39695),
            .I(N__39686));
    LocalMux I__8945 (
            .O(N__39692),
            .I(N__39683));
    Span4Mux_h I__8944 (
            .O(N__39689),
            .I(N__39680));
    Span4Mux_h I__8943 (
            .O(N__39686),
            .I(N__39675));
    Span4Mux_h I__8942 (
            .O(N__39683),
            .I(N__39675));
    Odrv4 I__8941 (
            .O(N__39680),
            .I(\c0.data_out_6_1 ));
    Odrv4 I__8940 (
            .O(N__39675),
            .I(\c0.data_out_6_1 ));
    InMux I__8939 (
            .O(N__39670),
            .I(N__39661));
    InMux I__8938 (
            .O(N__39669),
            .I(N__39661));
    InMux I__8937 (
            .O(N__39668),
            .I(N__39661));
    LocalMux I__8936 (
            .O(N__39661),
            .I(N__39657));
    InMux I__8935 (
            .O(N__39660),
            .I(N__39654));
    Sp12to4 I__8934 (
            .O(N__39657),
            .I(N__39651));
    LocalMux I__8933 (
            .O(N__39654),
            .I(data_out_frame2_7_0));
    Odrv12 I__8932 (
            .O(N__39651),
            .I(data_out_frame2_7_0));
    InMux I__8931 (
            .O(N__39646),
            .I(N__39643));
    LocalMux I__8930 (
            .O(N__39643),
            .I(N__39640));
    Odrv4 I__8929 (
            .O(N__39640),
            .I(\c0.n17346 ));
    InMux I__8928 (
            .O(N__39637),
            .I(N__39631));
    CascadeMux I__8927 (
            .O(N__39636),
            .I(N__39628));
    InMux I__8926 (
            .O(N__39635),
            .I(N__39623));
    InMux I__8925 (
            .O(N__39634),
            .I(N__39623));
    LocalMux I__8924 (
            .O(N__39631),
            .I(N__39619));
    InMux I__8923 (
            .O(N__39628),
            .I(N__39616));
    LocalMux I__8922 (
            .O(N__39623),
            .I(N__39613));
    InMux I__8921 (
            .O(N__39622),
            .I(N__39610));
    Span12Mux_h I__8920 (
            .O(N__39619),
            .I(N__39605));
    LocalMux I__8919 (
            .O(N__39616),
            .I(N__39605));
    Odrv4 I__8918 (
            .O(N__39613),
            .I(rand_data_26));
    LocalMux I__8917 (
            .O(N__39610),
            .I(rand_data_26));
    Odrv12 I__8916 (
            .O(N__39605),
            .I(rand_data_26));
    InMux I__8915 (
            .O(N__39598),
            .I(N__39594));
    InMux I__8914 (
            .O(N__39597),
            .I(N__39590));
    LocalMux I__8913 (
            .O(N__39594),
            .I(N__39586));
    InMux I__8912 (
            .O(N__39593),
            .I(N__39583));
    LocalMux I__8911 (
            .O(N__39590),
            .I(N__39580));
    InMux I__8910 (
            .O(N__39589),
            .I(N__39577));
    Span4Mux_h I__8909 (
            .O(N__39586),
            .I(N__39573));
    LocalMux I__8908 (
            .O(N__39583),
            .I(N__39568));
    Span4Mux_h I__8907 (
            .O(N__39580),
            .I(N__39568));
    LocalMux I__8906 (
            .O(N__39577),
            .I(N__39565));
    InMux I__8905 (
            .O(N__39576),
            .I(N__39562));
    Span4Mux_v I__8904 (
            .O(N__39573),
            .I(N__39559));
    Span4Mux_v I__8903 (
            .O(N__39568),
            .I(N__39554));
    Span4Mux_h I__8902 (
            .O(N__39565),
            .I(N__39554));
    LocalMux I__8901 (
            .O(N__39562),
            .I(data_out_frame2_14_2));
    Odrv4 I__8900 (
            .O(N__39559),
            .I(data_out_frame2_14_2));
    Odrv4 I__8899 (
            .O(N__39554),
            .I(data_out_frame2_14_2));
    CascadeMux I__8898 (
            .O(N__39547),
            .I(N__39542));
    InMux I__8897 (
            .O(N__39546),
            .I(N__39539));
    InMux I__8896 (
            .O(N__39545),
            .I(N__39534));
    InMux I__8895 (
            .O(N__39542),
            .I(N__39534));
    LocalMux I__8894 (
            .O(N__39539),
            .I(N__39529));
    LocalMux I__8893 (
            .O(N__39534),
            .I(N__39526));
    CascadeMux I__8892 (
            .O(N__39533),
            .I(N__39523));
    InMux I__8891 (
            .O(N__39532),
            .I(N__39519));
    Span4Mux_v I__8890 (
            .O(N__39529),
            .I(N__39514));
    Span4Mux_v I__8889 (
            .O(N__39526),
            .I(N__39514));
    InMux I__8888 (
            .O(N__39523),
            .I(N__39511));
    InMux I__8887 (
            .O(N__39522),
            .I(N__39508));
    LocalMux I__8886 (
            .O(N__39519),
            .I(N__39505));
    Odrv4 I__8885 (
            .O(N__39514),
            .I(rand_data_0));
    LocalMux I__8884 (
            .O(N__39511),
            .I(rand_data_0));
    LocalMux I__8883 (
            .O(N__39508),
            .I(rand_data_0));
    Odrv12 I__8882 (
            .O(N__39505),
            .I(rand_data_0));
    InMux I__8881 (
            .O(N__39496),
            .I(N__39491));
    CascadeMux I__8880 (
            .O(N__39495),
            .I(N__39488));
    InMux I__8879 (
            .O(N__39494),
            .I(N__39485));
    LocalMux I__8878 (
            .O(N__39491),
            .I(N__39482));
    InMux I__8877 (
            .O(N__39488),
            .I(N__39479));
    LocalMux I__8876 (
            .O(N__39485),
            .I(N__39474));
    Span4Mux_v I__8875 (
            .O(N__39482),
            .I(N__39469));
    LocalMux I__8874 (
            .O(N__39479),
            .I(N__39469));
    InMux I__8873 (
            .O(N__39478),
            .I(N__39464));
    InMux I__8872 (
            .O(N__39477),
            .I(N__39464));
    Span4Mux_v I__8871 (
            .O(N__39474),
            .I(N__39459));
    Span4Mux_v I__8870 (
            .O(N__39469),
            .I(N__39459));
    LocalMux I__8869 (
            .O(N__39464),
            .I(data_out_frame2_9_0));
    Odrv4 I__8868 (
            .O(N__39459),
            .I(data_out_frame2_9_0));
    InMux I__8867 (
            .O(N__39454),
            .I(N__39451));
    LocalMux I__8866 (
            .O(N__39451),
            .I(N__39448));
    Span4Mux_h I__8865 (
            .O(N__39448),
            .I(N__39445));
    Odrv4 I__8864 (
            .O(N__39445),
            .I(\c0.n32_adj_2297 ));
    InMux I__8863 (
            .O(N__39442),
            .I(N__39439));
    LocalMux I__8862 (
            .O(N__39439),
            .I(N__39436));
    Span4Mux_v I__8861 (
            .O(N__39436),
            .I(N__39431));
    InMux I__8860 (
            .O(N__39435),
            .I(N__39428));
    InMux I__8859 (
            .O(N__39434),
            .I(N__39425));
    Span4Mux_v I__8858 (
            .O(N__39431),
            .I(N__39422));
    LocalMux I__8857 (
            .O(N__39428),
            .I(N__39419));
    LocalMux I__8856 (
            .O(N__39425),
            .I(N__39416));
    Sp12to4 I__8855 (
            .O(N__39422),
            .I(N__39413));
    Span4Mux_h I__8854 (
            .O(N__39419),
            .I(N__39408));
    Span4Mux_h I__8853 (
            .O(N__39416),
            .I(N__39408));
    Odrv12 I__8852 (
            .O(N__39413),
            .I(\c0.n9814 ));
    Odrv4 I__8851 (
            .O(N__39408),
            .I(\c0.n9814 ));
    InMux I__8850 (
            .O(N__39403),
            .I(N__39400));
    LocalMux I__8849 (
            .O(N__39400),
            .I(N__39397));
    Span4Mux_h I__8848 (
            .O(N__39397),
            .I(N__39393));
    InMux I__8847 (
            .O(N__39396),
            .I(N__39390));
    Odrv4 I__8846 (
            .O(N__39393),
            .I(\c0.n16987 ));
    LocalMux I__8845 (
            .O(N__39390),
            .I(\c0.n16987 ));
    InMux I__8844 (
            .O(N__39385),
            .I(N__39382));
    LocalMux I__8843 (
            .O(N__39382),
            .I(N__39379));
    Odrv4 I__8842 (
            .O(N__39379),
            .I(\c0.n25_adj_2275 ));
    InMux I__8841 (
            .O(N__39376),
            .I(N__39369));
    InMux I__8840 (
            .O(N__39375),
            .I(N__39369));
    InMux I__8839 (
            .O(N__39374),
            .I(N__39365));
    LocalMux I__8838 (
            .O(N__39369),
            .I(N__39362));
    InMux I__8837 (
            .O(N__39368),
            .I(N__39359));
    LocalMux I__8836 (
            .O(N__39365),
            .I(N__39355));
    Span4Mux_v I__8835 (
            .O(N__39362),
            .I(N__39352));
    LocalMux I__8834 (
            .O(N__39359),
            .I(N__39349));
    InMux I__8833 (
            .O(N__39358),
            .I(N__39346));
    Span4Mux_s3_v I__8832 (
            .O(N__39355),
            .I(N__39343));
    Odrv4 I__8831 (
            .O(N__39352),
            .I(rand_data_17));
    Odrv4 I__8830 (
            .O(N__39349),
            .I(rand_data_17));
    LocalMux I__8829 (
            .O(N__39346),
            .I(rand_data_17));
    Odrv4 I__8828 (
            .O(N__39343),
            .I(rand_data_17));
    InMux I__8827 (
            .O(N__39334),
            .I(N__39330));
    InMux I__8826 (
            .O(N__39333),
            .I(N__39327));
    LocalMux I__8825 (
            .O(N__39330),
            .I(N__39322));
    LocalMux I__8824 (
            .O(N__39327),
            .I(N__39319));
    InMux I__8823 (
            .O(N__39326),
            .I(N__39314));
    InMux I__8822 (
            .O(N__39325),
            .I(N__39314));
    Span4Mux_v I__8821 (
            .O(N__39322),
            .I(N__39311));
    Odrv12 I__8820 (
            .O(N__39319),
            .I(data_out_frame2_6_4));
    LocalMux I__8819 (
            .O(N__39314),
            .I(data_out_frame2_6_4));
    Odrv4 I__8818 (
            .O(N__39311),
            .I(data_out_frame2_6_4));
    CascadeMux I__8817 (
            .O(N__39304),
            .I(\c0.n5_adj_2141_cascade_ ));
    InMux I__8816 (
            .O(N__39301),
            .I(N__39298));
    LocalMux I__8815 (
            .O(N__39298),
            .I(N__39295));
    Span4Mux_h I__8814 (
            .O(N__39295),
            .I(N__39292));
    Odrv4 I__8813 (
            .O(N__39292),
            .I(\c0.n17987 ));
    InMux I__8812 (
            .O(N__39289),
            .I(N__39286));
    LocalMux I__8811 (
            .O(N__39286),
            .I(N__39283));
    Span4Mux_h I__8810 (
            .O(N__39283),
            .I(N__39280));
    Odrv4 I__8809 (
            .O(N__39280),
            .I(\c0.n17951 ));
    InMux I__8808 (
            .O(N__39277),
            .I(N__39271));
    InMux I__8807 (
            .O(N__39276),
            .I(N__39268));
    InMux I__8806 (
            .O(N__39275),
            .I(N__39265));
    InMux I__8805 (
            .O(N__39274),
            .I(N__39262));
    LocalMux I__8804 (
            .O(N__39271),
            .I(N__39259));
    LocalMux I__8803 (
            .O(N__39268),
            .I(N__39256));
    LocalMux I__8802 (
            .O(N__39265),
            .I(N__39253));
    LocalMux I__8801 (
            .O(N__39262),
            .I(data_out_frame2_13_3));
    Odrv4 I__8800 (
            .O(N__39259),
            .I(data_out_frame2_13_3));
    Odrv4 I__8799 (
            .O(N__39256),
            .I(data_out_frame2_13_3));
    Odrv4 I__8798 (
            .O(N__39253),
            .I(data_out_frame2_13_3));
    CascadeMux I__8797 (
            .O(N__39244),
            .I(N__39241));
    InMux I__8796 (
            .O(N__39241),
            .I(N__39238));
    LocalMux I__8795 (
            .O(N__39238),
            .I(N__39235));
    Span4Mux_v I__8794 (
            .O(N__39235),
            .I(N__39232));
    Odrv4 I__8793 (
            .O(N__39232),
            .I(\c0.n17954 ));
    InMux I__8792 (
            .O(N__39229),
            .I(N__39226));
    LocalMux I__8791 (
            .O(N__39226),
            .I(N__39223));
    Span4Mux_h I__8790 (
            .O(N__39223),
            .I(N__39220));
    Span4Mux_v I__8789 (
            .O(N__39220),
            .I(N__39217));
    Odrv4 I__8788 (
            .O(N__39217),
            .I(\c0.n18056 ));
    InMux I__8787 (
            .O(N__39214),
            .I(N__39211));
    LocalMux I__8786 (
            .O(N__39211),
            .I(N__39207));
    InMux I__8785 (
            .O(N__39210),
            .I(N__39204));
    Span4Mux_h I__8784 (
            .O(N__39207),
            .I(N__39199));
    LocalMux I__8783 (
            .O(N__39204),
            .I(N__39195));
    InMux I__8782 (
            .O(N__39203),
            .I(N__39192));
    InMux I__8781 (
            .O(N__39202),
            .I(N__39189));
    Span4Mux_v I__8780 (
            .O(N__39199),
            .I(N__39186));
    InMux I__8779 (
            .O(N__39198),
            .I(N__39183));
    Span4Mux_v I__8778 (
            .O(N__39195),
            .I(N__39180));
    LocalMux I__8777 (
            .O(N__39192),
            .I(N__39175));
    LocalMux I__8776 (
            .O(N__39189),
            .I(N__39175));
    Span4Mux_h I__8775 (
            .O(N__39186),
            .I(N__39172));
    LocalMux I__8774 (
            .O(N__39183),
            .I(rand_data_28));
    Odrv4 I__8773 (
            .O(N__39180),
            .I(rand_data_28));
    Odrv12 I__8772 (
            .O(N__39175),
            .I(rand_data_28));
    Odrv4 I__8771 (
            .O(N__39172),
            .I(rand_data_28));
    InMux I__8770 (
            .O(N__39163),
            .I(N__39160));
    LocalMux I__8769 (
            .O(N__39160),
            .I(N__39156));
    CascadeMux I__8768 (
            .O(N__39159),
            .I(N__39153));
    Span4Mux_h I__8767 (
            .O(N__39156),
            .I(N__39148));
    InMux I__8766 (
            .O(N__39153),
            .I(N__39145));
    InMux I__8765 (
            .O(N__39152),
            .I(N__39140));
    InMux I__8764 (
            .O(N__39151),
            .I(N__39140));
    Odrv4 I__8763 (
            .O(N__39148),
            .I(data_out_frame2_15_2));
    LocalMux I__8762 (
            .O(N__39145),
            .I(data_out_frame2_15_2));
    LocalMux I__8761 (
            .O(N__39140),
            .I(data_out_frame2_15_2));
    InMux I__8760 (
            .O(N__39133),
            .I(N__39129));
    InMux I__8759 (
            .O(N__39132),
            .I(N__39123));
    LocalMux I__8758 (
            .O(N__39129),
            .I(N__39120));
    InMux I__8757 (
            .O(N__39128),
            .I(N__39117));
    InMux I__8756 (
            .O(N__39127),
            .I(N__39114));
    InMux I__8755 (
            .O(N__39126),
            .I(N__39111));
    LocalMux I__8754 (
            .O(N__39123),
            .I(N__39108));
    Span4Mux_v I__8753 (
            .O(N__39120),
            .I(N__39103));
    LocalMux I__8752 (
            .O(N__39117),
            .I(N__39103));
    LocalMux I__8751 (
            .O(N__39114),
            .I(data_out_frame2_16_1));
    LocalMux I__8750 (
            .O(N__39111),
            .I(data_out_frame2_16_1));
    Odrv12 I__8749 (
            .O(N__39108),
            .I(data_out_frame2_16_1));
    Odrv4 I__8748 (
            .O(N__39103),
            .I(data_out_frame2_16_1));
    CascadeMux I__8747 (
            .O(N__39094),
            .I(N__39091));
    InMux I__8746 (
            .O(N__39091),
            .I(N__39087));
    InMux I__8745 (
            .O(N__39090),
            .I(N__39084));
    LocalMux I__8744 (
            .O(N__39087),
            .I(N__39077));
    LocalMux I__8743 (
            .O(N__39084),
            .I(N__39077));
    CascadeMux I__8742 (
            .O(N__39083),
            .I(N__39074));
    InMux I__8741 (
            .O(N__39082),
            .I(N__39070));
    Span4Mux_v I__8740 (
            .O(N__39077),
            .I(N__39067));
    InMux I__8739 (
            .O(N__39074),
            .I(N__39064));
    InMux I__8738 (
            .O(N__39073),
            .I(N__39061));
    LocalMux I__8737 (
            .O(N__39070),
            .I(N__39058));
    Odrv4 I__8736 (
            .O(N__39067),
            .I(rand_data_20));
    LocalMux I__8735 (
            .O(N__39064),
            .I(rand_data_20));
    LocalMux I__8734 (
            .O(N__39061),
            .I(rand_data_20));
    Odrv12 I__8733 (
            .O(N__39058),
            .I(rand_data_20));
    InMux I__8732 (
            .O(N__39049),
            .I(N__39045));
    InMux I__8731 (
            .O(N__39048),
            .I(N__39042));
    LocalMux I__8730 (
            .O(N__39045),
            .I(N__39039));
    LocalMux I__8729 (
            .O(N__39042),
            .I(N__39035));
    Span4Mux_h I__8728 (
            .O(N__39039),
            .I(N__39032));
    InMux I__8727 (
            .O(N__39038),
            .I(N__39029));
    Odrv4 I__8726 (
            .O(N__39035),
            .I(\c0.n9749 ));
    Odrv4 I__8725 (
            .O(N__39032),
            .I(\c0.n9749 ));
    LocalMux I__8724 (
            .O(N__39029),
            .I(\c0.n9749 ));
    InMux I__8723 (
            .O(N__39022),
            .I(N__39018));
    InMux I__8722 (
            .O(N__39021),
            .I(N__39015));
    LocalMux I__8721 (
            .O(N__39018),
            .I(N__39010));
    LocalMux I__8720 (
            .O(N__39015),
            .I(N__39007));
    InMux I__8719 (
            .O(N__39014),
            .I(N__39004));
    InMux I__8718 (
            .O(N__39013),
            .I(N__39001));
    Span4Mux_v I__8717 (
            .O(N__39010),
            .I(N__38998));
    Span4Mux_h I__8716 (
            .O(N__39007),
            .I(N__38993));
    LocalMux I__8715 (
            .O(N__39004),
            .I(N__38993));
    LocalMux I__8714 (
            .O(N__39001),
            .I(data_out_frame2_5_1));
    Odrv4 I__8713 (
            .O(N__38998),
            .I(data_out_frame2_5_1));
    Odrv4 I__8712 (
            .O(N__38993),
            .I(data_out_frame2_5_1));
    CascadeMux I__8711 (
            .O(N__38986),
            .I(N__38983));
    InMux I__8710 (
            .O(N__38983),
            .I(N__38980));
    LocalMux I__8709 (
            .O(N__38980),
            .I(\c0.n9776 ));
    InMux I__8708 (
            .O(N__38977),
            .I(N__38973));
    InMux I__8707 (
            .O(N__38976),
            .I(N__38970));
    LocalMux I__8706 (
            .O(N__38973),
            .I(\c0.n9555 ));
    LocalMux I__8705 (
            .O(N__38970),
            .I(\c0.n9555 ));
    InMux I__8704 (
            .O(N__38965),
            .I(N__38962));
    LocalMux I__8703 (
            .O(N__38962),
            .I(N__38959));
    Span4Mux_h I__8702 (
            .O(N__38959),
            .I(N__38956));
    Odrv4 I__8701 (
            .O(N__38956),
            .I(\c0.n16946 ));
    CascadeMux I__8700 (
            .O(N__38953),
            .I(\c0.n22_adj_2207_cascade_ ));
    InMux I__8699 (
            .O(N__38950),
            .I(N__38947));
    LocalMux I__8698 (
            .O(N__38947),
            .I(N__38944));
    Span4Mux_h I__8697 (
            .O(N__38944),
            .I(N__38941));
    Odrv4 I__8696 (
            .O(N__38941),
            .I(\c0.n18_adj_2251 ));
    CascadeMux I__8695 (
            .O(N__38938),
            .I(\c0.n9892_cascade_ ));
    InMux I__8694 (
            .O(N__38935),
            .I(N__38932));
    LocalMux I__8693 (
            .O(N__38932),
            .I(N__38929));
    Odrv4 I__8692 (
            .O(N__38929),
            .I(\c0.n17079 ));
    InMux I__8691 (
            .O(N__38926),
            .I(N__38923));
    LocalMux I__8690 (
            .O(N__38923),
            .I(N__38920));
    Odrv4 I__8689 (
            .O(N__38920),
            .I(\c0.n20_adj_2202 ));
    CascadeMux I__8688 (
            .O(N__38917),
            .I(\c0.n17079_cascade_ ));
    InMux I__8687 (
            .O(N__38914),
            .I(N__38911));
    LocalMux I__8686 (
            .O(N__38911),
            .I(N__38908));
    Odrv12 I__8685 (
            .O(N__38908),
            .I(\c0.n24 ));
    InMux I__8684 (
            .O(N__38905),
            .I(N__38902));
    LocalMux I__8683 (
            .O(N__38902),
            .I(N__38899));
    Span4Mux_h I__8682 (
            .O(N__38899),
            .I(N__38896));
    Odrv4 I__8681 (
            .O(N__38896),
            .I(\c0.data_out_frame2_20_5 ));
    InMux I__8680 (
            .O(N__38893),
            .I(N__38887));
    InMux I__8679 (
            .O(N__38892),
            .I(N__38884));
    InMux I__8678 (
            .O(N__38891),
            .I(N__38881));
    InMux I__8677 (
            .O(N__38890),
            .I(N__38878));
    LocalMux I__8676 (
            .O(N__38887),
            .I(N__38873));
    LocalMux I__8675 (
            .O(N__38884),
            .I(N__38873));
    LocalMux I__8674 (
            .O(N__38881),
            .I(data_out_frame2_10_7));
    LocalMux I__8673 (
            .O(N__38878),
            .I(data_out_frame2_10_7));
    Odrv4 I__8672 (
            .O(N__38873),
            .I(data_out_frame2_10_7));
    CascadeMux I__8671 (
            .O(N__38866),
            .I(\c0.n15_adj_2320_cascade_ ));
    InMux I__8670 (
            .O(N__38863),
            .I(N__38859));
    InMux I__8669 (
            .O(N__38862),
            .I(N__38856));
    LocalMux I__8668 (
            .O(N__38859),
            .I(N__38851));
    LocalMux I__8667 (
            .O(N__38856),
            .I(N__38851));
    Odrv4 I__8666 (
            .O(N__38851),
            .I(\c0.n17088 ));
    InMux I__8665 (
            .O(N__38848),
            .I(N__38845));
    LocalMux I__8664 (
            .O(N__38845),
            .I(N__38842));
    Odrv12 I__8663 (
            .O(N__38842),
            .I(\c0.data_out_frame2_19_2 ));
    InMux I__8662 (
            .O(N__38839),
            .I(N__38836));
    LocalMux I__8661 (
            .O(N__38836),
            .I(\c0.n14_adj_2323 ));
    InMux I__8660 (
            .O(N__38833),
            .I(N__38829));
    InMux I__8659 (
            .O(N__38832),
            .I(N__38826));
    LocalMux I__8658 (
            .O(N__38829),
            .I(\c0.n17052 ));
    LocalMux I__8657 (
            .O(N__38826),
            .I(\c0.n17052 ));
    CascadeMux I__8656 (
            .O(N__38821),
            .I(N__38818));
    InMux I__8655 (
            .O(N__38818),
            .I(N__38815));
    LocalMux I__8654 (
            .O(N__38815),
            .I(N__38812));
    Span4Mux_h I__8653 (
            .O(N__38812),
            .I(N__38809));
    Odrv4 I__8652 (
            .O(N__38809),
            .I(\c0.n17121 ));
    InMux I__8651 (
            .O(N__38806),
            .I(N__38803));
    LocalMux I__8650 (
            .O(N__38803),
            .I(N__38800));
    Span4Mux_h I__8649 (
            .O(N__38800),
            .I(N__38797));
    Odrv4 I__8648 (
            .O(N__38797),
            .I(\c0.n19_adj_2254 ));
    CascadeMux I__8647 (
            .O(N__38794),
            .I(\c0.n21_adj_2255_cascade_ ));
    CascadeMux I__8646 (
            .O(N__38791),
            .I(N__38788));
    InMux I__8645 (
            .O(N__38788),
            .I(N__38785));
    LocalMux I__8644 (
            .O(N__38785),
            .I(N__38782));
    Odrv4 I__8643 (
            .O(N__38782),
            .I(\c0.data_out_frame2_20_3 ));
    InMux I__8642 (
            .O(N__38779),
            .I(N__38776));
    LocalMux I__8641 (
            .O(N__38776),
            .I(N__38770));
    InMux I__8640 (
            .O(N__38775),
            .I(N__38767));
    InMux I__8639 (
            .O(N__38774),
            .I(N__38762));
    InMux I__8638 (
            .O(N__38773),
            .I(N__38762));
    Span4Mux_h I__8637 (
            .O(N__38770),
            .I(N__38759));
    LocalMux I__8636 (
            .O(N__38767),
            .I(data_out_frame2_14_5));
    LocalMux I__8635 (
            .O(N__38762),
            .I(data_out_frame2_14_5));
    Odrv4 I__8634 (
            .O(N__38759),
            .I(data_out_frame2_14_5));
    InMux I__8633 (
            .O(N__38752),
            .I(N__38748));
    InMux I__8632 (
            .O(N__38751),
            .I(N__38745));
    LocalMux I__8631 (
            .O(N__38748),
            .I(N__38742));
    LocalMux I__8630 (
            .O(N__38745),
            .I(N__38739));
    Odrv4 I__8629 (
            .O(N__38742),
            .I(\c0.n17022 ));
    Odrv4 I__8628 (
            .O(N__38739),
            .I(\c0.n17022 ));
    InMux I__8627 (
            .O(N__38734),
            .I(N__38731));
    LocalMux I__8626 (
            .O(N__38731),
            .I(\c0.n26_adj_2273 ));
    CascadeMux I__8625 (
            .O(N__38728),
            .I(N__38725));
    InMux I__8624 (
            .O(N__38725),
            .I(N__38721));
    CascadeMux I__8623 (
            .O(N__38724),
            .I(N__38718));
    LocalMux I__8622 (
            .O(N__38721),
            .I(N__38714));
    InMux I__8621 (
            .O(N__38718),
            .I(N__38711));
    CascadeMux I__8620 (
            .O(N__38717),
            .I(N__38708));
    Span4Mux_h I__8619 (
            .O(N__38714),
            .I(N__38704));
    LocalMux I__8618 (
            .O(N__38711),
            .I(N__38701));
    InMux I__8617 (
            .O(N__38708),
            .I(N__38696));
    InMux I__8616 (
            .O(N__38707),
            .I(N__38696));
    Span4Mux_h I__8615 (
            .O(N__38704),
            .I(N__38693));
    Span4Mux_h I__8614 (
            .O(N__38701),
            .I(N__38690));
    LocalMux I__8613 (
            .O(N__38696),
            .I(\c0.data_out_frame2_0_5 ));
    Odrv4 I__8612 (
            .O(N__38693),
            .I(\c0.data_out_frame2_0_5 ));
    Odrv4 I__8611 (
            .O(N__38690),
            .I(\c0.data_out_frame2_0_5 ));
    InMux I__8610 (
            .O(N__38683),
            .I(N__38680));
    LocalMux I__8609 (
            .O(N__38680),
            .I(N__38676));
    InMux I__8608 (
            .O(N__38679),
            .I(N__38673));
    Odrv4 I__8607 (
            .O(N__38676),
            .I(\c0.n17103 ));
    LocalMux I__8606 (
            .O(N__38673),
            .I(\c0.n17103 ));
    InMux I__8605 (
            .O(N__38668),
            .I(N__38665));
    LocalMux I__8604 (
            .O(N__38665),
            .I(N__38661));
    InMux I__8603 (
            .O(N__38664),
            .I(N__38658));
    Span4Mux_v I__8602 (
            .O(N__38661),
            .I(N__38655));
    LocalMux I__8601 (
            .O(N__38658),
            .I(\c0.n17067 ));
    Odrv4 I__8600 (
            .O(N__38655),
            .I(\c0.n17067 ));
    InMux I__8599 (
            .O(N__38650),
            .I(N__38647));
    LocalMux I__8598 (
            .O(N__38647),
            .I(N__38644));
    Odrv4 I__8597 (
            .O(N__38644),
            .I(\c0.n17100 ));
    CascadeMux I__8596 (
            .O(N__38641),
            .I(N__38637));
    InMux I__8595 (
            .O(N__38640),
            .I(N__38634));
    InMux I__8594 (
            .O(N__38637),
            .I(N__38631));
    LocalMux I__8593 (
            .O(N__38634),
            .I(rand_setpoint_27));
    LocalMux I__8592 (
            .O(N__38631),
            .I(rand_setpoint_27));
    CascadeMux I__8591 (
            .O(N__38626),
            .I(N__38622));
    InMux I__8590 (
            .O(N__38625),
            .I(N__38619));
    InMux I__8589 (
            .O(N__38622),
            .I(N__38616));
    LocalMux I__8588 (
            .O(N__38619),
            .I(rand_setpoint_28));
    LocalMux I__8587 (
            .O(N__38616),
            .I(rand_setpoint_28));
    InMux I__8586 (
            .O(N__38611),
            .I(N__38608));
    LocalMux I__8585 (
            .O(N__38608),
            .I(N__38604));
    InMux I__8584 (
            .O(N__38607),
            .I(N__38601));
    Span4Mux_h I__8583 (
            .O(N__38604),
            .I(N__38597));
    LocalMux I__8582 (
            .O(N__38601),
            .I(N__38594));
    InMux I__8581 (
            .O(N__38600),
            .I(N__38591));
    Span4Mux_v I__8580 (
            .O(N__38597),
            .I(N__38586));
    Span4Mux_h I__8579 (
            .O(N__38594),
            .I(N__38586));
    LocalMux I__8578 (
            .O(N__38591),
            .I(data_out_frame2_7_1));
    Odrv4 I__8577 (
            .O(N__38586),
            .I(data_out_frame2_7_1));
    InMux I__8576 (
            .O(N__38581),
            .I(N__38577));
    InMux I__8575 (
            .O(N__38580),
            .I(N__38574));
    LocalMux I__8574 (
            .O(N__38577),
            .I(N__38571));
    LocalMux I__8573 (
            .O(N__38574),
            .I(N__38564));
    Span4Mux_h I__8572 (
            .O(N__38571),
            .I(N__38564));
    CascadeMux I__8571 (
            .O(N__38570),
            .I(N__38561));
    InMux I__8570 (
            .O(N__38569),
            .I(N__38558));
    Span4Mux_v I__8569 (
            .O(N__38564),
            .I(N__38555));
    InMux I__8568 (
            .O(N__38561),
            .I(N__38552));
    LocalMux I__8567 (
            .O(N__38558),
            .I(data_out_frame2_10_5));
    Odrv4 I__8566 (
            .O(N__38555),
            .I(data_out_frame2_10_5));
    LocalMux I__8565 (
            .O(N__38552),
            .I(data_out_frame2_10_5));
    InMux I__8564 (
            .O(N__38545),
            .I(N__38542));
    LocalMux I__8563 (
            .O(N__38542),
            .I(N__38538));
    InMux I__8562 (
            .O(N__38541),
            .I(N__38535));
    Span4Mux_v I__8561 (
            .O(N__38538),
            .I(N__38532));
    LocalMux I__8560 (
            .O(N__38535),
            .I(N__38529));
    Odrv4 I__8559 (
            .O(N__38532),
            .I(\c0.n9763 ));
    Odrv4 I__8558 (
            .O(N__38529),
            .I(\c0.n9763 ));
    InMux I__8557 (
            .O(N__38524),
            .I(N__38519));
    InMux I__8556 (
            .O(N__38523),
            .I(N__38515));
    InMux I__8555 (
            .O(N__38522),
            .I(N__38511));
    LocalMux I__8554 (
            .O(N__38519),
            .I(N__38508));
    InMux I__8553 (
            .O(N__38518),
            .I(N__38505));
    LocalMux I__8552 (
            .O(N__38515),
            .I(N__38502));
    InMux I__8551 (
            .O(N__38514),
            .I(N__38499));
    LocalMux I__8550 (
            .O(N__38511),
            .I(N__38494));
    Span4Mux_h I__8549 (
            .O(N__38508),
            .I(N__38494));
    LocalMux I__8548 (
            .O(N__38505),
            .I(data_out_frame2_8_2));
    Odrv12 I__8547 (
            .O(N__38502),
            .I(data_out_frame2_8_2));
    LocalMux I__8546 (
            .O(N__38499),
            .I(data_out_frame2_8_2));
    Odrv4 I__8545 (
            .O(N__38494),
            .I(data_out_frame2_8_2));
    InMux I__8544 (
            .O(N__38485),
            .I(N__38482));
    LocalMux I__8543 (
            .O(N__38482),
            .I(N__38479));
    Span4Mux_h I__8542 (
            .O(N__38479),
            .I(N__38476));
    Span4Mux_h I__8541 (
            .O(N__38476),
            .I(N__38473));
    Odrv4 I__8540 (
            .O(N__38473),
            .I(\c0.n9916 ));
    CascadeMux I__8539 (
            .O(N__38470),
            .I(N__38466));
    InMux I__8538 (
            .O(N__38469),
            .I(N__38463));
    InMux I__8537 (
            .O(N__38466),
            .I(N__38459));
    LocalMux I__8536 (
            .O(N__38463),
            .I(N__38456));
    InMux I__8535 (
            .O(N__38462),
            .I(N__38452));
    LocalMux I__8534 (
            .O(N__38459),
            .I(N__38447));
    Span4Mux_h I__8533 (
            .O(N__38456),
            .I(N__38447));
    InMux I__8532 (
            .O(N__38455),
            .I(N__38444));
    LocalMux I__8531 (
            .O(N__38452),
            .I(N__38441));
    Span4Mux_v I__8530 (
            .O(N__38447),
            .I(N__38436));
    LocalMux I__8529 (
            .O(N__38444),
            .I(N__38431));
    Span4Mux_h I__8528 (
            .O(N__38441),
            .I(N__38431));
    InMux I__8527 (
            .O(N__38440),
            .I(N__38426));
    InMux I__8526 (
            .O(N__38439),
            .I(N__38426));
    Odrv4 I__8525 (
            .O(N__38436),
            .I(data_out_frame2_12_4));
    Odrv4 I__8524 (
            .O(N__38431),
            .I(data_out_frame2_12_4));
    LocalMux I__8523 (
            .O(N__38426),
            .I(data_out_frame2_12_4));
    InMux I__8522 (
            .O(N__38419),
            .I(N__38416));
    LocalMux I__8521 (
            .O(N__38416),
            .I(N__38412));
    InMux I__8520 (
            .O(N__38415),
            .I(N__38409));
    Odrv12 I__8519 (
            .O(N__38412),
            .I(\c0.n17037 ));
    LocalMux I__8518 (
            .O(N__38409),
            .I(\c0.n17037 ));
    CascadeMux I__8517 (
            .O(N__38404),
            .I(\c0.n16933_cascade_ ));
    InMux I__8516 (
            .O(N__38401),
            .I(N__38398));
    LocalMux I__8515 (
            .O(N__38398),
            .I(\c0.n17_adj_2313 ));
    InMux I__8514 (
            .O(N__38395),
            .I(N__38392));
    LocalMux I__8513 (
            .O(N__38392),
            .I(N__38389));
    Odrv4 I__8512 (
            .O(N__38389),
            .I(\c0.n17960 ));
    InMux I__8511 (
            .O(N__38386),
            .I(N__38383));
    LocalMux I__8510 (
            .O(N__38383),
            .I(\c0.n18125 ));
    InMux I__8509 (
            .O(N__38380),
            .I(N__38376));
    InMux I__8508 (
            .O(N__38379),
            .I(N__38373));
    LocalMux I__8507 (
            .O(N__38376),
            .I(N__38370));
    LocalMux I__8506 (
            .O(N__38373),
            .I(N__38365));
    Span4Mux_s2_v I__8505 (
            .O(N__38370),
            .I(N__38365));
    Odrv4 I__8504 (
            .O(N__38365),
            .I(data_out_2_7));
    CascadeMux I__8503 (
            .O(N__38362),
            .I(N__38358));
    InMux I__8502 (
            .O(N__38361),
            .I(N__38355));
    InMux I__8501 (
            .O(N__38358),
            .I(N__38352));
    LocalMux I__8500 (
            .O(N__38355),
            .I(rand_setpoint_20));
    LocalMux I__8499 (
            .O(N__38352),
            .I(rand_setpoint_20));
    CascadeMux I__8498 (
            .O(N__38347),
            .I(N__38344));
    InMux I__8497 (
            .O(N__38344),
            .I(N__38341));
    LocalMux I__8496 (
            .O(N__38341),
            .I(N__38338));
    Span4Mux_h I__8495 (
            .O(N__38338),
            .I(N__38335));
    Odrv4 I__8494 (
            .O(N__38335),
            .I(\c0.n17518 ));
    CascadeMux I__8493 (
            .O(N__38332),
            .I(N__38328));
    InMux I__8492 (
            .O(N__38331),
            .I(N__38325));
    InMux I__8491 (
            .O(N__38328),
            .I(N__38322));
    LocalMux I__8490 (
            .O(N__38325),
            .I(rand_setpoint_19));
    LocalMux I__8489 (
            .O(N__38322),
            .I(rand_setpoint_19));
    CascadeMux I__8488 (
            .O(N__38317),
            .I(N__38314));
    InMux I__8487 (
            .O(N__38314),
            .I(N__38311));
    LocalMux I__8486 (
            .O(N__38311),
            .I(N__38308));
    Span4Mux_h I__8485 (
            .O(N__38308),
            .I(N__38305));
    Span4Mux_v I__8484 (
            .O(N__38305),
            .I(N__38302));
    Odrv4 I__8483 (
            .O(N__38302),
            .I(\c0.n17514 ));
    CascadeMux I__8482 (
            .O(N__38299),
            .I(N__38295));
    InMux I__8481 (
            .O(N__38298),
            .I(N__38292));
    InMux I__8480 (
            .O(N__38295),
            .I(N__38289));
    LocalMux I__8479 (
            .O(N__38292),
            .I(rand_setpoint_18));
    LocalMux I__8478 (
            .O(N__38289),
            .I(rand_setpoint_18));
    CascadeMux I__8477 (
            .O(N__38284),
            .I(N__38281));
    InMux I__8476 (
            .O(N__38281),
            .I(N__38278));
    LocalMux I__8475 (
            .O(N__38278),
            .I(N__38275));
    Odrv12 I__8474 (
            .O(N__38275),
            .I(\c0.n17507 ));
    CascadeMux I__8473 (
            .O(N__38272),
            .I(N__38268));
    InMux I__8472 (
            .O(N__38271),
            .I(N__38265));
    InMux I__8471 (
            .O(N__38268),
            .I(N__38262));
    LocalMux I__8470 (
            .O(N__38265),
            .I(rand_setpoint_17));
    LocalMux I__8469 (
            .O(N__38262),
            .I(rand_setpoint_17));
    CascadeMux I__8468 (
            .O(N__38257),
            .I(\c0.n17506_cascade_ ));
    InMux I__8467 (
            .O(N__38254),
            .I(N__38250));
    InMux I__8466 (
            .O(N__38253),
            .I(N__38247));
    LocalMux I__8465 (
            .O(N__38250),
            .I(rand_setpoint_26));
    LocalMux I__8464 (
            .O(N__38247),
            .I(rand_setpoint_26));
    CascadeMux I__8463 (
            .O(N__38242),
            .I(N__38238));
    CascadeMux I__8462 (
            .O(N__38241),
            .I(N__38235));
    InMux I__8461 (
            .O(N__38238),
            .I(N__38232));
    InMux I__8460 (
            .O(N__38235),
            .I(N__38229));
    LocalMux I__8459 (
            .O(N__38232),
            .I(rand_setpoint_29));
    LocalMux I__8458 (
            .O(N__38229),
            .I(rand_setpoint_29));
    CascadeMux I__8457 (
            .O(N__38224),
            .I(N__38220));
    InMux I__8456 (
            .O(N__38223),
            .I(N__38217));
    InMux I__8455 (
            .O(N__38220),
            .I(N__38214));
    LocalMux I__8454 (
            .O(N__38217),
            .I(rand_setpoint_24));
    LocalMux I__8453 (
            .O(N__38214),
            .I(rand_setpoint_24));
    CascadeMux I__8452 (
            .O(N__38209),
            .I(N__38206));
    InMux I__8451 (
            .O(N__38206),
            .I(N__38202));
    InMux I__8450 (
            .O(N__38205),
            .I(N__38199));
    LocalMux I__8449 (
            .O(N__38202),
            .I(rand_setpoint_7));
    LocalMux I__8448 (
            .O(N__38199),
            .I(rand_setpoint_7));
    CascadeMux I__8447 (
            .O(N__38194),
            .I(\c0.n8_adj_2169_cascade_ ));
    InMux I__8446 (
            .O(N__38191),
            .I(N__38188));
    LocalMux I__8445 (
            .O(N__38188),
            .I(N__38185));
    Span4Mux_h I__8444 (
            .O(N__38185),
            .I(N__38182));
    Odrv4 I__8443 (
            .O(N__38182),
            .I(n10_adj_2427));
    InMux I__8442 (
            .O(N__38179),
            .I(N__38176));
    LocalMux I__8441 (
            .O(N__38176),
            .I(\c0.n9496 ));
    CascadeMux I__8440 (
            .O(N__38173),
            .I(N__38170));
    InMux I__8439 (
            .O(N__38170),
            .I(N__38167));
    LocalMux I__8438 (
            .O(N__38167),
            .I(\c0.n9716 ));
    CascadeMux I__8437 (
            .O(N__38164),
            .I(N__38160));
    CascadeMux I__8436 (
            .O(N__38163),
            .I(N__38157));
    InMux I__8435 (
            .O(N__38160),
            .I(N__38154));
    InMux I__8434 (
            .O(N__38157),
            .I(N__38151));
    LocalMux I__8433 (
            .O(N__38154),
            .I(rand_setpoint_2));
    LocalMux I__8432 (
            .O(N__38151),
            .I(rand_setpoint_2));
    CascadeMux I__8431 (
            .O(N__38146),
            .I(N__38143));
    InMux I__8430 (
            .O(N__38143),
            .I(N__38140));
    LocalMux I__8429 (
            .O(N__38140),
            .I(N__38137));
    Span4Mux_v I__8428 (
            .O(N__38137),
            .I(N__38134));
    Span4Mux_h I__8427 (
            .O(N__38134),
            .I(N__38131));
    Odrv4 I__8426 (
            .O(N__38131),
            .I(\c0.n17594 ));
    CascadeMux I__8425 (
            .O(N__38128),
            .I(N__38125));
    InMux I__8424 (
            .O(N__38125),
            .I(N__38122));
    LocalMux I__8423 (
            .O(N__38122),
            .I(N__38119));
    Odrv12 I__8422 (
            .O(N__38119),
            .I(\c0.n8_adj_2176 ));
    InMux I__8421 (
            .O(N__38116),
            .I(N__38110));
    InMux I__8420 (
            .O(N__38115),
            .I(N__38110));
    LocalMux I__8419 (
            .O(N__38110),
            .I(\c0.data_out_1_2 ));
    InMux I__8418 (
            .O(N__38107),
            .I(N__38103));
    InMux I__8417 (
            .O(N__38106),
            .I(N__38098));
    LocalMux I__8416 (
            .O(N__38103),
            .I(N__38093));
    InMux I__8415 (
            .O(N__38102),
            .I(N__38088));
    InMux I__8414 (
            .O(N__38101),
            .I(N__38088));
    LocalMux I__8413 (
            .O(N__38098),
            .I(N__38085));
    InMux I__8412 (
            .O(N__38097),
            .I(N__38082));
    InMux I__8411 (
            .O(N__38096),
            .I(N__38079));
    Span4Mux_v I__8410 (
            .O(N__38093),
            .I(N__38072));
    LocalMux I__8409 (
            .O(N__38088),
            .I(N__38072));
    Span4Mux_h I__8408 (
            .O(N__38085),
            .I(N__38072));
    LocalMux I__8407 (
            .O(N__38082),
            .I(data_out_9_2));
    LocalMux I__8406 (
            .O(N__38079),
            .I(data_out_9_2));
    Odrv4 I__8405 (
            .O(N__38072),
            .I(data_out_9_2));
    CascadeMux I__8404 (
            .O(N__38065),
            .I(N__38061));
    CascadeMux I__8403 (
            .O(N__38064),
            .I(N__38058));
    InMux I__8402 (
            .O(N__38061),
            .I(N__38053));
    InMux I__8401 (
            .O(N__38058),
            .I(N__38053));
    LocalMux I__8400 (
            .O(N__38053),
            .I(N__38050));
    Sp12to4 I__8399 (
            .O(N__38050),
            .I(N__38047));
    Span12Mux_s7_v I__8398 (
            .O(N__38047),
            .I(N__38044));
    Odrv12 I__8397 (
            .O(N__38044),
            .I(\c0.n17064 ));
    CascadeMux I__8396 (
            .O(N__38041),
            .I(\c0.n12_adj_2289_cascade_ ));
    InMux I__8395 (
            .O(N__38038),
            .I(N__38035));
    LocalMux I__8394 (
            .O(N__38035),
            .I(N__38030));
    InMux I__8393 (
            .O(N__38034),
            .I(N__38026));
    InMux I__8392 (
            .O(N__38033),
            .I(N__38022));
    Span4Mux_h I__8391 (
            .O(N__38030),
            .I(N__38019));
    InMux I__8390 (
            .O(N__38029),
            .I(N__38016));
    LocalMux I__8389 (
            .O(N__38026),
            .I(N__38013));
    InMux I__8388 (
            .O(N__38025),
            .I(N__38010));
    LocalMux I__8387 (
            .O(N__38022),
            .I(N__38007));
    Odrv4 I__8386 (
            .O(N__38019),
            .I(\c0.data_out_7_6 ));
    LocalMux I__8385 (
            .O(N__38016),
            .I(\c0.data_out_7_6 ));
    Odrv12 I__8384 (
            .O(N__38013),
            .I(\c0.data_out_7_6 ));
    LocalMux I__8383 (
            .O(N__38010),
            .I(\c0.data_out_7_6 ));
    Odrv4 I__8382 (
            .O(N__38007),
            .I(\c0.data_out_7_6 ));
    CascadeMux I__8381 (
            .O(N__37996),
            .I(\c0.n9716_cascade_ ));
    InMux I__8380 (
            .O(N__37993),
            .I(N__37990));
    LocalMux I__8379 (
            .O(N__37990),
            .I(N__37986));
    InMux I__8378 (
            .O(N__37989),
            .I(N__37983));
    Span4Mux_v I__8377 (
            .O(N__37986),
            .I(N__37978));
    LocalMux I__8376 (
            .O(N__37983),
            .I(N__37978));
    Odrv4 I__8375 (
            .O(N__37978),
            .I(\c0.n9728 ));
    CascadeMux I__8374 (
            .O(N__37975),
            .I(\c0.n10_adj_2162_cascade_ ));
    InMux I__8373 (
            .O(N__37972),
            .I(N__37969));
    LocalMux I__8372 (
            .O(N__37969),
            .I(N__37966));
    Odrv12 I__8371 (
            .O(N__37966),
            .I(data_out_9__2__N_367));
    CascadeMux I__8370 (
            .O(N__37963),
            .I(data_out_9__2__N_367_cascade_));
    CascadeMux I__8369 (
            .O(N__37960),
            .I(\c0.n6_adj_2306_cascade_ ));
    InMux I__8368 (
            .O(N__37957),
            .I(N__37954));
    LocalMux I__8367 (
            .O(N__37954),
            .I(N__37950));
    InMux I__8366 (
            .O(N__37953),
            .I(N__37947));
    Span4Mux_v I__8365 (
            .O(N__37950),
            .I(N__37940));
    LocalMux I__8364 (
            .O(N__37947),
            .I(N__37940));
    InMux I__8363 (
            .O(N__37946),
            .I(N__37937));
    InMux I__8362 (
            .O(N__37945),
            .I(N__37933));
    Span4Mux_v I__8361 (
            .O(N__37940),
            .I(N__37930));
    LocalMux I__8360 (
            .O(N__37937),
            .I(N__37927));
    InMux I__8359 (
            .O(N__37936),
            .I(N__37924));
    LocalMux I__8358 (
            .O(N__37933),
            .I(N__37921));
    Odrv4 I__8357 (
            .O(N__37930),
            .I(rand_data_27));
    Odrv4 I__8356 (
            .O(N__37927),
            .I(rand_data_27));
    LocalMux I__8355 (
            .O(N__37924),
            .I(rand_data_27));
    Odrv12 I__8354 (
            .O(N__37921),
            .I(rand_data_27));
    InMux I__8353 (
            .O(N__37912),
            .I(N__37905));
    InMux I__8352 (
            .O(N__37911),
            .I(N__37905));
    InMux I__8351 (
            .O(N__37910),
            .I(N__37902));
    LocalMux I__8350 (
            .O(N__37905),
            .I(N__37898));
    LocalMux I__8349 (
            .O(N__37902),
            .I(N__37893));
    InMux I__8348 (
            .O(N__37901),
            .I(N__37890));
    Span4Mux_v I__8347 (
            .O(N__37898),
            .I(N__37887));
    InMux I__8346 (
            .O(N__37897),
            .I(N__37884));
    InMux I__8345 (
            .O(N__37896),
            .I(N__37881));
    Span12Mux_h I__8344 (
            .O(N__37893),
            .I(N__37876));
    LocalMux I__8343 (
            .O(N__37890),
            .I(N__37876));
    Odrv4 I__8342 (
            .O(N__37887),
            .I(rand_data_9));
    LocalMux I__8341 (
            .O(N__37884),
            .I(rand_data_9));
    LocalMux I__8340 (
            .O(N__37881),
            .I(rand_data_9));
    Odrv12 I__8339 (
            .O(N__37876),
            .I(rand_data_9));
    InMux I__8338 (
            .O(N__37867),
            .I(N__37864));
    LocalMux I__8337 (
            .O(N__37864),
            .I(N__37860));
    InMux I__8336 (
            .O(N__37863),
            .I(N__37857));
    Span4Mux_v I__8335 (
            .O(N__37860),
            .I(N__37854));
    LocalMux I__8334 (
            .O(N__37857),
            .I(data_out_frame2_17_1));
    Odrv4 I__8333 (
            .O(N__37854),
            .I(data_out_frame2_17_1));
    InMux I__8332 (
            .O(N__37849),
            .I(N__37844));
    InMux I__8331 (
            .O(N__37848),
            .I(N__37839));
    InMux I__8330 (
            .O(N__37847),
            .I(N__37839));
    LocalMux I__8329 (
            .O(N__37844),
            .I(N__37834));
    LocalMux I__8328 (
            .O(N__37839),
            .I(N__37831));
    InMux I__8327 (
            .O(N__37838),
            .I(N__37828));
    InMux I__8326 (
            .O(N__37837),
            .I(N__37825));
    Span4Mux_v I__8325 (
            .O(N__37834),
            .I(N__37822));
    Span12Mux_v I__8324 (
            .O(N__37831),
            .I(N__37819));
    LocalMux I__8323 (
            .O(N__37828),
            .I(N__37816));
    LocalMux I__8322 (
            .O(N__37825),
            .I(data_out_frame2_10_4));
    Odrv4 I__8321 (
            .O(N__37822),
            .I(data_out_frame2_10_4));
    Odrv12 I__8320 (
            .O(N__37819),
            .I(data_out_frame2_10_4));
    Odrv4 I__8319 (
            .O(N__37816),
            .I(data_out_frame2_10_4));
    CascadeMux I__8318 (
            .O(N__37807),
            .I(N__37804));
    InMux I__8317 (
            .O(N__37804),
            .I(N__37801));
    LocalMux I__8316 (
            .O(N__37801),
            .I(\c0.n10_adj_2191 ));
    InMux I__8315 (
            .O(N__37798),
            .I(N__37795));
    LocalMux I__8314 (
            .O(N__37795),
            .I(N__37792));
    Odrv12 I__8313 (
            .O(N__37792),
            .I(\c0.n14 ));
    CascadeMux I__8312 (
            .O(N__37789),
            .I(N__37786));
    InMux I__8311 (
            .O(N__37786),
            .I(N__37783));
    LocalMux I__8310 (
            .O(N__37783),
            .I(N__37780));
    Span4Mux_h I__8309 (
            .O(N__37780),
            .I(N__37777));
    Span4Mux_v I__8308 (
            .O(N__37777),
            .I(N__37774));
    Odrv4 I__8307 (
            .O(N__37774),
            .I(\c0.n17528 ));
    InMux I__8306 (
            .O(N__37771),
            .I(N__37768));
    LocalMux I__8305 (
            .O(N__37768),
            .I(N__37763));
    InMux I__8304 (
            .O(N__37767),
            .I(N__37760));
    InMux I__8303 (
            .O(N__37766),
            .I(N__37757));
    Span4Mux_h I__8302 (
            .O(N__37763),
            .I(N__37753));
    LocalMux I__8301 (
            .O(N__37760),
            .I(N__37748));
    LocalMux I__8300 (
            .O(N__37757),
            .I(N__37748));
    InMux I__8299 (
            .O(N__37756),
            .I(N__37745));
    Odrv4 I__8298 (
            .O(N__37753),
            .I(data_out_frame2_15_4));
    Odrv4 I__8297 (
            .O(N__37748),
            .I(data_out_frame2_15_4));
    LocalMux I__8296 (
            .O(N__37745),
            .I(data_out_frame2_15_4));
    CascadeMux I__8295 (
            .O(N__37738),
            .I(N__37733));
    InMux I__8294 (
            .O(N__37737),
            .I(N__37728));
    InMux I__8293 (
            .O(N__37736),
            .I(N__37725));
    InMux I__8292 (
            .O(N__37733),
            .I(N__37722));
    InMux I__8291 (
            .O(N__37732),
            .I(N__37719));
    InMux I__8290 (
            .O(N__37731),
            .I(N__37716));
    LocalMux I__8289 (
            .O(N__37728),
            .I(N__37713));
    LocalMux I__8288 (
            .O(N__37725),
            .I(N__37708));
    LocalMux I__8287 (
            .O(N__37722),
            .I(N__37708));
    LocalMux I__8286 (
            .O(N__37719),
            .I(N__37703));
    LocalMux I__8285 (
            .O(N__37716),
            .I(N__37703));
    Span4Mux_v I__8284 (
            .O(N__37713),
            .I(N__37698));
    Span4Mux_h I__8283 (
            .O(N__37708),
            .I(N__37698));
    Odrv12 I__8282 (
            .O(N__37703),
            .I(data_out_frame2_12_5));
    Odrv4 I__8281 (
            .O(N__37698),
            .I(data_out_frame2_12_5));
    InMux I__8280 (
            .O(N__37693),
            .I(N__37689));
    InMux I__8279 (
            .O(N__37692),
            .I(N__37686));
    LocalMux I__8278 (
            .O(N__37689),
            .I(N__37683));
    LocalMux I__8277 (
            .O(N__37686),
            .I(N__37680));
    Span4Mux_h I__8276 (
            .O(N__37683),
            .I(N__37675));
    Span4Mux_h I__8275 (
            .O(N__37680),
            .I(N__37675));
    Odrv4 I__8274 (
            .O(N__37675),
            .I(\c0.n17049 ));
    CascadeMux I__8273 (
            .O(N__37672),
            .I(N__37669));
    InMux I__8272 (
            .O(N__37669),
            .I(N__37665));
    CascadeMux I__8271 (
            .O(N__37668),
            .I(N__37661));
    LocalMux I__8270 (
            .O(N__37665),
            .I(N__37658));
    InMux I__8269 (
            .O(N__37664),
            .I(N__37653));
    InMux I__8268 (
            .O(N__37661),
            .I(N__37653));
    Span4Mux_h I__8267 (
            .O(N__37658),
            .I(N__37648));
    LocalMux I__8266 (
            .O(N__37653),
            .I(N__37645));
    InMux I__8265 (
            .O(N__37652),
            .I(N__37642));
    InMux I__8264 (
            .O(N__37651),
            .I(N__37639));
    Span4Mux_v I__8263 (
            .O(N__37648),
            .I(N__37636));
    Span4Mux_h I__8262 (
            .O(N__37645),
            .I(N__37631));
    LocalMux I__8261 (
            .O(N__37642),
            .I(N__37631));
    LocalMux I__8260 (
            .O(N__37639),
            .I(data_out_frame2_5_2));
    Odrv4 I__8259 (
            .O(N__37636),
            .I(data_out_frame2_5_2));
    Odrv4 I__8258 (
            .O(N__37631),
            .I(data_out_frame2_5_2));
    InMux I__8257 (
            .O(N__37624),
            .I(N__37620));
    InMux I__8256 (
            .O(N__37623),
            .I(N__37617));
    LocalMux I__8255 (
            .O(N__37620),
            .I(N__37614));
    LocalMux I__8254 (
            .O(N__37617),
            .I(N__37611));
    Odrv4 I__8253 (
            .O(N__37614),
            .I(\c0.n9865 ));
    Odrv4 I__8252 (
            .O(N__37611),
            .I(\c0.n9865 ));
    InMux I__8251 (
            .O(N__37606),
            .I(N__37603));
    LocalMux I__8250 (
            .O(N__37603),
            .I(N__37600));
    Odrv4 I__8249 (
            .O(N__37600),
            .I(\c0.n16908 ));
    CascadeMux I__8248 (
            .O(N__37597),
            .I(\c0.n16908_cascade_ ));
    InMux I__8247 (
            .O(N__37594),
            .I(N__37591));
    LocalMux I__8246 (
            .O(N__37591),
            .I(\c0.n6_adj_2286 ));
    InMux I__8245 (
            .O(N__37588),
            .I(N__37584));
    InMux I__8244 (
            .O(N__37587),
            .I(N__37581));
    LocalMux I__8243 (
            .O(N__37584),
            .I(N__37574));
    LocalMux I__8242 (
            .O(N__37581),
            .I(N__37574));
    InMux I__8241 (
            .O(N__37580),
            .I(N__37571));
    InMux I__8240 (
            .O(N__37579),
            .I(N__37568));
    Span4Mux_v I__8239 (
            .O(N__37574),
            .I(N__37565));
    LocalMux I__8238 (
            .O(N__37571),
            .I(N__37562));
    LocalMux I__8237 (
            .O(N__37568),
            .I(data_out_frame2_14_4));
    Odrv4 I__8236 (
            .O(N__37565),
            .I(data_out_frame2_14_4));
    Odrv12 I__8235 (
            .O(N__37562),
            .I(data_out_frame2_14_4));
    InMux I__8234 (
            .O(N__37555),
            .I(N__37549));
    InMux I__8233 (
            .O(N__37554),
            .I(N__37545));
    InMux I__8232 (
            .O(N__37553),
            .I(N__37542));
    InMux I__8231 (
            .O(N__37552),
            .I(N__37535));
    LocalMux I__8230 (
            .O(N__37549),
            .I(N__37532));
    InMux I__8229 (
            .O(N__37548),
            .I(N__37529));
    LocalMux I__8228 (
            .O(N__37545),
            .I(N__37524));
    LocalMux I__8227 (
            .O(N__37542),
            .I(N__37524));
    InMux I__8226 (
            .O(N__37541),
            .I(N__37519));
    InMux I__8225 (
            .O(N__37540),
            .I(N__37519));
    InMux I__8224 (
            .O(N__37539),
            .I(N__37516));
    InMux I__8223 (
            .O(N__37538),
            .I(N__37513));
    LocalMux I__8222 (
            .O(N__37535),
            .I(N__37508));
    Span4Mux_h I__8221 (
            .O(N__37532),
            .I(N__37508));
    LocalMux I__8220 (
            .O(N__37529),
            .I(N__37505));
    Span4Mux_v I__8219 (
            .O(N__37524),
            .I(N__37498));
    LocalMux I__8218 (
            .O(N__37519),
            .I(N__37498));
    LocalMux I__8217 (
            .O(N__37516),
            .I(N__37498));
    LocalMux I__8216 (
            .O(N__37513),
            .I(N__37495));
    Span4Mux_h I__8215 (
            .O(N__37508),
            .I(N__37492));
    Odrv12 I__8214 (
            .O(N__37505),
            .I(\c0.n5543 ));
    Odrv4 I__8213 (
            .O(N__37498),
            .I(\c0.n5543 ));
    Odrv4 I__8212 (
            .O(N__37495),
            .I(\c0.n5543 ));
    Odrv4 I__8211 (
            .O(N__37492),
            .I(\c0.n5543 ));
    CascadeMux I__8210 (
            .O(N__37483),
            .I(N__37480));
    InMux I__8209 (
            .O(N__37480),
            .I(N__37473));
    InMux I__8208 (
            .O(N__37479),
            .I(N__37467));
    InMux I__8207 (
            .O(N__37478),
            .I(N__37467));
    InMux I__8206 (
            .O(N__37477),
            .I(N__37462));
    InMux I__8205 (
            .O(N__37476),
            .I(N__37462));
    LocalMux I__8204 (
            .O(N__37473),
            .I(N__37459));
    InMux I__8203 (
            .O(N__37472),
            .I(N__37456));
    LocalMux I__8202 (
            .O(N__37467),
            .I(N__37444));
    LocalMux I__8201 (
            .O(N__37462),
            .I(N__37444));
    Span4Mux_v I__8200 (
            .O(N__37459),
            .I(N__37444));
    LocalMux I__8199 (
            .O(N__37456),
            .I(N__37444));
    InMux I__8198 (
            .O(N__37455),
            .I(N__37439));
    InMux I__8197 (
            .O(N__37454),
            .I(N__37439));
    InMux I__8196 (
            .O(N__37453),
            .I(N__37436));
    Span4Mux_v I__8195 (
            .O(N__37444),
            .I(N__37427));
    LocalMux I__8194 (
            .O(N__37439),
            .I(N__37422));
    LocalMux I__8193 (
            .O(N__37436),
            .I(N__37422));
    InMux I__8192 (
            .O(N__37435),
            .I(N__37417));
    InMux I__8191 (
            .O(N__37434),
            .I(N__37417));
    InMux I__8190 (
            .O(N__37433),
            .I(N__37414));
    InMux I__8189 (
            .O(N__37432),
            .I(N__37409));
    InMux I__8188 (
            .O(N__37431),
            .I(N__37409));
    InMux I__8187 (
            .O(N__37430),
            .I(N__37406));
    Sp12to4 I__8186 (
            .O(N__37427),
            .I(N__37403));
    Span4Mux_h I__8185 (
            .O(N__37422),
            .I(N__37400));
    LocalMux I__8184 (
            .O(N__37417),
            .I(\c0.n5545 ));
    LocalMux I__8183 (
            .O(N__37414),
            .I(\c0.n5545 ));
    LocalMux I__8182 (
            .O(N__37409),
            .I(\c0.n5545 ));
    LocalMux I__8181 (
            .O(N__37406),
            .I(\c0.n5545 ));
    Odrv12 I__8180 (
            .O(N__37403),
            .I(\c0.n5545 ));
    Odrv4 I__8179 (
            .O(N__37400),
            .I(\c0.n5545 ));
    InMux I__8178 (
            .O(N__37387),
            .I(N__37384));
    LocalMux I__8177 (
            .O(N__37384),
            .I(N__37379));
    InMux I__8176 (
            .O(N__37383),
            .I(N__37376));
    InMux I__8175 (
            .O(N__37382),
            .I(N__37373));
    Span4Mux_h I__8174 (
            .O(N__37379),
            .I(N__37370));
    LocalMux I__8173 (
            .O(N__37376),
            .I(N__37367));
    LocalMux I__8172 (
            .O(N__37373),
            .I(N__37364));
    Span4Mux_h I__8171 (
            .O(N__37370),
            .I(N__37361));
    Odrv12 I__8170 (
            .O(N__37367),
            .I(n31));
    Odrv4 I__8169 (
            .O(N__37364),
            .I(n31));
    Odrv4 I__8168 (
            .O(N__37361),
            .I(n31));
    InMux I__8167 (
            .O(N__37354),
            .I(N__37350));
    CascadeMux I__8166 (
            .O(N__37353),
            .I(N__37345));
    LocalMux I__8165 (
            .O(N__37350),
            .I(N__37340));
    InMux I__8164 (
            .O(N__37349),
            .I(N__37337));
    InMux I__8163 (
            .O(N__37348),
            .I(N__37334));
    InMux I__8162 (
            .O(N__37345),
            .I(N__37329));
    InMux I__8161 (
            .O(N__37344),
            .I(N__37329));
    InMux I__8160 (
            .O(N__37343),
            .I(N__37326));
    Span4Mux_v I__8159 (
            .O(N__37340),
            .I(N__37323));
    LocalMux I__8158 (
            .O(N__37337),
            .I(rand_data_4));
    LocalMux I__8157 (
            .O(N__37334),
            .I(rand_data_4));
    LocalMux I__8156 (
            .O(N__37329),
            .I(rand_data_4));
    LocalMux I__8155 (
            .O(N__37326),
            .I(rand_data_4));
    Odrv4 I__8154 (
            .O(N__37323),
            .I(rand_data_4));
    CascadeMux I__8153 (
            .O(N__37312),
            .I(n10197_cascade_));
    InMux I__8152 (
            .O(N__37309),
            .I(N__37306));
    LocalMux I__8151 (
            .O(N__37306),
            .I(N__37299));
    CascadeMux I__8150 (
            .O(N__37305),
            .I(N__37296));
    InMux I__8149 (
            .O(N__37304),
            .I(N__37293));
    InMux I__8148 (
            .O(N__37303),
            .I(N__37290));
    InMux I__8147 (
            .O(N__37302),
            .I(N__37287));
    Span4Mux_h I__8146 (
            .O(N__37299),
            .I(N__37284));
    InMux I__8145 (
            .O(N__37296),
            .I(N__37281));
    LocalMux I__8144 (
            .O(N__37293),
            .I(N__37276));
    LocalMux I__8143 (
            .O(N__37290),
            .I(N__37276));
    LocalMux I__8142 (
            .O(N__37287),
            .I(data_out_frame2_9_3));
    Odrv4 I__8141 (
            .O(N__37284),
            .I(data_out_frame2_9_3));
    LocalMux I__8140 (
            .O(N__37281),
            .I(data_out_frame2_9_3));
    Odrv4 I__8139 (
            .O(N__37276),
            .I(data_out_frame2_9_3));
    CascadeMux I__8138 (
            .O(N__37267),
            .I(\c0.n17085_cascade_ ));
    InMux I__8137 (
            .O(N__37264),
            .I(N__37260));
    InMux I__8136 (
            .O(N__37263),
            .I(N__37257));
    LocalMux I__8135 (
            .O(N__37260),
            .I(N__37254));
    LocalMux I__8134 (
            .O(N__37257),
            .I(N__37251));
    Span4Mux_h I__8133 (
            .O(N__37254),
            .I(N__37248));
    Odrv12 I__8132 (
            .O(N__37251),
            .I(\c0.n17073 ));
    Odrv4 I__8131 (
            .O(N__37248),
            .I(\c0.n17073 ));
    InMux I__8130 (
            .O(N__37243),
            .I(N__37240));
    LocalMux I__8129 (
            .O(N__37240),
            .I(N__37237));
    Span4Mux_h I__8128 (
            .O(N__37237),
            .I(N__37233));
    InMux I__8127 (
            .O(N__37236),
            .I(N__37230));
    Span4Mux_v I__8126 (
            .O(N__37233),
            .I(N__37227));
    LocalMux I__8125 (
            .O(N__37230),
            .I(data_out_frame2_18_4));
    Odrv4 I__8124 (
            .O(N__37227),
            .I(data_out_frame2_18_4));
    InMux I__8123 (
            .O(N__37222),
            .I(N__37219));
    LocalMux I__8122 (
            .O(N__37219),
            .I(N__37216));
    Odrv4 I__8121 (
            .O(N__37216),
            .I(\c0.data_out_frame2_19_4 ));
    InMux I__8120 (
            .O(N__37213),
            .I(N__37210));
    LocalMux I__8119 (
            .O(N__37210),
            .I(N__37207));
    Span4Mux_h I__8118 (
            .O(N__37207),
            .I(N__37203));
    InMux I__8117 (
            .O(N__37206),
            .I(N__37200));
    Odrv4 I__8116 (
            .O(N__37203),
            .I(\c0.n9707 ));
    LocalMux I__8115 (
            .O(N__37200),
            .I(\c0.n9707 ));
    InMux I__8114 (
            .O(N__37195),
            .I(N__37192));
    LocalMux I__8113 (
            .O(N__37192),
            .I(N__37188));
    InMux I__8112 (
            .O(N__37191),
            .I(N__37185));
    Span4Mux_v I__8111 (
            .O(N__37188),
            .I(N__37180));
    LocalMux I__8110 (
            .O(N__37185),
            .I(N__37180));
    Sp12to4 I__8109 (
            .O(N__37180),
            .I(N__37177));
    Odrv12 I__8108 (
            .O(N__37177),
            .I(\c0.n16963 ));
    InMux I__8107 (
            .O(N__37174),
            .I(N__37171));
    LocalMux I__8106 (
            .O(N__37171),
            .I(\c0.n9579 ));
    CascadeMux I__8105 (
            .O(N__37168),
            .I(\c0.n9579_cascade_ ));
    InMux I__8104 (
            .O(N__37165),
            .I(N__37162));
    LocalMux I__8103 (
            .O(N__37162),
            .I(N__37159));
    Odrv12 I__8102 (
            .O(N__37159),
            .I(\c0.n10_adj_2307 ));
    InMux I__8101 (
            .O(N__37156),
            .I(N__37153));
    LocalMux I__8100 (
            .O(N__37153),
            .I(\c0.n17957 ));
    InMux I__8099 (
            .O(N__37150),
            .I(N__37144));
    InMux I__8098 (
            .O(N__37149),
            .I(N__37141));
    InMux I__8097 (
            .O(N__37148),
            .I(N__37138));
    InMux I__8096 (
            .O(N__37147),
            .I(N__37135));
    LocalMux I__8095 (
            .O(N__37144),
            .I(data_out_frame2_6_0));
    LocalMux I__8094 (
            .O(N__37141),
            .I(data_out_frame2_6_0));
    LocalMux I__8093 (
            .O(N__37138),
            .I(data_out_frame2_6_0));
    LocalMux I__8092 (
            .O(N__37135),
            .I(data_out_frame2_6_0));
    CascadeMux I__8091 (
            .O(N__37126),
            .I(N__37123));
    InMux I__8090 (
            .O(N__37123),
            .I(N__37120));
    LocalMux I__8089 (
            .O(N__37120),
            .I(\c0.n5_adj_2334 ));
    InMux I__8088 (
            .O(N__37117),
            .I(N__37113));
    CascadeMux I__8087 (
            .O(N__37116),
            .I(N__37110));
    LocalMux I__8086 (
            .O(N__37113),
            .I(N__37106));
    InMux I__8085 (
            .O(N__37110),
            .I(N__37102));
    InMux I__8084 (
            .O(N__37109),
            .I(N__37099));
    Sp12to4 I__8083 (
            .O(N__37106),
            .I(N__37096));
    InMux I__8082 (
            .O(N__37105),
            .I(N__37093));
    LocalMux I__8081 (
            .O(N__37102),
            .I(N__37090));
    LocalMux I__8080 (
            .O(N__37099),
            .I(\c0.data_out_frame2_0_1 ));
    Odrv12 I__8079 (
            .O(N__37096),
            .I(\c0.data_out_frame2_0_1 ));
    LocalMux I__8078 (
            .O(N__37093),
            .I(\c0.data_out_frame2_0_1 ));
    Odrv4 I__8077 (
            .O(N__37090),
            .I(\c0.data_out_frame2_0_1 ));
    InMux I__8076 (
            .O(N__37081),
            .I(N__37078));
    LocalMux I__8075 (
            .O(N__37078),
            .I(N__37074));
    CascadeMux I__8074 (
            .O(N__37077),
            .I(N__37071));
    Span4Mux_h I__8073 (
            .O(N__37074),
            .I(N__37068));
    InMux I__8072 (
            .O(N__37071),
            .I(N__37065));
    Odrv4 I__8071 (
            .O(N__37068),
            .I(\c0.n17124 ));
    LocalMux I__8070 (
            .O(N__37065),
            .I(\c0.n17124 ));
    InMux I__8069 (
            .O(N__37060),
            .I(N__37057));
    LocalMux I__8068 (
            .O(N__37057),
            .I(\c0.n14_adj_2264 ));
    CascadeMux I__8067 (
            .O(N__37054),
            .I(N__37050));
    InMux I__8066 (
            .O(N__37053),
            .I(N__37047));
    InMux I__8065 (
            .O(N__37050),
            .I(N__37044));
    LocalMux I__8064 (
            .O(N__37047),
            .I(N__37036));
    LocalMux I__8063 (
            .O(N__37044),
            .I(N__37036));
    InMux I__8062 (
            .O(N__37043),
            .I(N__37033));
    InMux I__8061 (
            .O(N__37042),
            .I(N__37028));
    InMux I__8060 (
            .O(N__37041),
            .I(N__37028));
    Odrv4 I__8059 (
            .O(N__37036),
            .I(data_out_frame2_16_2));
    LocalMux I__8058 (
            .O(N__37033),
            .I(data_out_frame2_16_2));
    LocalMux I__8057 (
            .O(N__37028),
            .I(data_out_frame2_16_2));
    InMux I__8056 (
            .O(N__37021),
            .I(N__37018));
    LocalMux I__8055 (
            .O(N__37018),
            .I(N__37015));
    Span4Mux_v I__8054 (
            .O(N__37015),
            .I(N__37012));
    Span4Mux_h I__8053 (
            .O(N__37012),
            .I(N__37009));
    Span4Mux_h I__8052 (
            .O(N__37009),
            .I(N__37006));
    Odrv4 I__8051 (
            .O(N__37006),
            .I(\c0.n17031 ));
    InMux I__8050 (
            .O(N__37003),
            .I(N__37000));
    LocalMux I__8049 (
            .O(N__37000),
            .I(N__36997));
    Span4Mux_h I__8048 (
            .O(N__36997),
            .I(N__36994));
    Odrv4 I__8047 (
            .O(N__36994),
            .I(\c0.n17091 ));
    CascadeMux I__8046 (
            .O(N__36991),
            .I(\c0.n17031_cascade_ ));
    InMux I__8045 (
            .O(N__36988),
            .I(N__36984));
    InMux I__8044 (
            .O(N__36987),
            .I(N__36981));
    LocalMux I__8043 (
            .O(N__36984),
            .I(N__36978));
    LocalMux I__8042 (
            .O(N__36981),
            .I(N__36975));
    Span4Mux_h I__8041 (
            .O(N__36978),
            .I(N__36972));
    Odrv4 I__8040 (
            .O(N__36975),
            .I(\c0.n9692 ));
    Odrv4 I__8039 (
            .O(N__36972),
            .I(\c0.n9692 ));
    InMux I__8038 (
            .O(N__36967),
            .I(N__36964));
    LocalMux I__8037 (
            .O(N__36964),
            .I(\c0.n17085 ));
    InMux I__8036 (
            .O(N__36961),
            .I(N__36958));
    LocalMux I__8035 (
            .O(N__36958),
            .I(\c0.n18_adj_2331 ));
    CascadeMux I__8034 (
            .O(N__36955),
            .I(\c0.n17100_cascade_ ));
    CascadeMux I__8033 (
            .O(N__36952),
            .I(\c0.n16_adj_2332_cascade_ ));
    InMux I__8032 (
            .O(N__36949),
            .I(N__36946));
    LocalMux I__8031 (
            .O(N__36946),
            .I(\c0.n20_adj_2333 ));
    CascadeMux I__8030 (
            .O(N__36943),
            .I(N__36940));
    InMux I__8029 (
            .O(N__36940),
            .I(N__36937));
    LocalMux I__8028 (
            .O(N__36937),
            .I(N__36934));
    Span4Mux_h I__8027 (
            .O(N__36934),
            .I(N__36931));
    Odrv4 I__8026 (
            .O(N__36931),
            .I(\c0.data_out_frame2_19_0 ));
    InMux I__8025 (
            .O(N__36928),
            .I(N__36925));
    LocalMux I__8024 (
            .O(N__36925),
            .I(\c0.n9886 ));
    CascadeMux I__8023 (
            .O(N__36922),
            .I(\c0.n12_adj_2263_cascade_ ));
    InMux I__8022 (
            .O(N__36919),
            .I(N__36916));
    LocalMux I__8021 (
            .O(N__36916),
            .I(N__36913));
    Span4Mux_h I__8020 (
            .O(N__36913),
            .I(N__36910));
    Odrv4 I__8019 (
            .O(N__36910),
            .I(\c0.data_out_frame2_20_2 ));
    InMux I__8018 (
            .O(N__36907),
            .I(N__36904));
    LocalMux I__8017 (
            .O(N__36904),
            .I(N__36901));
    Span4Mux_v I__8016 (
            .O(N__36901),
            .I(N__36898));
    Odrv4 I__8015 (
            .O(N__36898),
            .I(\c0.n17112 ));
    CascadeMux I__8014 (
            .O(N__36895),
            .I(\c0.n16_adj_2312_cascade_ ));
    CascadeMux I__8013 (
            .O(N__36892),
            .I(N__36889));
    InMux I__8012 (
            .O(N__36889),
            .I(N__36885));
    InMux I__8011 (
            .O(N__36888),
            .I(N__36882));
    LocalMux I__8010 (
            .O(N__36885),
            .I(\c0.n17097 ));
    LocalMux I__8009 (
            .O(N__36882),
            .I(\c0.n17097 ));
    InMux I__8008 (
            .O(N__36877),
            .I(n15586));
    InMux I__8007 (
            .O(N__36874),
            .I(n15587));
    CascadeMux I__8006 (
            .O(N__36871),
            .I(N__36867));
    InMux I__8005 (
            .O(N__36870),
            .I(N__36864));
    InMux I__8004 (
            .O(N__36867),
            .I(N__36861));
    LocalMux I__8003 (
            .O(N__36864),
            .I(rand_setpoint_30));
    LocalMux I__8002 (
            .O(N__36861),
            .I(rand_setpoint_30));
    InMux I__8001 (
            .O(N__36856),
            .I(n15588));
    InMux I__8000 (
            .O(N__36853),
            .I(n15589));
    InMux I__7999 (
            .O(N__36850),
            .I(N__36846));
    InMux I__7998 (
            .O(N__36849),
            .I(N__36843));
    LocalMux I__7997 (
            .O(N__36846),
            .I(rand_setpoint_31));
    LocalMux I__7996 (
            .O(N__36843),
            .I(rand_setpoint_31));
    InMux I__7995 (
            .O(N__36838),
            .I(N__36835));
    LocalMux I__7994 (
            .O(N__36835),
            .I(N__36832));
    Span4Mux_v I__7993 (
            .O(N__36832),
            .I(N__36829));
    Span4Mux_h I__7992 (
            .O(N__36829),
            .I(N__36824));
    CascadeMux I__7991 (
            .O(N__36828),
            .I(N__36821));
    InMux I__7990 (
            .O(N__36827),
            .I(N__36817));
    Span4Mux_v I__7989 (
            .O(N__36824),
            .I(N__36814));
    InMux I__7988 (
            .O(N__36821),
            .I(N__36811));
    InMux I__7987 (
            .O(N__36820),
            .I(N__36808));
    LocalMux I__7986 (
            .O(N__36817),
            .I(N__36803));
    Span4Mux_v I__7985 (
            .O(N__36814),
            .I(N__36803));
    LocalMux I__7984 (
            .O(N__36811),
            .I(\c0.data_out_7_4 ));
    LocalMux I__7983 (
            .O(N__36808),
            .I(\c0.data_out_7_4 ));
    Odrv4 I__7982 (
            .O(N__36803),
            .I(\c0.data_out_7_4 ));
    CascadeMux I__7981 (
            .O(N__36796),
            .I(\c0.n22_adj_2357_cascade_ ));
    InMux I__7980 (
            .O(N__36793),
            .I(N__36790));
    LocalMux I__7979 (
            .O(N__36790),
            .I(N__36787));
    Span12Mux_v I__7978 (
            .O(N__36787),
            .I(N__36784));
    Odrv12 I__7977 (
            .O(N__36784),
            .I(\c0.tx2.r_Tx_Data_3 ));
    InMux I__7976 (
            .O(N__36781),
            .I(N__36778));
    LocalMux I__7975 (
            .O(N__36778),
            .I(N__36775));
    Span4Mux_h I__7974 (
            .O(N__36775),
            .I(N__36772));
    Odrv4 I__7973 (
            .O(N__36772),
            .I(\c0.n6_adj_2187 ));
    InMux I__7972 (
            .O(N__36769),
            .I(N__36766));
    LocalMux I__7971 (
            .O(N__36766),
            .I(\c0.n18128 ));
    CascadeMux I__7970 (
            .O(N__36763),
            .I(N__36760));
    InMux I__7969 (
            .O(N__36760),
            .I(N__36757));
    LocalMux I__7968 (
            .O(N__36757),
            .I(N__36753));
    CascadeMux I__7967 (
            .O(N__36756),
            .I(N__36750));
    Span4Mux_h I__7966 (
            .O(N__36753),
            .I(N__36747));
    InMux I__7965 (
            .O(N__36750),
            .I(N__36744));
    Span4Mux_v I__7964 (
            .O(N__36747),
            .I(N__36741));
    LocalMux I__7963 (
            .O(N__36744),
            .I(\c0.n16936 ));
    Odrv4 I__7962 (
            .O(N__36741),
            .I(\c0.n16936 ));
    InMux I__7961 (
            .O(N__36736),
            .I(N__36732));
    CascadeMux I__7960 (
            .O(N__36735),
            .I(N__36728));
    LocalMux I__7959 (
            .O(N__36732),
            .I(N__36725));
    InMux I__7958 (
            .O(N__36731),
            .I(N__36722));
    InMux I__7957 (
            .O(N__36728),
            .I(N__36719));
    Span4Mux_h I__7956 (
            .O(N__36725),
            .I(N__36715));
    LocalMux I__7955 (
            .O(N__36722),
            .I(N__36712));
    LocalMux I__7954 (
            .O(N__36719),
            .I(N__36709));
    InMux I__7953 (
            .O(N__36718),
            .I(N__36705));
    Span4Mux_v I__7952 (
            .O(N__36715),
            .I(N__36702));
    Span4Mux_h I__7951 (
            .O(N__36712),
            .I(N__36699));
    Span4Mux_v I__7950 (
            .O(N__36709),
            .I(N__36696));
    InMux I__7949 (
            .O(N__36708),
            .I(N__36693));
    LocalMux I__7948 (
            .O(N__36705),
            .I(N__36690));
    Odrv4 I__7947 (
            .O(N__36702),
            .I(rand_data_19));
    Odrv4 I__7946 (
            .O(N__36699),
            .I(rand_data_19));
    Odrv4 I__7945 (
            .O(N__36696),
            .I(rand_data_19));
    LocalMux I__7944 (
            .O(N__36693),
            .I(rand_data_19));
    Odrv12 I__7943 (
            .O(N__36690),
            .I(rand_data_19));
    InMux I__7942 (
            .O(N__36679),
            .I(n15577));
    InMux I__7941 (
            .O(N__36676),
            .I(n15578));
    InMux I__7940 (
            .O(N__36673),
            .I(n15579));
    CascadeMux I__7939 (
            .O(N__36670),
            .I(N__36666));
    InMux I__7938 (
            .O(N__36669),
            .I(N__36663));
    InMux I__7937 (
            .O(N__36666),
            .I(N__36660));
    LocalMux I__7936 (
            .O(N__36663),
            .I(rand_setpoint_22));
    LocalMux I__7935 (
            .O(N__36660),
            .I(rand_setpoint_22));
    InMux I__7934 (
            .O(N__36655),
            .I(n15580));
    InMux I__7933 (
            .O(N__36652),
            .I(n15581));
    InMux I__7932 (
            .O(N__36649),
            .I(bfn_13_32_0_));
    CascadeMux I__7931 (
            .O(N__36646),
            .I(N__36642));
    InMux I__7930 (
            .O(N__36645),
            .I(N__36639));
    InMux I__7929 (
            .O(N__36642),
            .I(N__36636));
    LocalMux I__7928 (
            .O(N__36639),
            .I(rand_setpoint_25));
    LocalMux I__7927 (
            .O(N__36636),
            .I(rand_setpoint_25));
    InMux I__7926 (
            .O(N__36631),
            .I(n15583));
    InMux I__7925 (
            .O(N__36628),
            .I(n15584));
    InMux I__7924 (
            .O(N__36625),
            .I(n15585));
    InMux I__7923 (
            .O(N__36622),
            .I(N__36616));
    CascadeMux I__7922 (
            .O(N__36621),
            .I(N__36613));
    InMux I__7921 (
            .O(N__36620),
            .I(N__36610));
    InMux I__7920 (
            .O(N__36619),
            .I(N__36606));
    LocalMux I__7919 (
            .O(N__36616),
            .I(N__36603));
    InMux I__7918 (
            .O(N__36613),
            .I(N__36600));
    LocalMux I__7917 (
            .O(N__36610),
            .I(N__36597));
    InMux I__7916 (
            .O(N__36609),
            .I(N__36593));
    LocalMux I__7915 (
            .O(N__36606),
            .I(N__36590));
    Span4Mux_v I__7914 (
            .O(N__36603),
            .I(N__36587));
    LocalMux I__7913 (
            .O(N__36600),
            .I(N__36582));
    Sp12to4 I__7912 (
            .O(N__36597),
            .I(N__36582));
    InMux I__7911 (
            .O(N__36596),
            .I(N__36579));
    LocalMux I__7910 (
            .O(N__36593),
            .I(N__36576));
    Odrv4 I__7909 (
            .O(N__36590),
            .I(rand_data_10));
    Odrv4 I__7908 (
            .O(N__36587),
            .I(rand_data_10));
    Odrv12 I__7907 (
            .O(N__36582),
            .I(rand_data_10));
    LocalMux I__7906 (
            .O(N__36579),
            .I(rand_data_10));
    Odrv12 I__7905 (
            .O(N__36576),
            .I(rand_data_10));
    InMux I__7904 (
            .O(N__36565),
            .I(n15568));
    InMux I__7903 (
            .O(N__36562),
            .I(N__36559));
    LocalMux I__7902 (
            .O(N__36559),
            .I(N__36556));
    Span4Mux_s2_v I__7901 (
            .O(N__36556),
            .I(N__36552));
    CascadeMux I__7900 (
            .O(N__36555),
            .I(N__36549));
    Sp12to4 I__7899 (
            .O(N__36552),
            .I(N__36546));
    InMux I__7898 (
            .O(N__36549),
            .I(N__36543));
    Odrv12 I__7897 (
            .O(N__36546),
            .I(rand_setpoint_11));
    LocalMux I__7896 (
            .O(N__36543),
            .I(rand_setpoint_11));
    InMux I__7895 (
            .O(N__36538),
            .I(n15569));
    InMux I__7894 (
            .O(N__36535),
            .I(N__36532));
    LocalMux I__7893 (
            .O(N__36532),
            .I(N__36529));
    Span4Mux_h I__7892 (
            .O(N__36529),
            .I(N__36525));
    InMux I__7891 (
            .O(N__36528),
            .I(N__36522));
    Odrv4 I__7890 (
            .O(N__36525),
            .I(rand_setpoint_12));
    LocalMux I__7889 (
            .O(N__36522),
            .I(rand_setpoint_12));
    InMux I__7888 (
            .O(N__36517),
            .I(n15570));
    InMux I__7887 (
            .O(N__36514),
            .I(N__36511));
    LocalMux I__7886 (
            .O(N__36511),
            .I(N__36508));
    Span4Mux_h I__7885 (
            .O(N__36508),
            .I(N__36504));
    InMux I__7884 (
            .O(N__36507),
            .I(N__36501));
    Odrv4 I__7883 (
            .O(N__36504),
            .I(rand_setpoint_13));
    LocalMux I__7882 (
            .O(N__36501),
            .I(rand_setpoint_13));
    InMux I__7881 (
            .O(N__36496),
            .I(n15571));
    InMux I__7880 (
            .O(N__36493),
            .I(N__36489));
    CascadeMux I__7879 (
            .O(N__36492),
            .I(N__36486));
    LocalMux I__7878 (
            .O(N__36489),
            .I(N__36483));
    InMux I__7877 (
            .O(N__36486),
            .I(N__36480));
    Odrv4 I__7876 (
            .O(N__36483),
            .I(rand_setpoint_14));
    LocalMux I__7875 (
            .O(N__36480),
            .I(rand_setpoint_14));
    InMux I__7874 (
            .O(N__36475),
            .I(n15572));
    InMux I__7873 (
            .O(N__36472),
            .I(N__36469));
    LocalMux I__7872 (
            .O(N__36469),
            .I(N__36466));
    Span4Mux_s2_v I__7871 (
            .O(N__36466),
            .I(N__36462));
    InMux I__7870 (
            .O(N__36465),
            .I(N__36459));
    Odrv4 I__7869 (
            .O(N__36462),
            .I(rand_setpoint_15));
    LocalMux I__7868 (
            .O(N__36459),
            .I(rand_setpoint_15));
    InMux I__7867 (
            .O(N__36454),
            .I(n15573));
    InMux I__7866 (
            .O(N__36451),
            .I(bfn_13_31_0_));
    InMux I__7865 (
            .O(N__36448),
            .I(n15575));
    InMux I__7864 (
            .O(N__36445),
            .I(n15576));
    InMux I__7863 (
            .O(N__36442),
            .I(N__36436));
    InMux I__7862 (
            .O(N__36441),
            .I(N__36433));
    InMux I__7861 (
            .O(N__36440),
            .I(N__36428));
    InMux I__7860 (
            .O(N__36439),
            .I(N__36428));
    LocalMux I__7859 (
            .O(N__36436),
            .I(N__36425));
    LocalMux I__7858 (
            .O(N__36433),
            .I(N__36419));
    LocalMux I__7857 (
            .O(N__36428),
            .I(N__36419));
    Span4Mux_h I__7856 (
            .O(N__36425),
            .I(N__36415));
    InMux I__7855 (
            .O(N__36424),
            .I(N__36412));
    Span4Mux_v I__7854 (
            .O(N__36419),
            .I(N__36409));
    InMux I__7853 (
            .O(N__36418),
            .I(N__36406));
    Sp12to4 I__7852 (
            .O(N__36415),
            .I(N__36401));
    LocalMux I__7851 (
            .O(N__36412),
            .I(N__36401));
    Odrv4 I__7850 (
            .O(N__36409),
            .I(rand_data_2));
    LocalMux I__7849 (
            .O(N__36406),
            .I(rand_data_2));
    Odrv12 I__7848 (
            .O(N__36401),
            .I(rand_data_2));
    InMux I__7847 (
            .O(N__36394),
            .I(n15560));
    CascadeMux I__7846 (
            .O(N__36391),
            .I(N__36387));
    InMux I__7845 (
            .O(N__36390),
            .I(N__36384));
    InMux I__7844 (
            .O(N__36387),
            .I(N__36381));
    LocalMux I__7843 (
            .O(N__36384),
            .I(rand_setpoint_3));
    LocalMux I__7842 (
            .O(N__36381),
            .I(rand_setpoint_3));
    InMux I__7841 (
            .O(N__36376),
            .I(n15561));
    CascadeMux I__7840 (
            .O(N__36373),
            .I(N__36369));
    InMux I__7839 (
            .O(N__36372),
            .I(N__36366));
    InMux I__7838 (
            .O(N__36369),
            .I(N__36363));
    LocalMux I__7837 (
            .O(N__36366),
            .I(rand_setpoint_4));
    LocalMux I__7836 (
            .O(N__36363),
            .I(rand_setpoint_4));
    InMux I__7835 (
            .O(N__36358),
            .I(n15562));
    InMux I__7834 (
            .O(N__36355),
            .I(n15563));
    InMux I__7833 (
            .O(N__36352),
            .I(n15564));
    InMux I__7832 (
            .O(N__36349),
            .I(n15565));
    CascadeMux I__7831 (
            .O(N__36346),
            .I(N__36343));
    InMux I__7830 (
            .O(N__36343),
            .I(N__36340));
    LocalMux I__7829 (
            .O(N__36340),
            .I(N__36336));
    CascadeMux I__7828 (
            .O(N__36339),
            .I(N__36333));
    Span4Mux_s2_v I__7827 (
            .O(N__36336),
            .I(N__36330));
    InMux I__7826 (
            .O(N__36333),
            .I(N__36327));
    Odrv4 I__7825 (
            .O(N__36330),
            .I(rand_setpoint_8));
    LocalMux I__7824 (
            .O(N__36327),
            .I(rand_setpoint_8));
    InMux I__7823 (
            .O(N__36322),
            .I(bfn_13_30_0_));
    CascadeMux I__7822 (
            .O(N__36319),
            .I(N__36316));
    InMux I__7821 (
            .O(N__36316),
            .I(N__36313));
    LocalMux I__7820 (
            .O(N__36313),
            .I(N__36309));
    CascadeMux I__7819 (
            .O(N__36312),
            .I(N__36306));
    Span4Mux_h I__7818 (
            .O(N__36309),
            .I(N__36303));
    InMux I__7817 (
            .O(N__36306),
            .I(N__36300));
    Odrv4 I__7816 (
            .O(N__36303),
            .I(rand_setpoint_9));
    LocalMux I__7815 (
            .O(N__36300),
            .I(rand_setpoint_9));
    InMux I__7814 (
            .O(N__36295),
            .I(n15567));
    InMux I__7813 (
            .O(N__36292),
            .I(n15552));
    InMux I__7812 (
            .O(N__36289),
            .I(n15553));
    InMux I__7811 (
            .O(N__36286),
            .I(n15554));
    InMux I__7810 (
            .O(N__36283),
            .I(n15555));
    InMux I__7809 (
            .O(N__36280),
            .I(n15556));
    InMux I__7808 (
            .O(N__36277),
            .I(n15557));
    InMux I__7807 (
            .O(N__36274),
            .I(n15558));
    InMux I__7806 (
            .O(N__36271),
            .I(N__36268));
    LocalMux I__7805 (
            .O(N__36268),
            .I(N__36264));
    CascadeMux I__7804 (
            .O(N__36267),
            .I(N__36261));
    Span4Mux_h I__7803 (
            .O(N__36264),
            .I(N__36258));
    InMux I__7802 (
            .O(N__36261),
            .I(N__36255));
    Odrv4 I__7801 (
            .O(N__36258),
            .I(rand_setpoint_0));
    LocalMux I__7800 (
            .O(N__36255),
            .I(rand_setpoint_0));
    InMux I__7799 (
            .O(N__36250),
            .I(N__36246));
    InMux I__7798 (
            .O(N__36249),
            .I(N__36242));
    LocalMux I__7797 (
            .O(N__36246),
            .I(N__36239));
    InMux I__7796 (
            .O(N__36245),
            .I(N__36236));
    LocalMux I__7795 (
            .O(N__36242),
            .I(N__36233));
    Span4Mux_v I__7794 (
            .O(N__36239),
            .I(N__36228));
    LocalMux I__7793 (
            .O(N__36236),
            .I(N__36225));
    Sp12to4 I__7792 (
            .O(N__36233),
            .I(N__36221));
    InMux I__7791 (
            .O(N__36232),
            .I(N__36218));
    InMux I__7790 (
            .O(N__36231),
            .I(N__36215));
    Sp12to4 I__7789 (
            .O(N__36228),
            .I(N__36212));
    Span4Mux_h I__7788 (
            .O(N__36225),
            .I(N__36209));
    InMux I__7787 (
            .O(N__36224),
            .I(N__36206));
    Span12Mux_h I__7786 (
            .O(N__36221),
            .I(N__36201));
    LocalMux I__7785 (
            .O(N__36218),
            .I(N__36201));
    LocalMux I__7784 (
            .O(N__36215),
            .I(rand_data_1));
    Odrv12 I__7783 (
            .O(N__36212),
            .I(rand_data_1));
    Odrv4 I__7782 (
            .O(N__36209),
            .I(rand_data_1));
    LocalMux I__7781 (
            .O(N__36206),
            .I(rand_data_1));
    Odrv12 I__7780 (
            .O(N__36201),
            .I(rand_data_1));
    InMux I__7779 (
            .O(N__36190),
            .I(n15559));
    InMux I__7778 (
            .O(N__36187),
            .I(bfn_13_27_0_));
    InMux I__7777 (
            .O(N__36184),
            .I(n15544));
    InMux I__7776 (
            .O(N__36181),
            .I(n15545));
    InMux I__7775 (
            .O(N__36178),
            .I(n15546));
    InMux I__7774 (
            .O(N__36175),
            .I(n15547));
    InMux I__7773 (
            .O(N__36172),
            .I(n15548));
    InMux I__7772 (
            .O(N__36169),
            .I(n15549));
    InMux I__7771 (
            .O(N__36166),
            .I(n15550));
    InMux I__7770 (
            .O(N__36163),
            .I(bfn_13_28_0_));
    InMux I__7769 (
            .O(N__36160),
            .I(n15533));
    InMux I__7768 (
            .O(N__36157),
            .I(n15534));
    InMux I__7767 (
            .O(N__36154),
            .I(bfn_13_26_0_));
    InMux I__7766 (
            .O(N__36151),
            .I(n15536));
    InMux I__7765 (
            .O(N__36148),
            .I(n15537));
    InMux I__7764 (
            .O(N__36145),
            .I(n15538));
    InMux I__7763 (
            .O(N__36142),
            .I(n15539));
    InMux I__7762 (
            .O(N__36139),
            .I(n15540));
    InMux I__7761 (
            .O(N__36136),
            .I(n15541));
    InMux I__7760 (
            .O(N__36133),
            .I(n15542));
    InMux I__7759 (
            .O(N__36130),
            .I(N__36127));
    LocalMux I__7758 (
            .O(N__36127),
            .I(N__36124));
    Span4Mux_v I__7757 (
            .O(N__36124),
            .I(N__36121));
    Odrv4 I__7756 (
            .O(N__36121),
            .I(\c0.n17981 ));
    CascadeMux I__7755 (
            .O(N__36118),
            .I(\c0.n17984_cascade_ ));
    InMux I__7754 (
            .O(N__36115),
            .I(N__36112));
    LocalMux I__7753 (
            .O(N__36112),
            .I(\c0.n22_adj_2354 ));
    CascadeMux I__7752 (
            .O(N__36109),
            .I(N__36105));
    CascadeMux I__7751 (
            .O(N__36108),
            .I(N__36102));
    InMux I__7750 (
            .O(N__36105),
            .I(N__36097));
    InMux I__7749 (
            .O(N__36102),
            .I(N__36097));
    LocalMux I__7748 (
            .O(N__36097),
            .I(data_out_frame2_17_5));
    InMux I__7747 (
            .O(N__36094),
            .I(bfn_13_25_0_));
    InMux I__7746 (
            .O(N__36091),
            .I(n15528));
    InMux I__7745 (
            .O(N__36088),
            .I(n15529));
    InMux I__7744 (
            .O(N__36085),
            .I(n15530));
    InMux I__7743 (
            .O(N__36082),
            .I(n15531));
    InMux I__7742 (
            .O(N__36079),
            .I(n15532));
    InMux I__7741 (
            .O(N__36076),
            .I(N__36070));
    InMux I__7740 (
            .O(N__36075),
            .I(N__36066));
    InMux I__7739 (
            .O(N__36074),
            .I(N__36061));
    InMux I__7738 (
            .O(N__36073),
            .I(N__36061));
    LocalMux I__7737 (
            .O(N__36070),
            .I(N__36058));
    InMux I__7736 (
            .O(N__36069),
            .I(N__36055));
    LocalMux I__7735 (
            .O(N__36066),
            .I(N__36052));
    LocalMux I__7734 (
            .O(N__36061),
            .I(data_out_frame2_15_3));
    Odrv4 I__7733 (
            .O(N__36058),
            .I(data_out_frame2_15_3));
    LocalMux I__7732 (
            .O(N__36055),
            .I(data_out_frame2_15_3));
    Odrv4 I__7731 (
            .O(N__36052),
            .I(data_out_frame2_15_3));
    InMux I__7730 (
            .O(N__36043),
            .I(N__36038));
    InMux I__7729 (
            .O(N__36042),
            .I(N__36033));
    InMux I__7728 (
            .O(N__36041),
            .I(N__36033));
    LocalMux I__7727 (
            .O(N__36038),
            .I(data_out_frame2_13_4));
    LocalMux I__7726 (
            .O(N__36033),
            .I(data_out_frame2_13_4));
    InMux I__7725 (
            .O(N__36028),
            .I(N__36025));
    LocalMux I__7724 (
            .O(N__36025),
            .I(N__36022));
    Span4Mux_h I__7723 (
            .O(N__36022),
            .I(N__36019));
    Odrv4 I__7722 (
            .O(N__36019),
            .I(\c0.n11 ));
    InMux I__7721 (
            .O(N__36016),
            .I(N__36013));
    LocalMux I__7720 (
            .O(N__36013),
            .I(N__36010));
    Odrv12 I__7719 (
            .O(N__36010),
            .I(\c0.n9810 ));
    InMux I__7718 (
            .O(N__36007),
            .I(N__36004));
    LocalMux I__7717 (
            .O(N__36004),
            .I(N__36001));
    Span4Mux_h I__7716 (
            .O(N__36001),
            .I(N__35998));
    Odrv4 I__7715 (
            .O(N__35998),
            .I(\c0.n17_adj_2193 ));
    CascadeMux I__7714 (
            .O(N__35995),
            .I(\c0.n16_cascade_ ));
    CascadeMux I__7713 (
            .O(N__35992),
            .I(\c0.n17112_cascade_ ));
    CascadeMux I__7712 (
            .O(N__35989),
            .I(\c0.n14_adj_2308_cascade_ ));
    CascadeMux I__7711 (
            .O(N__35986),
            .I(N__35983));
    InMux I__7710 (
            .O(N__35983),
            .I(N__35980));
    LocalMux I__7709 (
            .O(N__35980),
            .I(N__35977));
    Span12Mux_h I__7708 (
            .O(N__35977),
            .I(N__35974));
    Odrv12 I__7707 (
            .O(N__35974),
            .I(\c0.data_out_frame2_19_5 ));
    InMux I__7706 (
            .O(N__35971),
            .I(N__35968));
    LocalMux I__7705 (
            .O(N__35968),
            .I(N__35965));
    Span4Mux_v I__7704 (
            .O(N__35965),
            .I(N__35962));
    Odrv4 I__7703 (
            .O(N__35962),
            .I(\c0.n17933 ));
    InMux I__7702 (
            .O(N__35959),
            .I(N__35956));
    LocalMux I__7701 (
            .O(N__35956),
            .I(N__35953));
    Odrv4 I__7700 (
            .O(N__35953),
            .I(\c0.n5_adj_2317 ));
    InMux I__7699 (
            .O(N__35950),
            .I(N__35947));
    LocalMux I__7698 (
            .O(N__35947),
            .I(N__35944));
    Odrv4 I__7697 (
            .O(N__35944),
            .I(\c0.n16957 ));
    CascadeMux I__7696 (
            .O(N__35941),
            .I(N__35938));
    InMux I__7695 (
            .O(N__35938),
            .I(N__35934));
    InMux I__7694 (
            .O(N__35937),
            .I(N__35931));
    LocalMux I__7693 (
            .O(N__35934),
            .I(N__35928));
    LocalMux I__7692 (
            .O(N__35931),
            .I(N__35925));
    Span4Mux_h I__7691 (
            .O(N__35928),
            .I(N__35922));
    Odrv4 I__7690 (
            .O(N__35925),
            .I(\c0.n17106 ));
    Odrv4 I__7689 (
            .O(N__35922),
            .I(\c0.n17106 ));
    CascadeMux I__7688 (
            .O(N__35917),
            .I(\c0.n16957_cascade_ ));
    InMux I__7687 (
            .O(N__35914),
            .I(N__35911));
    LocalMux I__7686 (
            .O(N__35911),
            .I(\c0.n15_adj_2269 ));
    CascadeMux I__7685 (
            .O(N__35908),
            .I(N__35905));
    InMux I__7684 (
            .O(N__35905),
            .I(N__35902));
    LocalMux I__7683 (
            .O(N__35902),
            .I(N__35899));
    Span4Mux_v I__7682 (
            .O(N__35899),
            .I(N__35896));
    Odrv4 I__7681 (
            .O(N__35896),
            .I(\c0.data_out_frame2_20_1 ));
    InMux I__7680 (
            .O(N__35893),
            .I(N__35887));
    InMux I__7679 (
            .O(N__35892),
            .I(N__35887));
    LocalMux I__7678 (
            .O(N__35887),
            .I(\c0.n17061 ));
    InMux I__7677 (
            .O(N__35884),
            .I(N__35881));
    LocalMux I__7676 (
            .O(N__35881),
            .I(N__35878));
    Odrv4 I__7675 (
            .O(N__35878),
            .I(\c0.data_out_frame2_20_0 ));
    InMux I__7674 (
            .O(N__35875),
            .I(N__35870));
    InMux I__7673 (
            .O(N__35874),
            .I(N__35866));
    InMux I__7672 (
            .O(N__35873),
            .I(N__35863));
    LocalMux I__7671 (
            .O(N__35870),
            .I(N__35860));
    InMux I__7670 (
            .O(N__35869),
            .I(N__35857));
    LocalMux I__7669 (
            .O(N__35866),
            .I(N__35854));
    LocalMux I__7668 (
            .O(N__35863),
            .I(N__35846));
    Span4Mux_h I__7667 (
            .O(N__35860),
            .I(N__35846));
    LocalMux I__7666 (
            .O(N__35857),
            .I(N__35846));
    Span4Mux_v I__7665 (
            .O(N__35854),
            .I(N__35843));
    InMux I__7664 (
            .O(N__35853),
            .I(N__35840));
    Span4Mux_v I__7663 (
            .O(N__35846),
            .I(N__35837));
    Odrv4 I__7662 (
            .O(N__35843),
            .I(\c0.data_out_frame2_0_2 ));
    LocalMux I__7661 (
            .O(N__35840),
            .I(\c0.data_out_frame2_0_2 ));
    Odrv4 I__7660 (
            .O(N__35837),
            .I(\c0.data_out_frame2_0_2 ));
    InMux I__7659 (
            .O(N__35830),
            .I(N__35827));
    LocalMux I__7658 (
            .O(N__35827),
            .I(N__35824));
    Span4Mux_h I__7657 (
            .O(N__35824),
            .I(N__35821));
    Odrv4 I__7656 (
            .O(N__35821),
            .I(\c0.n17578 ));
    InMux I__7655 (
            .O(N__35818),
            .I(N__35815));
    LocalMux I__7654 (
            .O(N__35815),
            .I(N__35811));
    CascadeMux I__7653 (
            .O(N__35814),
            .I(N__35806));
    Span4Mux_v I__7652 (
            .O(N__35811),
            .I(N__35803));
    InMux I__7651 (
            .O(N__35810),
            .I(N__35800));
    InMux I__7650 (
            .O(N__35809),
            .I(N__35797));
    InMux I__7649 (
            .O(N__35806),
            .I(N__35794));
    Span4Mux_h I__7648 (
            .O(N__35803),
            .I(N__35791));
    LocalMux I__7647 (
            .O(N__35800),
            .I(N__35788));
    LocalMux I__7646 (
            .O(N__35797),
            .I(\c0.data_out_frame2_0_4 ));
    LocalMux I__7645 (
            .O(N__35794),
            .I(\c0.data_out_frame2_0_4 ));
    Odrv4 I__7644 (
            .O(N__35791),
            .I(\c0.data_out_frame2_0_4 ));
    Odrv4 I__7643 (
            .O(N__35788),
            .I(\c0.data_out_frame2_0_4 ));
    InMux I__7642 (
            .O(N__35779),
            .I(N__35776));
    LocalMux I__7641 (
            .O(N__35776),
            .I(\c0.n6_adj_2335 ));
    CascadeMux I__7640 (
            .O(N__35773),
            .I(N__35769));
    CascadeMux I__7639 (
            .O(N__35772),
            .I(N__35764));
    InMux I__7638 (
            .O(N__35769),
            .I(N__35753));
    InMux I__7637 (
            .O(N__35768),
            .I(N__35753));
    InMux I__7636 (
            .O(N__35767),
            .I(N__35753));
    InMux I__7635 (
            .O(N__35764),
            .I(N__35746));
    InMux I__7634 (
            .O(N__35763),
            .I(N__35746));
    InMux I__7633 (
            .O(N__35762),
            .I(N__35746));
    InMux I__7632 (
            .O(N__35761),
            .I(N__35742));
    CascadeMux I__7631 (
            .O(N__35760),
            .I(N__35739));
    LocalMux I__7630 (
            .O(N__35753),
            .I(N__35734));
    LocalMux I__7629 (
            .O(N__35746),
            .I(N__35734));
    InMux I__7628 (
            .O(N__35745),
            .I(N__35731));
    LocalMux I__7627 (
            .O(N__35742),
            .I(N__35728));
    InMux I__7626 (
            .O(N__35739),
            .I(N__35725));
    Span4Mux_s3_v I__7625 (
            .O(N__35734),
            .I(N__35722));
    LocalMux I__7624 (
            .O(N__35731),
            .I(N__35717));
    Span4Mux_v I__7623 (
            .O(N__35728),
            .I(N__35717));
    LocalMux I__7622 (
            .O(N__35725),
            .I(N__35714));
    Span4Mux_h I__7621 (
            .O(N__35722),
            .I(N__35711));
    Span4Mux_h I__7620 (
            .O(N__35717),
            .I(N__35708));
    Odrv12 I__7619 (
            .O(N__35714),
            .I(\c0.n10181 ));
    Odrv4 I__7618 (
            .O(N__35711),
            .I(\c0.n10181 ));
    Odrv4 I__7617 (
            .O(N__35708),
            .I(\c0.n10181 ));
    InMux I__7616 (
            .O(N__35701),
            .I(N__35697));
    InMux I__7615 (
            .O(N__35700),
            .I(N__35694));
    LocalMux I__7614 (
            .O(N__35697),
            .I(N__35691));
    LocalMux I__7613 (
            .O(N__35694),
            .I(\c0.data_out_6_6 ));
    Odrv4 I__7612 (
            .O(N__35691),
            .I(\c0.data_out_6_6 ));
    InMux I__7611 (
            .O(N__35686),
            .I(N__35683));
    LocalMux I__7610 (
            .O(N__35683),
            .I(\c0.n5_adj_2300 ));
    CascadeMux I__7609 (
            .O(N__35680),
            .I(\c0.n17555_cascade_ ));
    InMux I__7608 (
            .O(N__35677),
            .I(N__35674));
    LocalMux I__7607 (
            .O(N__35674),
            .I(N__35671));
    Odrv4 I__7606 (
            .O(N__35671),
            .I(\c0.n18035 ));
    InMux I__7605 (
            .O(N__35668),
            .I(N__35665));
    LocalMux I__7604 (
            .O(N__35665),
            .I(N__35662));
    Odrv4 I__7603 (
            .O(N__35662),
            .I(\c0.n17569 ));
    InMux I__7602 (
            .O(N__35659),
            .I(N__35656));
    LocalMux I__7601 (
            .O(N__35656),
            .I(\c0.n16912 ));
    InMux I__7600 (
            .O(N__35653),
            .I(N__35650));
    LocalMux I__7599 (
            .O(N__35650),
            .I(N__35647));
    Span4Mux_h I__7598 (
            .O(N__35647),
            .I(N__35644));
    Odrv4 I__7597 (
            .O(N__35644),
            .I(\c0.n21 ));
    InMux I__7596 (
            .O(N__35641),
            .I(N__35638));
    LocalMux I__7595 (
            .O(N__35638),
            .I(\c0.n17588 ));
    CascadeMux I__7594 (
            .O(N__35635),
            .I(N__35632));
    InMux I__7593 (
            .O(N__35632),
            .I(N__35629));
    LocalMux I__7592 (
            .O(N__35629),
            .I(N__35626));
    Span4Mux_s3_v I__7591 (
            .O(N__35626),
            .I(N__35623));
    Odrv4 I__7590 (
            .O(N__35623),
            .I(\c0.n1 ));
    CascadeMux I__7589 (
            .O(N__35620),
            .I(n18038_cascade_));
    CascadeMux I__7588 (
            .O(N__35617),
            .I(N__35612));
    CascadeMux I__7587 (
            .O(N__35616),
            .I(N__35609));
    InMux I__7586 (
            .O(N__35615),
            .I(N__35606));
    InMux I__7585 (
            .O(N__35612),
            .I(N__35599));
    InMux I__7584 (
            .O(N__35609),
            .I(N__35596));
    LocalMux I__7583 (
            .O(N__35606),
            .I(N__35593));
    InMux I__7582 (
            .O(N__35605),
            .I(N__35590));
    InMux I__7581 (
            .O(N__35604),
            .I(N__35587));
    InMux I__7580 (
            .O(N__35603),
            .I(N__35584));
    InMux I__7579 (
            .O(N__35602),
            .I(N__35581));
    LocalMux I__7578 (
            .O(N__35599),
            .I(N__35576));
    LocalMux I__7577 (
            .O(N__35596),
            .I(N__35576));
    Span4Mux_s3_v I__7576 (
            .O(N__35593),
            .I(N__35571));
    LocalMux I__7575 (
            .O(N__35590),
            .I(N__35571));
    LocalMux I__7574 (
            .O(N__35587),
            .I(N__35568));
    LocalMux I__7573 (
            .O(N__35584),
            .I(N__35565));
    LocalMux I__7572 (
            .O(N__35581),
            .I(N__35561));
    Span4Mux_h I__7571 (
            .O(N__35576),
            .I(N__35556));
    Span4Mux_h I__7570 (
            .O(N__35571),
            .I(N__35556));
    Span4Mux_v I__7569 (
            .O(N__35568),
            .I(N__35551));
    Span4Mux_s1_v I__7568 (
            .O(N__35565),
            .I(N__35551));
    InMux I__7567 (
            .O(N__35564),
            .I(N__35548));
    Span4Mux_v I__7566 (
            .O(N__35561),
            .I(N__35545));
    Span4Mux_h I__7565 (
            .O(N__35556),
            .I(N__35542));
    Span4Mux_h I__7564 (
            .O(N__35551),
            .I(N__35539));
    LocalMux I__7563 (
            .O(N__35548),
            .I(N__35534));
    Sp12to4 I__7562 (
            .O(N__35545),
            .I(N__35534));
    Odrv4 I__7561 (
            .O(N__35542),
            .I(n8730));
    Odrv4 I__7560 (
            .O(N__35539),
            .I(n8730));
    Odrv12 I__7559 (
            .O(N__35534),
            .I(n8730));
    CascadeMux I__7558 (
            .O(N__35527),
            .I(n10_adj_2413_cascade_));
    CascadeMux I__7557 (
            .O(N__35524),
            .I(N__35515));
    InMux I__7556 (
            .O(N__35523),
            .I(N__35512));
    InMux I__7555 (
            .O(N__35522),
            .I(N__35508));
    InMux I__7554 (
            .O(N__35521),
            .I(N__35505));
    InMux I__7553 (
            .O(N__35520),
            .I(N__35500));
    InMux I__7552 (
            .O(N__35519),
            .I(N__35500));
    InMux I__7551 (
            .O(N__35518),
            .I(N__35497));
    InMux I__7550 (
            .O(N__35515),
            .I(N__35494));
    LocalMux I__7549 (
            .O(N__35512),
            .I(N__35491));
    InMux I__7548 (
            .O(N__35511),
            .I(N__35487));
    LocalMux I__7547 (
            .O(N__35508),
            .I(N__35484));
    LocalMux I__7546 (
            .O(N__35505),
            .I(N__35479));
    LocalMux I__7545 (
            .O(N__35500),
            .I(N__35479));
    LocalMux I__7544 (
            .O(N__35497),
            .I(N__35472));
    LocalMux I__7543 (
            .O(N__35494),
            .I(N__35472));
    Span4Mux_h I__7542 (
            .O(N__35491),
            .I(N__35472));
    InMux I__7541 (
            .O(N__35490),
            .I(N__35468));
    LocalMux I__7540 (
            .O(N__35487),
            .I(N__35465));
    Span4Mux_s1_v I__7539 (
            .O(N__35484),
            .I(N__35460));
    Span4Mux_v I__7538 (
            .O(N__35479),
            .I(N__35460));
    Span4Mux_h I__7537 (
            .O(N__35472),
            .I(N__35457));
    InMux I__7536 (
            .O(N__35471),
            .I(N__35454));
    LocalMux I__7535 (
            .O(N__35468),
            .I(byte_transmit_counter_4));
    Odrv4 I__7534 (
            .O(N__35465),
            .I(byte_transmit_counter_4));
    Odrv4 I__7533 (
            .O(N__35460),
            .I(byte_transmit_counter_4));
    Odrv4 I__7532 (
            .O(N__35457),
            .I(byte_transmit_counter_4));
    LocalMux I__7531 (
            .O(N__35454),
            .I(byte_transmit_counter_4));
    InMux I__7530 (
            .O(N__35443),
            .I(N__35440));
    LocalMux I__7529 (
            .O(N__35440),
            .I(N__35437));
    Span4Mux_s3_h I__7528 (
            .O(N__35437),
            .I(N__35434));
    Span4Mux_h I__7527 (
            .O(N__35434),
            .I(N__35430));
    InMux I__7526 (
            .O(N__35433),
            .I(N__35427));
    Span4Mux_h I__7525 (
            .O(N__35430),
            .I(N__35424));
    LocalMux I__7524 (
            .O(N__35427),
            .I(r_Tx_Data_6));
    Odrv4 I__7523 (
            .O(N__35424),
            .I(r_Tx_Data_6));
    InMux I__7522 (
            .O(N__35419),
            .I(N__35416));
    LocalMux I__7521 (
            .O(N__35416),
            .I(N__35413));
    Span4Mux_s1_v I__7520 (
            .O(N__35413),
            .I(N__35410));
    Odrv4 I__7519 (
            .O(N__35410),
            .I(\c0.data_out_1_1 ));
    CascadeMux I__7518 (
            .O(N__35407),
            .I(\c0.n8_adj_2348_cascade_ ));
    InMux I__7517 (
            .O(N__35404),
            .I(N__35401));
    LocalMux I__7516 (
            .O(N__35401),
            .I(N__35398));
    Span4Mux_h I__7515 (
            .O(N__35398),
            .I(N__35395));
    Odrv4 I__7514 (
            .O(N__35395),
            .I(\c0.n17900 ));
    CascadeMux I__7513 (
            .O(N__35392),
            .I(N__35387));
    CascadeMux I__7512 (
            .O(N__35391),
            .I(N__35382));
    CascadeMux I__7511 (
            .O(N__35390),
            .I(N__35377));
    InMux I__7510 (
            .O(N__35387),
            .I(N__35374));
    InMux I__7509 (
            .O(N__35386),
            .I(N__35369));
    InMux I__7508 (
            .O(N__35385),
            .I(N__35369));
    InMux I__7507 (
            .O(N__35382),
            .I(N__35360));
    InMux I__7506 (
            .O(N__35381),
            .I(N__35360));
    InMux I__7505 (
            .O(N__35380),
            .I(N__35360));
    InMux I__7504 (
            .O(N__35377),
            .I(N__35360));
    LocalMux I__7503 (
            .O(N__35374),
            .I(N__35357));
    LocalMux I__7502 (
            .O(N__35369),
            .I(r_Bit_Index_1_adj_2456));
    LocalMux I__7501 (
            .O(N__35360),
            .I(r_Bit_Index_1_adj_2456));
    Odrv4 I__7500 (
            .O(N__35357),
            .I(r_Bit_Index_1_adj_2456));
    InMux I__7499 (
            .O(N__35350),
            .I(N__35344));
    InMux I__7498 (
            .O(N__35349),
            .I(N__35335));
    InMux I__7497 (
            .O(N__35348),
            .I(N__35335));
    InMux I__7496 (
            .O(N__35347),
            .I(N__35335));
    LocalMux I__7495 (
            .O(N__35344),
            .I(N__35332));
    InMux I__7494 (
            .O(N__35343),
            .I(N__35329));
    InMux I__7493 (
            .O(N__35342),
            .I(N__35326));
    LocalMux I__7492 (
            .O(N__35335),
            .I(N__35321));
    Span4Mux_v I__7491 (
            .O(N__35332),
            .I(N__35321));
    LocalMux I__7490 (
            .O(N__35329),
            .I(r_Bit_Index_0_adj_2457));
    LocalMux I__7489 (
            .O(N__35326),
            .I(r_Bit_Index_0_adj_2457));
    Odrv4 I__7488 (
            .O(N__35321),
            .I(r_Bit_Index_0_adj_2457));
    InMux I__7487 (
            .O(N__35314),
            .I(N__35311));
    LocalMux I__7486 (
            .O(N__35311),
            .I(N__35308));
    Odrv4 I__7485 (
            .O(N__35308),
            .I(\c0.tx2.n17903 ));
    InMux I__7484 (
            .O(N__35305),
            .I(N__35301));
    InMux I__7483 (
            .O(N__35304),
            .I(N__35298));
    LocalMux I__7482 (
            .O(N__35301),
            .I(\c0.n16975 ));
    LocalMux I__7481 (
            .O(N__35298),
            .I(\c0.n16975 ));
    CascadeMux I__7480 (
            .O(N__35293),
            .I(\c0.n16978_cascade_ ));
    InMux I__7479 (
            .O(N__35290),
            .I(N__35287));
    LocalMux I__7478 (
            .O(N__35287),
            .I(N__35283));
    InMux I__7477 (
            .O(N__35286),
            .I(N__35280));
    Span4Mux_v I__7476 (
            .O(N__35283),
            .I(N__35277));
    LocalMux I__7475 (
            .O(N__35280),
            .I(data_out_0_3));
    Odrv4 I__7474 (
            .O(N__35277),
            .I(data_out_0_3));
    InMux I__7473 (
            .O(N__35272),
            .I(N__35268));
    InMux I__7472 (
            .O(N__35271),
            .I(N__35265));
    LocalMux I__7471 (
            .O(N__35268),
            .I(data_out_2_2));
    LocalMux I__7470 (
            .O(N__35265),
            .I(data_out_2_2));
    InMux I__7469 (
            .O(N__35260),
            .I(N__35257));
    LocalMux I__7468 (
            .O(N__35257),
            .I(N__35254));
    Span4Mux_v I__7467 (
            .O(N__35254),
            .I(N__35251));
    Odrv4 I__7466 (
            .O(N__35251),
            .I(\c0.n2_adj_2291 ));
    InMux I__7465 (
            .O(N__35248),
            .I(N__35242));
    InMux I__7464 (
            .O(N__35247),
            .I(N__35242));
    LocalMux I__7463 (
            .O(N__35242),
            .I(data_out_3_2));
    CascadeMux I__7462 (
            .O(N__35239),
            .I(N__35233));
    InMux I__7461 (
            .O(N__35238),
            .I(N__35227));
    InMux I__7460 (
            .O(N__35237),
            .I(N__35227));
    InMux I__7459 (
            .O(N__35236),
            .I(N__35224));
    InMux I__7458 (
            .O(N__35233),
            .I(N__35219));
    InMux I__7457 (
            .O(N__35232),
            .I(N__35219));
    LocalMux I__7456 (
            .O(N__35227),
            .I(N__35216));
    LocalMux I__7455 (
            .O(N__35224),
            .I(N__35212));
    LocalMux I__7454 (
            .O(N__35219),
            .I(N__35209));
    Span4Mux_v I__7453 (
            .O(N__35216),
            .I(N__35206));
    InMux I__7452 (
            .O(N__35215),
            .I(N__35203));
    Span4Mux_h I__7451 (
            .O(N__35212),
            .I(N__35200));
    Span4Mux_v I__7450 (
            .O(N__35209),
            .I(N__35197));
    Span4Mux_h I__7449 (
            .O(N__35206),
            .I(N__35194));
    LocalMux I__7448 (
            .O(N__35203),
            .I(data_out_frame2_9_4));
    Odrv4 I__7447 (
            .O(N__35200),
            .I(data_out_frame2_9_4));
    Odrv4 I__7446 (
            .O(N__35197),
            .I(data_out_frame2_9_4));
    Odrv4 I__7445 (
            .O(N__35194),
            .I(data_out_frame2_9_4));
    InMux I__7444 (
            .O(N__35185),
            .I(N__35182));
    LocalMux I__7443 (
            .O(N__35182),
            .I(N__35179));
    Sp12to4 I__7442 (
            .O(N__35179),
            .I(N__35176));
    Odrv12 I__7441 (
            .O(N__35176),
            .I(\c0.n9_adj_2347 ));
    InMux I__7440 (
            .O(N__35173),
            .I(N__35170));
    LocalMux I__7439 (
            .O(N__35170),
            .I(\c0.n17897 ));
    InMux I__7438 (
            .O(N__35167),
            .I(N__35160));
    InMux I__7437 (
            .O(N__35166),
            .I(N__35160));
    InMux I__7436 (
            .O(N__35165),
            .I(N__35156));
    LocalMux I__7435 (
            .O(N__35160),
            .I(N__35153));
    InMux I__7434 (
            .O(N__35159),
            .I(N__35150));
    LocalMux I__7433 (
            .O(N__35156),
            .I(data_out_frame2_10_2));
    Odrv4 I__7432 (
            .O(N__35153),
            .I(data_out_frame2_10_2));
    LocalMux I__7431 (
            .O(N__35150),
            .I(data_out_frame2_10_2));
    InMux I__7430 (
            .O(N__35143),
            .I(N__35140));
    LocalMux I__7429 (
            .O(N__35140),
            .I(N__35137));
    Odrv4 I__7428 (
            .O(N__35137),
            .I(\c0.n12_adj_2305 ));
    InMux I__7427 (
            .O(N__35134),
            .I(N__35131));
    LocalMux I__7426 (
            .O(N__35131),
            .I(\c0.n17990 ));
    CascadeMux I__7425 (
            .O(N__35128),
            .I(\c0.n17993_cascade_ ));
    InMux I__7424 (
            .O(N__35125),
            .I(N__35122));
    LocalMux I__7423 (
            .O(N__35122),
            .I(\c0.n17894 ));
    CascadeMux I__7422 (
            .O(N__35119),
            .I(\c0.n17393_cascade_ ));
    InMux I__7421 (
            .O(N__35116),
            .I(N__35113));
    LocalMux I__7420 (
            .O(N__35113),
            .I(N__35110));
    Odrv4 I__7419 (
            .O(N__35110),
            .I(\c0.n17571 ));
    CascadeMux I__7418 (
            .O(N__35107),
            .I(\c0.n17963_cascade_ ));
    CascadeMux I__7417 (
            .O(N__35104),
            .I(\c0.n17966_cascade_ ));
    InMux I__7416 (
            .O(N__35101),
            .I(N__35098));
    LocalMux I__7415 (
            .O(N__35098),
            .I(N__35095));
    Span4Mux_v I__7414 (
            .O(N__35095),
            .I(N__35092));
    Odrv4 I__7413 (
            .O(N__35092),
            .I(\c0.tx2.r_Tx_Data_5 ));
    InMux I__7412 (
            .O(N__35089),
            .I(N__35086));
    LocalMux I__7411 (
            .O(N__35086),
            .I(N__35082));
    InMux I__7410 (
            .O(N__35085),
            .I(N__35079));
    Span4Mux_v I__7409 (
            .O(N__35082),
            .I(N__35076));
    LocalMux I__7408 (
            .O(N__35079),
            .I(data_out_0_5));
    Odrv4 I__7407 (
            .O(N__35076),
            .I(data_out_0_5));
    CascadeMux I__7406 (
            .O(N__35071),
            .I(N__35068));
    InMux I__7405 (
            .O(N__35068),
            .I(N__35065));
    LocalMux I__7404 (
            .O(N__35065),
            .I(N__35059));
    InMux I__7403 (
            .O(N__35064),
            .I(N__35056));
    InMux I__7402 (
            .O(N__35063),
            .I(N__35053));
    InMux I__7401 (
            .O(N__35062),
            .I(N__35050));
    Span4Mux_h I__7400 (
            .O(N__35059),
            .I(N__35047));
    LocalMux I__7399 (
            .O(N__35056),
            .I(data_out_frame2_5_3));
    LocalMux I__7398 (
            .O(N__35053),
            .I(data_out_frame2_5_3));
    LocalMux I__7397 (
            .O(N__35050),
            .I(data_out_frame2_5_3));
    Odrv4 I__7396 (
            .O(N__35047),
            .I(data_out_frame2_5_3));
    InMux I__7395 (
            .O(N__35038),
            .I(N__35031));
    InMux I__7394 (
            .O(N__35037),
            .I(N__35028));
    InMux I__7393 (
            .O(N__35036),
            .I(N__35025));
    InMux I__7392 (
            .O(N__35035),
            .I(N__35022));
    InMux I__7391 (
            .O(N__35034),
            .I(N__35019));
    LocalMux I__7390 (
            .O(N__35031),
            .I(N__35014));
    LocalMux I__7389 (
            .O(N__35028),
            .I(N__35005));
    LocalMux I__7388 (
            .O(N__35025),
            .I(N__35005));
    LocalMux I__7387 (
            .O(N__35022),
            .I(N__35005));
    LocalMux I__7386 (
            .O(N__35019),
            .I(N__35005));
    InMux I__7385 (
            .O(N__35018),
            .I(N__35001));
    InMux I__7384 (
            .O(N__35017),
            .I(N__34998));
    Span4Mux_h I__7383 (
            .O(N__35014),
            .I(N__34993));
    Span4Mux_v I__7382 (
            .O(N__35005),
            .I(N__34993));
    InMux I__7381 (
            .O(N__35004),
            .I(N__34990));
    LocalMux I__7380 (
            .O(N__35001),
            .I(\c0.n16148 ));
    LocalMux I__7379 (
            .O(N__34998),
            .I(\c0.n16148 ));
    Odrv4 I__7378 (
            .O(N__34993),
            .I(\c0.n16148 ));
    LocalMux I__7377 (
            .O(N__34990),
            .I(\c0.n16148 ));
    CascadeMux I__7376 (
            .O(N__34981),
            .I(\c0.n17331_cascade_ ));
    InMux I__7375 (
            .O(N__34978),
            .I(N__34973));
    InMux I__7374 (
            .O(N__34977),
            .I(N__34970));
    InMux I__7373 (
            .O(N__34976),
            .I(N__34967));
    LocalMux I__7372 (
            .O(N__34973),
            .I(N__34964));
    LocalMux I__7371 (
            .O(N__34970),
            .I(N__34961));
    LocalMux I__7370 (
            .O(N__34967),
            .I(N__34958));
    Span4Mux_v I__7369 (
            .O(N__34964),
            .I(N__34953));
    Span4Mux_h I__7368 (
            .O(N__34961),
            .I(N__34950));
    Span4Mux_h I__7367 (
            .O(N__34958),
            .I(N__34947));
    InMux I__7366 (
            .O(N__34957),
            .I(N__34944));
    InMux I__7365 (
            .O(N__34956),
            .I(N__34941));
    Odrv4 I__7364 (
            .O(N__34953),
            .I(\c0.n15846 ));
    Odrv4 I__7363 (
            .O(N__34950),
            .I(\c0.n15846 ));
    Odrv4 I__7362 (
            .O(N__34947),
            .I(\c0.n15846 ));
    LocalMux I__7361 (
            .O(N__34944),
            .I(\c0.n15846 ));
    LocalMux I__7360 (
            .O(N__34941),
            .I(\c0.n15846 ));
    InMux I__7359 (
            .O(N__34930),
            .I(N__34927));
    LocalMux I__7358 (
            .O(N__34927),
            .I(\c0.n17891 ));
    InMux I__7357 (
            .O(N__34924),
            .I(N__34921));
    LocalMux I__7356 (
            .O(N__34921),
            .I(N__34918));
    Odrv4 I__7355 (
            .O(N__34918),
            .I(\c0.n17939 ));
    InMux I__7354 (
            .O(N__34915),
            .I(N__34909));
    InMux I__7353 (
            .O(N__34914),
            .I(N__34906));
    InMux I__7352 (
            .O(N__34913),
            .I(N__34903));
    InMux I__7351 (
            .O(N__34912),
            .I(N__34900));
    LocalMux I__7350 (
            .O(N__34909),
            .I(data_out_frame2_6_3));
    LocalMux I__7349 (
            .O(N__34906),
            .I(data_out_frame2_6_3));
    LocalMux I__7348 (
            .O(N__34903),
            .I(data_out_frame2_6_3));
    LocalMux I__7347 (
            .O(N__34900),
            .I(data_out_frame2_6_3));
    CascadeMux I__7346 (
            .O(N__34891),
            .I(N__34888));
    InMux I__7345 (
            .O(N__34888),
            .I(N__34885));
    LocalMux I__7344 (
            .O(N__34885),
            .I(N__34882));
    Span4Mux_v I__7343 (
            .O(N__34882),
            .I(N__34879));
    Odrv4 I__7342 (
            .O(N__34879),
            .I(\c0.n16_adj_2197 ));
    InMux I__7341 (
            .O(N__34876),
            .I(N__34873));
    LocalMux I__7340 (
            .O(N__34873),
            .I(N__34870));
    Odrv4 I__7339 (
            .O(N__34870),
            .I(\c0.n22_adj_2194 ));
    InMux I__7338 (
            .O(N__34867),
            .I(N__34864));
    LocalMux I__7337 (
            .O(N__34864),
            .I(N__34861));
    Odrv4 I__7336 (
            .O(N__34861),
            .I(\c0.n9754 ));
    CascadeMux I__7335 (
            .O(N__34858),
            .I(\c0.n9901_cascade_ ));
    InMux I__7334 (
            .O(N__34855),
            .I(N__34852));
    LocalMux I__7333 (
            .O(N__34852),
            .I(\c0.n6_adj_2201 ));
    InMux I__7332 (
            .O(N__34849),
            .I(N__34846));
    LocalMux I__7331 (
            .O(N__34846),
            .I(\c0.n17942 ));
    CascadeMux I__7330 (
            .O(N__34843),
            .I(N__34840));
    InMux I__7329 (
            .O(N__34840),
            .I(N__34837));
    LocalMux I__7328 (
            .O(N__34837),
            .I(N__34834));
    Span4Mux_h I__7327 (
            .O(N__34834),
            .I(N__34831));
    Odrv4 I__7326 (
            .O(N__34831),
            .I(\c0.n17560 ));
    CascadeMux I__7325 (
            .O(N__34828),
            .I(\c0.n17301_cascade_ ));
    CascadeMux I__7324 (
            .O(N__34825),
            .I(\c0.n17303_cascade_ ));
    InMux I__7323 (
            .O(N__34822),
            .I(N__34819));
    LocalMux I__7322 (
            .O(N__34819),
            .I(N__34816));
    Span4Mux_h I__7321 (
            .O(N__34816),
            .I(N__34813));
    Span4Mux_v I__7320 (
            .O(N__34813),
            .I(N__34810));
    Odrv4 I__7319 (
            .O(N__34810),
            .I(\c0.tx2.r_Tx_Data_0 ));
    InMux I__7318 (
            .O(N__34807),
            .I(N__34803));
    InMux I__7317 (
            .O(N__34806),
            .I(N__34800));
    LocalMux I__7316 (
            .O(N__34803),
            .I(N__34797));
    LocalMux I__7315 (
            .O(N__34800),
            .I(data_out_frame2_18_0));
    Odrv4 I__7314 (
            .O(N__34797),
            .I(data_out_frame2_18_0));
    InMux I__7313 (
            .O(N__34792),
            .I(N__34789));
    LocalMux I__7312 (
            .O(N__34789),
            .I(N__34786));
    Span4Mux_v I__7311 (
            .O(N__34786),
            .I(N__34782));
    InMux I__7310 (
            .O(N__34785),
            .I(N__34779));
    Span4Mux_h I__7309 (
            .O(N__34782),
            .I(N__34776));
    LocalMux I__7308 (
            .O(N__34779),
            .I(data_out_frame2_17_0));
    Odrv4 I__7307 (
            .O(N__34776),
            .I(data_out_frame2_17_0));
    CascadeMux I__7306 (
            .O(N__34771),
            .I(\c0.n18101_cascade_ ));
    CascadeMux I__7305 (
            .O(N__34768),
            .I(\c0.n18104_cascade_ ));
    InMux I__7304 (
            .O(N__34765),
            .I(N__34762));
    LocalMux I__7303 (
            .O(N__34762),
            .I(\c0.n22_adj_2337 ));
    InMux I__7302 (
            .O(N__34759),
            .I(\c0.n15618 ));
    InMux I__7301 (
            .O(N__34756),
            .I(N__34753));
    LocalMux I__7300 (
            .O(N__34753),
            .I(N__34749));
    InMux I__7299 (
            .O(N__34752),
            .I(N__34746));
    Span4Mux_h I__7298 (
            .O(N__34749),
            .I(N__34743));
    LocalMux I__7297 (
            .O(N__34746),
            .I(\c0.byte_transmit_counter2_5 ));
    Odrv4 I__7296 (
            .O(N__34743),
            .I(\c0.byte_transmit_counter2_5 ));
    InMux I__7295 (
            .O(N__34738),
            .I(\c0.n15619 ));
    CascadeMux I__7294 (
            .O(N__34735),
            .I(N__34732));
    InMux I__7293 (
            .O(N__34732),
            .I(N__34729));
    LocalMux I__7292 (
            .O(N__34729),
            .I(N__34725));
    InMux I__7291 (
            .O(N__34728),
            .I(N__34722));
    Span4Mux_h I__7290 (
            .O(N__34725),
            .I(N__34719));
    LocalMux I__7289 (
            .O(N__34722),
            .I(\c0.byte_transmit_counter2_6 ));
    Odrv4 I__7288 (
            .O(N__34719),
            .I(\c0.byte_transmit_counter2_6 ));
    InMux I__7287 (
            .O(N__34714),
            .I(\c0.n15620 ));
    InMux I__7286 (
            .O(N__34711),
            .I(\c0.n15621 ));
    InMux I__7285 (
            .O(N__34708),
            .I(N__34705));
    LocalMux I__7284 (
            .O(N__34705),
            .I(N__34701));
    InMux I__7283 (
            .O(N__34704),
            .I(N__34698));
    Span4Mux_h I__7282 (
            .O(N__34701),
            .I(N__34695));
    LocalMux I__7281 (
            .O(N__34698),
            .I(\c0.byte_transmit_counter2_7 ));
    Odrv4 I__7280 (
            .O(N__34695),
            .I(\c0.byte_transmit_counter2_7 ));
    CEMux I__7279 (
            .O(N__34690),
            .I(N__34687));
    LocalMux I__7278 (
            .O(N__34687),
            .I(N__34684));
    Span4Mux_h I__7277 (
            .O(N__34684),
            .I(N__34680));
    InMux I__7276 (
            .O(N__34683),
            .I(N__34677));
    Odrv4 I__7275 (
            .O(N__34680),
            .I(\c0.n10052 ));
    LocalMux I__7274 (
            .O(N__34677),
            .I(\c0.n10052 ));
    SRMux I__7273 (
            .O(N__34672),
            .I(N__34669));
    LocalMux I__7272 (
            .O(N__34669),
            .I(N__34666));
    Odrv12 I__7271 (
            .O(N__34666),
            .I(\c0.n10297 ));
    InMux I__7270 (
            .O(N__34663),
            .I(N__34656));
    InMux I__7269 (
            .O(N__34662),
            .I(N__34638));
    InMux I__7268 (
            .O(N__34661),
            .I(N__34635));
    InMux I__7267 (
            .O(N__34660),
            .I(N__34632));
    InMux I__7266 (
            .O(N__34659),
            .I(N__34629));
    LocalMux I__7265 (
            .O(N__34656),
            .I(N__34626));
    InMux I__7264 (
            .O(N__34655),
            .I(N__34623));
    InMux I__7263 (
            .O(N__34654),
            .I(N__34620));
    InMux I__7262 (
            .O(N__34653),
            .I(N__34617));
    InMux I__7261 (
            .O(N__34652),
            .I(N__34614));
    InMux I__7260 (
            .O(N__34651),
            .I(N__34610));
    InMux I__7259 (
            .O(N__34650),
            .I(N__34607));
    InMux I__7258 (
            .O(N__34649),
            .I(N__34604));
    InMux I__7257 (
            .O(N__34648),
            .I(N__34601));
    InMux I__7256 (
            .O(N__34647),
            .I(N__34598));
    InMux I__7255 (
            .O(N__34646),
            .I(N__34595));
    InMux I__7254 (
            .O(N__34645),
            .I(N__34592));
    InMux I__7253 (
            .O(N__34644),
            .I(N__34589));
    InMux I__7252 (
            .O(N__34643),
            .I(N__34586));
    InMux I__7251 (
            .O(N__34642),
            .I(N__34583));
    InMux I__7250 (
            .O(N__34641),
            .I(N__34580));
    LocalMux I__7249 (
            .O(N__34638),
            .I(N__34577));
    LocalMux I__7248 (
            .O(N__34635),
            .I(N__34574));
    LocalMux I__7247 (
            .O(N__34632),
            .I(N__34565));
    LocalMux I__7246 (
            .O(N__34629),
            .I(N__34565));
    Span4Mux_s1_h I__7245 (
            .O(N__34626),
            .I(N__34565));
    LocalMux I__7244 (
            .O(N__34623),
            .I(N__34565));
    LocalMux I__7243 (
            .O(N__34620),
            .I(N__34555));
    LocalMux I__7242 (
            .O(N__34617),
            .I(N__34550));
    LocalMux I__7241 (
            .O(N__34614),
            .I(N__34550));
    InMux I__7240 (
            .O(N__34613),
            .I(N__34547));
    LocalMux I__7239 (
            .O(N__34610),
            .I(N__34544));
    LocalMux I__7238 (
            .O(N__34607),
            .I(N__34537));
    LocalMux I__7237 (
            .O(N__34604),
            .I(N__34537));
    LocalMux I__7236 (
            .O(N__34601),
            .I(N__34537));
    LocalMux I__7235 (
            .O(N__34598),
            .I(N__34530));
    LocalMux I__7234 (
            .O(N__34595),
            .I(N__34530));
    LocalMux I__7233 (
            .O(N__34592),
            .I(N__34530));
    LocalMux I__7232 (
            .O(N__34589),
            .I(N__34527));
    LocalMux I__7231 (
            .O(N__34586),
            .I(N__34524));
    LocalMux I__7230 (
            .O(N__34583),
            .I(N__34521));
    LocalMux I__7229 (
            .O(N__34580),
            .I(N__34516));
    Span4Mux_v I__7228 (
            .O(N__34577),
            .I(N__34516));
    Span4Mux_v I__7227 (
            .O(N__34574),
            .I(N__34511));
    Span4Mux_v I__7226 (
            .O(N__34565),
            .I(N__34511));
    InMux I__7225 (
            .O(N__34564),
            .I(N__34508));
    InMux I__7224 (
            .O(N__34563),
            .I(N__34505));
    InMux I__7223 (
            .O(N__34562),
            .I(N__34502));
    InMux I__7222 (
            .O(N__34561),
            .I(N__34499));
    InMux I__7221 (
            .O(N__34560),
            .I(N__34496));
    InMux I__7220 (
            .O(N__34559),
            .I(N__34493));
    InMux I__7219 (
            .O(N__34558),
            .I(N__34490));
    Span4Mux_h I__7218 (
            .O(N__34555),
            .I(N__34485));
    Span4Mux_v I__7217 (
            .O(N__34550),
            .I(N__34485));
    LocalMux I__7216 (
            .O(N__34547),
            .I(N__34476));
    Span4Mux_h I__7215 (
            .O(N__34544),
            .I(N__34476));
    Span4Mux_v I__7214 (
            .O(N__34537),
            .I(N__34476));
    Span4Mux_v I__7213 (
            .O(N__34530),
            .I(N__34476));
    Span4Mux_v I__7212 (
            .O(N__34527),
            .I(N__34467));
    Span4Mux_v I__7211 (
            .O(N__34524),
            .I(N__34467));
    Span4Mux_v I__7210 (
            .O(N__34521),
            .I(N__34467));
    Span4Mux_h I__7209 (
            .O(N__34516),
            .I(N__34467));
    Span4Mux_h I__7208 (
            .O(N__34511),
            .I(N__34464));
    LocalMux I__7207 (
            .O(N__34508),
            .I(\c0.n7 ));
    LocalMux I__7206 (
            .O(N__34505),
            .I(\c0.n7 ));
    LocalMux I__7205 (
            .O(N__34502),
            .I(\c0.n7 ));
    LocalMux I__7204 (
            .O(N__34499),
            .I(\c0.n7 ));
    LocalMux I__7203 (
            .O(N__34496),
            .I(\c0.n7 ));
    LocalMux I__7202 (
            .O(N__34493),
            .I(\c0.n7 ));
    LocalMux I__7201 (
            .O(N__34490),
            .I(\c0.n7 ));
    Odrv4 I__7200 (
            .O(N__34485),
            .I(\c0.n7 ));
    Odrv4 I__7199 (
            .O(N__34476),
            .I(\c0.n7 ));
    Odrv4 I__7198 (
            .O(N__34467),
            .I(\c0.n7 ));
    Odrv4 I__7197 (
            .O(N__34464),
            .I(\c0.n7 ));
    CascadeMux I__7196 (
            .O(N__34441),
            .I(N__34438));
    InMux I__7195 (
            .O(N__34438),
            .I(N__34435));
    LocalMux I__7194 (
            .O(N__34435),
            .I(N__34432));
    Span4Mux_h I__7193 (
            .O(N__34432),
            .I(N__34427));
    InMux I__7192 (
            .O(N__34431),
            .I(N__34424));
    InMux I__7191 (
            .O(N__34430),
            .I(N__34421));
    Span4Mux_h I__7190 (
            .O(N__34427),
            .I(N__34418));
    LocalMux I__7189 (
            .O(N__34424),
            .I(\c0.FRAME_MATCHER_state_9 ));
    LocalMux I__7188 (
            .O(N__34421),
            .I(\c0.FRAME_MATCHER_state_9 ));
    Odrv4 I__7187 (
            .O(N__34418),
            .I(\c0.FRAME_MATCHER_state_9 ));
    SRMux I__7186 (
            .O(N__34411),
            .I(N__34408));
    LocalMux I__7185 (
            .O(N__34408),
            .I(\c0.n16455 ));
    InMux I__7184 (
            .O(N__34405),
            .I(N__34402));
    LocalMux I__7183 (
            .O(N__34402),
            .I(\c0.n17927 ));
    CascadeMux I__7182 (
            .O(N__34399),
            .I(N__34396));
    InMux I__7181 (
            .O(N__34396),
            .I(N__34393));
    LocalMux I__7180 (
            .O(N__34393),
            .I(N__34389));
    InMux I__7179 (
            .O(N__34392),
            .I(N__34386));
    Span4Mux_v I__7178 (
            .O(N__34389),
            .I(N__34383));
    LocalMux I__7177 (
            .O(N__34386),
            .I(data_out_frame2_17_2));
    Odrv4 I__7176 (
            .O(N__34383),
            .I(data_out_frame2_17_2));
    CascadeMux I__7175 (
            .O(N__34378),
            .I(\c0.n17930_cascade_ ));
    InMux I__7174 (
            .O(N__34375),
            .I(N__34372));
    LocalMux I__7173 (
            .O(N__34372),
            .I(\c0.n22_adj_2358 ));
    CascadeMux I__7172 (
            .O(N__34369),
            .I(N__34366));
    InMux I__7171 (
            .O(N__34366),
            .I(N__34363));
    LocalMux I__7170 (
            .O(N__34363),
            .I(\c0.n17936 ));
    CascadeMux I__7169 (
            .O(N__34360),
            .I(\c0.n17456_cascade_ ));
    CEMux I__7168 (
            .O(N__34357),
            .I(N__34352));
    CascadeMux I__7167 (
            .O(N__34356),
            .I(N__34349));
    InMux I__7166 (
            .O(N__34355),
            .I(N__34345));
    LocalMux I__7165 (
            .O(N__34352),
            .I(N__34342));
    InMux I__7164 (
            .O(N__34349),
            .I(N__34339));
    InMux I__7163 (
            .O(N__34348),
            .I(N__34336));
    LocalMux I__7162 (
            .O(N__34345),
            .I(N__34333));
    Span4Mux_s2_v I__7161 (
            .O(N__34342),
            .I(N__34330));
    LocalMux I__7160 (
            .O(N__34339),
            .I(\c0.n10054 ));
    LocalMux I__7159 (
            .O(N__34336),
            .I(\c0.n10054 ));
    Odrv4 I__7158 (
            .O(N__34333),
            .I(\c0.n10054 ));
    Odrv4 I__7157 (
            .O(N__34330),
            .I(\c0.n10054 ));
    InMux I__7156 (
            .O(N__34321),
            .I(N__34318));
    LocalMux I__7155 (
            .O(N__34318),
            .I(N__34314));
    InMux I__7154 (
            .O(N__34317),
            .I(N__34311));
    Span4Mux_h I__7153 (
            .O(N__34314),
            .I(N__34304));
    LocalMux I__7152 (
            .O(N__34311),
            .I(N__34304));
    InMux I__7151 (
            .O(N__34310),
            .I(N__34299));
    InMux I__7150 (
            .O(N__34309),
            .I(N__34299));
    Span4Mux_h I__7149 (
            .O(N__34304),
            .I(N__34294));
    LocalMux I__7148 (
            .O(N__34299),
            .I(N__34294));
    Odrv4 I__7147 (
            .O(N__34294),
            .I(n9361));
    InMux I__7146 (
            .O(N__34291),
            .I(N__34288));
    LocalMux I__7145 (
            .O(N__34288),
            .I(N__34285));
    Odrv12 I__7144 (
            .O(N__34285),
            .I(n17154));
    InMux I__7143 (
            .O(N__34282),
            .I(N__34277));
    InMux I__7142 (
            .O(N__34281),
            .I(N__34272));
    InMux I__7141 (
            .O(N__34280),
            .I(N__34269));
    LocalMux I__7140 (
            .O(N__34277),
            .I(N__34266));
    InMux I__7139 (
            .O(N__34276),
            .I(N__34263));
    InMux I__7138 (
            .O(N__34275),
            .I(N__34259));
    LocalMux I__7137 (
            .O(N__34272),
            .I(N__34256));
    LocalMux I__7136 (
            .O(N__34269),
            .I(N__34249));
    Span4Mux_v I__7135 (
            .O(N__34266),
            .I(N__34249));
    LocalMux I__7134 (
            .O(N__34263),
            .I(N__34249));
    InMux I__7133 (
            .O(N__34262),
            .I(N__34243));
    LocalMux I__7132 (
            .O(N__34259),
            .I(N__34238));
    Span12Mux_v I__7131 (
            .O(N__34256),
            .I(N__34238));
    Span4Mux_v I__7130 (
            .O(N__34249),
            .I(N__34235));
    InMux I__7129 (
            .O(N__34248),
            .I(N__34228));
    InMux I__7128 (
            .O(N__34247),
            .I(N__34228));
    InMux I__7127 (
            .O(N__34246),
            .I(N__34228));
    LocalMux I__7126 (
            .O(N__34243),
            .I(FRAME_MATCHER_state_0));
    Odrv12 I__7125 (
            .O(N__34238),
            .I(FRAME_MATCHER_state_0));
    Odrv4 I__7124 (
            .O(N__34235),
            .I(FRAME_MATCHER_state_0));
    LocalMux I__7123 (
            .O(N__34228),
            .I(FRAME_MATCHER_state_0));
    InMux I__7122 (
            .O(N__34219),
            .I(N__34216));
    LocalMux I__7121 (
            .O(N__34216),
            .I(N__34213));
    Span4Mux_h I__7120 (
            .O(N__34213),
            .I(N__34210));
    Odrv4 I__7119 (
            .O(N__34210),
            .I(\c0.tx2_transmit_N_1997 ));
    InMux I__7118 (
            .O(N__34207),
            .I(\c0.n15615 ));
    InMux I__7117 (
            .O(N__34204),
            .I(\c0.n15616 ));
    InMux I__7116 (
            .O(N__34201),
            .I(\c0.n15617 ));
    InMux I__7115 (
            .O(N__34198),
            .I(N__34189));
    InMux I__7114 (
            .O(N__34197),
            .I(N__34189));
    InMux I__7113 (
            .O(N__34196),
            .I(N__34186));
    InMux I__7112 (
            .O(N__34195),
            .I(N__34181));
    InMux I__7111 (
            .O(N__34194),
            .I(N__34181));
    LocalMux I__7110 (
            .O(N__34189),
            .I(N__34176));
    LocalMux I__7109 (
            .O(N__34186),
            .I(N__34176));
    LocalMux I__7108 (
            .O(N__34181),
            .I(\c0.data_out_7_7 ));
    Odrv4 I__7107 (
            .O(N__34176),
            .I(\c0.data_out_7_7 ));
    CascadeMux I__7106 (
            .O(N__34171),
            .I(\c0.n5_adj_2188_cascade_ ));
    InMux I__7105 (
            .O(N__34168),
            .I(N__34165));
    LocalMux I__7104 (
            .O(N__34165),
            .I(\c0.n18041 ));
    InMux I__7103 (
            .O(N__34162),
            .I(N__34159));
    LocalMux I__7102 (
            .O(N__34159),
            .I(\c0.n5_adj_2208 ));
    CascadeMux I__7101 (
            .O(N__34156),
            .I(\c0.n17543_cascade_ ));
    InMux I__7100 (
            .O(N__34153),
            .I(N__34150));
    LocalMux I__7099 (
            .O(N__34150),
            .I(\c0.n18011 ));
    InMux I__7098 (
            .O(N__34147),
            .I(N__34144));
    LocalMux I__7097 (
            .O(N__34144),
            .I(\c0.n17445 ));
    InMux I__7096 (
            .O(N__34141),
            .I(N__34137));
    CascadeMux I__7095 (
            .O(N__34140),
            .I(N__34134));
    LocalMux I__7094 (
            .O(N__34137),
            .I(N__34130));
    InMux I__7093 (
            .O(N__34134),
            .I(N__34127));
    InMux I__7092 (
            .O(N__34133),
            .I(N__34124));
    Span4Mux_h I__7091 (
            .O(N__34130),
            .I(N__34121));
    LocalMux I__7090 (
            .O(N__34127),
            .I(\c0.data_out_7_5 ));
    LocalMux I__7089 (
            .O(N__34124),
            .I(\c0.data_out_7_5 ));
    Odrv4 I__7088 (
            .O(N__34121),
            .I(\c0.data_out_7_5 ));
    CascadeMux I__7087 (
            .O(N__34114),
            .I(N__34111));
    InMux I__7086 (
            .O(N__34111),
            .I(N__34108));
    LocalMux I__7085 (
            .O(N__34108),
            .I(N__34105));
    Odrv4 I__7084 (
            .O(N__34105),
            .I(\c0.n26 ));
    InMux I__7083 (
            .O(N__34102),
            .I(N__34099));
    LocalMux I__7082 (
            .O(N__34099),
            .I(N__34096));
    Odrv12 I__7081 (
            .O(N__34096),
            .I(n18032));
    InMux I__7080 (
            .O(N__34093),
            .I(N__34090));
    LocalMux I__7079 (
            .O(N__34090),
            .I(n10));
    CascadeMux I__7078 (
            .O(N__34087),
            .I(N__34084));
    InMux I__7077 (
            .O(N__34084),
            .I(N__34081));
    LocalMux I__7076 (
            .O(N__34081),
            .I(N__34078));
    Odrv4 I__7075 (
            .O(N__34078),
            .I(\c0.n5_adj_2142 ));
    InMux I__7074 (
            .O(N__34075),
            .I(N__34071));
    InMux I__7073 (
            .O(N__34074),
            .I(N__34068));
    LocalMux I__7072 (
            .O(N__34071),
            .I(N__34065));
    LocalMux I__7071 (
            .O(N__34068),
            .I(data_out_3_0));
    Odrv4 I__7070 (
            .O(N__34065),
            .I(data_out_3_0));
    InMux I__7069 (
            .O(N__34060),
            .I(N__34057));
    LocalMux I__7068 (
            .O(N__34057),
            .I(N__34054));
    Span4Mux_v I__7067 (
            .O(N__34054),
            .I(N__34050));
    InMux I__7066 (
            .O(N__34053),
            .I(N__34047));
    Span4Mux_h I__7065 (
            .O(N__34050),
            .I(N__34044));
    LocalMux I__7064 (
            .O(N__34047),
            .I(\c0.data_out_3_6 ));
    Odrv4 I__7063 (
            .O(N__34044),
            .I(\c0.data_out_3_6 ));
    CascadeMux I__7062 (
            .O(N__34039),
            .I(\c0.n10054_cascade_ ));
    InMux I__7061 (
            .O(N__34036),
            .I(N__34032));
    InMux I__7060 (
            .O(N__34035),
            .I(N__34029));
    LocalMux I__7059 (
            .O(N__34032),
            .I(data_out_3_5));
    LocalMux I__7058 (
            .O(N__34029),
            .I(data_out_3_5));
    CascadeMux I__7057 (
            .O(N__34024),
            .I(N__34021));
    InMux I__7056 (
            .O(N__34021),
            .I(N__34017));
    InMux I__7055 (
            .O(N__34020),
            .I(N__34014));
    LocalMux I__7054 (
            .O(N__34017),
            .I(data_out_2_5));
    LocalMux I__7053 (
            .O(N__34014),
            .I(data_out_2_5));
    CascadeMux I__7052 (
            .O(N__34009),
            .I(N__34006));
    InMux I__7051 (
            .O(N__34006),
            .I(N__34003));
    LocalMux I__7050 (
            .O(N__34003),
            .I(N__34000));
    Span4Mux_h I__7049 (
            .O(N__34000),
            .I(N__33997));
    Span4Mux_h I__7048 (
            .O(N__33997),
            .I(N__33994));
    Odrv4 I__7047 (
            .O(N__33994),
            .I(\c0.n9530 ));
    CascadeMux I__7046 (
            .O(N__33991),
            .I(N__33988));
    InMux I__7045 (
            .O(N__33988),
            .I(N__33984));
    InMux I__7044 (
            .O(N__33987),
            .I(N__33981));
    LocalMux I__7043 (
            .O(N__33984),
            .I(data_out_1_6));
    LocalMux I__7042 (
            .O(N__33981),
            .I(data_out_1_6));
    InMux I__7041 (
            .O(N__33976),
            .I(N__33973));
    LocalMux I__7040 (
            .O(N__33973),
            .I(N__33969));
    InMux I__7039 (
            .O(N__33972),
            .I(N__33966));
    Span4Mux_h I__7038 (
            .O(N__33969),
            .I(N__33963));
    LocalMux I__7037 (
            .O(N__33966),
            .I(data_out_2_0));
    Odrv4 I__7036 (
            .O(N__33963),
            .I(data_out_2_0));
    InMux I__7035 (
            .O(N__33958),
            .I(N__33955));
    LocalMux I__7034 (
            .O(N__33955),
            .I(N__33952));
    Odrv12 I__7033 (
            .O(N__33952),
            .I(\c0.n9509 ));
    InMux I__7032 (
            .O(N__33949),
            .I(N__33946));
    LocalMux I__7031 (
            .O(N__33946),
            .I(N__33943));
    Span4Mux_h I__7030 (
            .O(N__33943),
            .I(N__33940));
    Odrv4 I__7029 (
            .O(N__33940),
            .I(\c0.tx2.r_Tx_Data_1 ));
    InMux I__7028 (
            .O(N__33937),
            .I(N__33934));
    LocalMux I__7027 (
            .O(N__33934),
            .I(N__33931));
    Span4Mux_v I__7026 (
            .O(N__33931),
            .I(N__33928));
    Odrv4 I__7025 (
            .O(N__33928),
            .I(\c0.n17548 ));
    InMux I__7024 (
            .O(N__33925),
            .I(N__33922));
    LocalMux I__7023 (
            .O(N__33922),
            .I(N__33919));
    Odrv12 I__7022 (
            .O(N__33919),
            .I(\c0.n17589 ));
    InMux I__7021 (
            .O(N__33916),
            .I(N__33913));
    LocalMux I__7020 (
            .O(N__33913),
            .I(N__33910));
    Odrv4 I__7019 (
            .O(N__33910),
            .I(\c0.n2_adj_2298 ));
    CascadeMux I__7018 (
            .O(N__33907),
            .I(\c0.n18029_cascade_ ));
    InMux I__7017 (
            .O(N__33904),
            .I(N__33901));
    LocalMux I__7016 (
            .O(N__33901),
            .I(N__33898));
    Odrv4 I__7015 (
            .O(N__33898),
            .I(\c0.n8_adj_2138 ));
    CascadeMux I__7014 (
            .O(N__33895),
            .I(N__33892));
    InMux I__7013 (
            .O(N__33892),
            .I(N__33889));
    LocalMux I__7012 (
            .O(N__33889),
            .I(\c0.n5_adj_2299 ));
    CascadeMux I__7011 (
            .O(N__33886),
            .I(N__33882));
    CascadeMux I__7010 (
            .O(N__33885),
            .I(N__33877));
    InMux I__7009 (
            .O(N__33882),
            .I(N__33871));
    InMux I__7008 (
            .O(N__33881),
            .I(N__33866));
    InMux I__7007 (
            .O(N__33880),
            .I(N__33866));
    InMux I__7006 (
            .O(N__33877),
            .I(N__33863));
    CascadeMux I__7005 (
            .O(N__33876),
            .I(N__33860));
    CascadeMux I__7004 (
            .O(N__33875),
            .I(N__33855));
    CascadeMux I__7003 (
            .O(N__33874),
            .I(N__33852));
    LocalMux I__7002 (
            .O(N__33871),
            .I(N__33849));
    LocalMux I__7001 (
            .O(N__33866),
            .I(N__33844));
    LocalMux I__7000 (
            .O(N__33863),
            .I(N__33844));
    InMux I__6999 (
            .O(N__33860),
            .I(N__33841));
    CascadeMux I__6998 (
            .O(N__33859),
            .I(N__33838));
    InMux I__6997 (
            .O(N__33858),
            .I(N__33835));
    InMux I__6996 (
            .O(N__33855),
            .I(N__33829));
    InMux I__6995 (
            .O(N__33852),
            .I(N__33829));
    Span4Mux_v I__6994 (
            .O(N__33849),
            .I(N__33822));
    Span4Mux_s2_v I__6993 (
            .O(N__33844),
            .I(N__33822));
    LocalMux I__6992 (
            .O(N__33841),
            .I(N__33822));
    InMux I__6991 (
            .O(N__33838),
            .I(N__33819));
    LocalMux I__6990 (
            .O(N__33835),
            .I(N__33816));
    InMux I__6989 (
            .O(N__33834),
            .I(N__33813));
    LocalMux I__6988 (
            .O(N__33829),
            .I(N__33810));
    Span4Mux_h I__6987 (
            .O(N__33822),
            .I(N__33807));
    LocalMux I__6986 (
            .O(N__33819),
            .I(N__33798));
    Span12Mux_s5_v I__6985 (
            .O(N__33816),
            .I(N__33798));
    LocalMux I__6984 (
            .O(N__33813),
            .I(N__33798));
    Span12Mux_s2_h I__6983 (
            .O(N__33810),
            .I(N__33798));
    Span4Mux_h I__6982 (
            .O(N__33807),
            .I(N__33795));
    Odrv12 I__6981 (
            .O(N__33798),
            .I(r_SM_Main_0_adj_2441));
    Odrv4 I__6980 (
            .O(N__33795),
            .I(r_SM_Main_0_adj_2441));
    InMux I__6979 (
            .O(N__33790),
            .I(N__33787));
    LocalMux I__6978 (
            .O(N__33787),
            .I(N__33784));
    Span4Mux_h I__6977 (
            .O(N__33784),
            .I(N__33781));
    Span4Mux_h I__6976 (
            .O(N__33781),
            .I(N__33777));
    InMux I__6975 (
            .O(N__33780),
            .I(N__33774));
    Span4Mux_h I__6974 (
            .O(N__33777),
            .I(N__33771));
    LocalMux I__6973 (
            .O(N__33774),
            .I(\c0.rx.r_SM_Main_2_N_2096_0 ));
    Odrv4 I__6972 (
            .O(N__33771),
            .I(\c0.rx.r_SM_Main_2_N_2096_0 ));
    CascadeMux I__6971 (
            .O(N__33766),
            .I(N__33760));
    CascadeMux I__6970 (
            .O(N__33765),
            .I(N__33755));
    InMux I__6969 (
            .O(N__33764),
            .I(N__33748));
    InMux I__6968 (
            .O(N__33763),
            .I(N__33748));
    InMux I__6967 (
            .O(N__33760),
            .I(N__33741));
    InMux I__6966 (
            .O(N__33759),
            .I(N__33741));
    InMux I__6965 (
            .O(N__33758),
            .I(N__33738));
    InMux I__6964 (
            .O(N__33755),
            .I(N__33735));
    InMux I__6963 (
            .O(N__33754),
            .I(N__33732));
    InMux I__6962 (
            .O(N__33753),
            .I(N__33728));
    LocalMux I__6961 (
            .O(N__33748),
            .I(N__33725));
    InMux I__6960 (
            .O(N__33747),
            .I(N__33722));
    InMux I__6959 (
            .O(N__33746),
            .I(N__33719));
    LocalMux I__6958 (
            .O(N__33741),
            .I(N__33716));
    LocalMux I__6957 (
            .O(N__33738),
            .I(N__33713));
    LocalMux I__6956 (
            .O(N__33735),
            .I(N__33710));
    LocalMux I__6955 (
            .O(N__33732),
            .I(N__33707));
    InMux I__6954 (
            .O(N__33731),
            .I(N__33704));
    LocalMux I__6953 (
            .O(N__33728),
            .I(N__33699));
    Span4Mux_v I__6952 (
            .O(N__33725),
            .I(N__33699));
    LocalMux I__6951 (
            .O(N__33722),
            .I(N__33696));
    LocalMux I__6950 (
            .O(N__33719),
            .I(N__33689));
    Span4Mux_h I__6949 (
            .O(N__33716),
            .I(N__33689));
    Span4Mux_v I__6948 (
            .O(N__33713),
            .I(N__33689));
    Span4Mux_v I__6947 (
            .O(N__33710),
            .I(N__33684));
    Span4Mux_s2_v I__6946 (
            .O(N__33707),
            .I(N__33684));
    LocalMux I__6945 (
            .O(N__33704),
            .I(N__33681));
    Span4Mux_v I__6944 (
            .O(N__33699),
            .I(N__33676));
    Span4Mux_s2_v I__6943 (
            .O(N__33696),
            .I(N__33676));
    Span4Mux_v I__6942 (
            .O(N__33689),
            .I(N__33671));
    Span4Mux_h I__6941 (
            .O(N__33684),
            .I(N__33671));
    Span4Mux_v I__6940 (
            .O(N__33681),
            .I(N__33666));
    Span4Mux_h I__6939 (
            .O(N__33676),
            .I(N__33666));
    Odrv4 I__6938 (
            .O(N__33671),
            .I(r_Rx_Data));
    Odrv4 I__6937 (
            .O(N__33666),
            .I(r_Rx_Data));
    InMux I__6936 (
            .O(N__33661),
            .I(N__33658));
    LocalMux I__6935 (
            .O(N__33658),
            .I(n1));
    InMux I__6934 (
            .O(N__33655),
            .I(N__33652));
    LocalMux I__6933 (
            .O(N__33652),
            .I(N__33649));
    Span4Mux_v I__6932 (
            .O(N__33649),
            .I(N__33646));
    Odrv4 I__6931 (
            .O(N__33646),
            .I(\c0.n17915 ));
    CascadeMux I__6930 (
            .O(N__33643),
            .I(N__33640));
    InMux I__6929 (
            .O(N__33640),
            .I(N__33634));
    InMux I__6928 (
            .O(N__33639),
            .I(N__33634));
    LocalMux I__6927 (
            .O(N__33634),
            .I(data_out_frame2_18_1));
    CascadeMux I__6926 (
            .O(N__33631),
            .I(\c0.n17909_cascade_ ));
    InMux I__6925 (
            .O(N__33628),
            .I(N__33625));
    LocalMux I__6924 (
            .O(N__33625),
            .I(N__33622));
    Odrv4 I__6923 (
            .O(N__33622),
            .I(\c0.n6 ));
    InMux I__6922 (
            .O(N__33619),
            .I(N__33616));
    LocalMux I__6921 (
            .O(N__33616),
            .I(\c0.n18107 ));
    CascadeMux I__6920 (
            .O(N__33613),
            .I(N__33610));
    InMux I__6919 (
            .O(N__33610),
            .I(N__33607));
    LocalMux I__6918 (
            .O(N__33607),
            .I(N__33604));
    Odrv12 I__6917 (
            .O(N__33604),
            .I(\c0.n17579 ));
    InMux I__6916 (
            .O(N__33601),
            .I(N__33598));
    LocalMux I__6915 (
            .O(N__33598),
            .I(\c0.n17912 ));
    InMux I__6914 (
            .O(N__33595),
            .I(N__33592));
    LocalMux I__6913 (
            .O(N__33592),
            .I(\c0.n18110 ));
    CascadeMux I__6912 (
            .O(N__33589),
            .I(\c0.n22_adj_2359_cascade_ ));
    InMux I__6911 (
            .O(N__33586),
            .I(N__33583));
    LocalMux I__6910 (
            .O(N__33583),
            .I(\c0.n9758 ));
    SRMux I__6909 (
            .O(N__33580),
            .I(N__33577));
    LocalMux I__6908 (
            .O(N__33577),
            .I(N__33574));
    Span4Mux_h I__6907 (
            .O(N__33574),
            .I(N__33571));
    Odrv4 I__6906 (
            .O(N__33571),
            .I(\c0.n13496 ));
    CascadeMux I__6905 (
            .O(N__33568),
            .I(N__33565));
    InMux I__6904 (
            .O(N__33565),
            .I(N__33561));
    CascadeMux I__6903 (
            .O(N__33564),
            .I(N__33558));
    LocalMux I__6902 (
            .O(N__33561),
            .I(N__33553));
    InMux I__6901 (
            .O(N__33558),
            .I(N__33548));
    InMux I__6900 (
            .O(N__33557),
            .I(N__33548));
    InMux I__6899 (
            .O(N__33556),
            .I(N__33545));
    Span4Mux_v I__6898 (
            .O(N__33553),
            .I(N__33538));
    LocalMux I__6897 (
            .O(N__33548),
            .I(N__33538));
    LocalMux I__6896 (
            .O(N__33545),
            .I(N__33538));
    Odrv4 I__6895 (
            .O(N__33538),
            .I(data_out_frame2_7_3));
    InMux I__6894 (
            .O(N__33535),
            .I(N__33527));
    InMux I__6893 (
            .O(N__33534),
            .I(N__33524));
    InMux I__6892 (
            .O(N__33533),
            .I(N__33518));
    InMux I__6891 (
            .O(N__33532),
            .I(N__33512));
    InMux I__6890 (
            .O(N__33531),
            .I(N__33509));
    InMux I__6889 (
            .O(N__33530),
            .I(N__33506));
    LocalMux I__6888 (
            .O(N__33527),
            .I(N__33501));
    LocalMux I__6887 (
            .O(N__33524),
            .I(N__33501));
    InMux I__6886 (
            .O(N__33523),
            .I(N__33494));
    InMux I__6885 (
            .O(N__33522),
            .I(N__33494));
    InMux I__6884 (
            .O(N__33521),
            .I(N__33494));
    LocalMux I__6883 (
            .O(N__33518),
            .I(N__33490));
    InMux I__6882 (
            .O(N__33517),
            .I(N__33487));
    InMux I__6881 (
            .O(N__33516),
            .I(N__33482));
    InMux I__6880 (
            .O(N__33515),
            .I(N__33482));
    LocalMux I__6879 (
            .O(N__33512),
            .I(N__33479));
    LocalMux I__6878 (
            .O(N__33509),
            .I(N__33467));
    LocalMux I__6877 (
            .O(N__33506),
            .I(N__33467));
    Span4Mux_h I__6876 (
            .O(N__33501),
            .I(N__33467));
    LocalMux I__6875 (
            .O(N__33494),
            .I(N__33467));
    InMux I__6874 (
            .O(N__33493),
            .I(N__33464));
    Sp12to4 I__6873 (
            .O(N__33490),
            .I(N__33455));
    LocalMux I__6872 (
            .O(N__33487),
            .I(N__33455));
    LocalMux I__6871 (
            .O(N__33482),
            .I(N__33455));
    Span12Mux_v I__6870 (
            .O(N__33479),
            .I(N__33455));
    InMux I__6869 (
            .O(N__33478),
            .I(N__33450));
    InMux I__6868 (
            .O(N__33477),
            .I(N__33450));
    InMux I__6867 (
            .O(N__33476),
            .I(N__33447));
    Span4Mux_v I__6866 (
            .O(N__33467),
            .I(N__33444));
    LocalMux I__6865 (
            .O(N__33464),
            .I(FRAME_MATCHER_state_2));
    Odrv12 I__6864 (
            .O(N__33455),
            .I(FRAME_MATCHER_state_2));
    LocalMux I__6863 (
            .O(N__33450),
            .I(FRAME_MATCHER_state_2));
    LocalMux I__6862 (
            .O(N__33447),
            .I(FRAME_MATCHER_state_2));
    Odrv4 I__6861 (
            .O(N__33444),
            .I(FRAME_MATCHER_state_2));
    CascadeMux I__6860 (
            .O(N__33433),
            .I(N__33430));
    InMux I__6859 (
            .O(N__33430),
            .I(N__33426));
    InMux I__6858 (
            .O(N__33429),
            .I(N__33422));
    LocalMux I__6857 (
            .O(N__33426),
            .I(N__33419));
    InMux I__6856 (
            .O(N__33425),
            .I(N__33416));
    LocalMux I__6855 (
            .O(N__33422),
            .I(N__33413));
    Span4Mux_v I__6854 (
            .O(N__33419),
            .I(N__33409));
    LocalMux I__6853 (
            .O(N__33416),
            .I(N__33406));
    Span4Mux_h I__6852 (
            .O(N__33413),
            .I(N__33403));
    InMux I__6851 (
            .O(N__33412),
            .I(N__33398));
    Span4Mux_v I__6850 (
            .O(N__33409),
            .I(N__33392));
    Span4Mux_v I__6849 (
            .O(N__33406),
            .I(N__33392));
    Sp12to4 I__6848 (
            .O(N__33403),
            .I(N__33389));
    InMux I__6847 (
            .O(N__33402),
            .I(N__33386));
    InMux I__6846 (
            .O(N__33401),
            .I(N__33383));
    LocalMux I__6845 (
            .O(N__33398),
            .I(N__33380));
    InMux I__6844 (
            .O(N__33397),
            .I(N__33377));
    Sp12to4 I__6843 (
            .O(N__33392),
            .I(N__33372));
    Span12Mux_v I__6842 (
            .O(N__33389),
            .I(N__33372));
    LocalMux I__6841 (
            .O(N__33386),
            .I(N__33365));
    LocalMux I__6840 (
            .O(N__33383),
            .I(N__33365));
    Span4Mux_v I__6839 (
            .O(N__33380),
            .I(N__33365));
    LocalMux I__6838 (
            .O(N__33377),
            .I(\c0.FRAME_MATCHER_state_3 ));
    Odrv12 I__6837 (
            .O(N__33372),
            .I(\c0.FRAME_MATCHER_state_3 ));
    Odrv4 I__6836 (
            .O(N__33365),
            .I(\c0.FRAME_MATCHER_state_3 ));
    InMux I__6835 (
            .O(N__33358),
            .I(N__33353));
    InMux I__6834 (
            .O(N__33357),
            .I(N__33349));
    InMux I__6833 (
            .O(N__33356),
            .I(N__33346));
    LocalMux I__6832 (
            .O(N__33353),
            .I(N__33343));
    InMux I__6831 (
            .O(N__33352),
            .I(N__33340));
    LocalMux I__6830 (
            .O(N__33349),
            .I(N__33335));
    LocalMux I__6829 (
            .O(N__33346),
            .I(N__33335));
    Span4Mux_h I__6828 (
            .O(N__33343),
            .I(N__33328));
    LocalMux I__6827 (
            .O(N__33340),
            .I(N__33328));
    Span4Mux_v I__6826 (
            .O(N__33335),
            .I(N__33328));
    Span4Mux_h I__6825 (
            .O(N__33328),
            .I(N__33325));
    Odrv4 I__6824 (
            .O(N__33325),
            .I(\c0.n62 ));
    InMux I__6823 (
            .O(N__33322),
            .I(N__33316));
    InMux I__6822 (
            .O(N__33321),
            .I(N__33313));
    InMux I__6821 (
            .O(N__33320),
            .I(N__33310));
    InMux I__6820 (
            .O(N__33319),
            .I(N__33307));
    LocalMux I__6819 (
            .O(N__33316),
            .I(N__33304));
    LocalMux I__6818 (
            .O(N__33313),
            .I(\c0.n13464 ));
    LocalMux I__6817 (
            .O(N__33310),
            .I(\c0.n13464 ));
    LocalMux I__6816 (
            .O(N__33307),
            .I(\c0.n13464 ));
    Odrv12 I__6815 (
            .O(N__33304),
            .I(\c0.n13464 ));
    CascadeMux I__6814 (
            .O(N__33295),
            .I(\c0.n2_adj_2330_cascade_ ));
    SRMux I__6813 (
            .O(N__33292),
            .I(N__33289));
    LocalMux I__6812 (
            .O(N__33289),
            .I(N__33286));
    Span4Mux_h I__6811 (
            .O(N__33286),
            .I(N__33283));
    Odrv4 I__6810 (
            .O(N__33283),
            .I(\c0.n16377 ));
    InMux I__6809 (
            .O(N__33280),
            .I(N__33273));
    InMux I__6808 (
            .O(N__33279),
            .I(N__33270));
    InMux I__6807 (
            .O(N__33278),
            .I(N__33262));
    InMux I__6806 (
            .O(N__33277),
            .I(N__33251));
    InMux I__6805 (
            .O(N__33276),
            .I(N__33248));
    LocalMux I__6804 (
            .O(N__33273),
            .I(N__33242));
    LocalMux I__6803 (
            .O(N__33270),
            .I(N__33242));
    InMux I__6802 (
            .O(N__33269),
            .I(N__33239));
    InMux I__6801 (
            .O(N__33268),
            .I(N__33236));
    InMux I__6800 (
            .O(N__33267),
            .I(N__33233));
    InMux I__6799 (
            .O(N__33266),
            .I(N__33230));
    InMux I__6798 (
            .O(N__33265),
            .I(N__33227));
    LocalMux I__6797 (
            .O(N__33262),
            .I(N__33222));
    InMux I__6796 (
            .O(N__33261),
            .I(N__33219));
    InMux I__6795 (
            .O(N__33260),
            .I(N__33216));
    InMux I__6794 (
            .O(N__33259),
            .I(N__33213));
    InMux I__6793 (
            .O(N__33258),
            .I(N__33210));
    InMux I__6792 (
            .O(N__33257),
            .I(N__33205));
    InMux I__6791 (
            .O(N__33256),
            .I(N__33202));
    InMux I__6790 (
            .O(N__33255),
            .I(N__33199));
    InMux I__6789 (
            .O(N__33254),
            .I(N__33196));
    LocalMux I__6788 (
            .O(N__33251),
            .I(N__33190));
    LocalMux I__6787 (
            .O(N__33248),
            .I(N__33190));
    InMux I__6786 (
            .O(N__33247),
            .I(N__33187));
    Span4Mux_v I__6785 (
            .O(N__33242),
            .I(N__33168));
    LocalMux I__6784 (
            .O(N__33239),
            .I(N__33168));
    LocalMux I__6783 (
            .O(N__33236),
            .I(N__33168));
    LocalMux I__6782 (
            .O(N__33233),
            .I(N__33168));
    LocalMux I__6781 (
            .O(N__33230),
            .I(N__33168));
    LocalMux I__6780 (
            .O(N__33227),
            .I(N__33168));
    InMux I__6779 (
            .O(N__33226),
            .I(N__33165));
    InMux I__6778 (
            .O(N__33225),
            .I(N__33162));
    Span4Mux_v I__6777 (
            .O(N__33222),
            .I(N__33150));
    LocalMux I__6776 (
            .O(N__33219),
            .I(N__33150));
    LocalMux I__6775 (
            .O(N__33216),
            .I(N__33150));
    LocalMux I__6774 (
            .O(N__33213),
            .I(N__33150));
    LocalMux I__6773 (
            .O(N__33210),
            .I(N__33150));
    InMux I__6772 (
            .O(N__33209),
            .I(N__33147));
    InMux I__6771 (
            .O(N__33208),
            .I(N__33144));
    LocalMux I__6770 (
            .O(N__33205),
            .I(N__33135));
    LocalMux I__6769 (
            .O(N__33202),
            .I(N__33135));
    LocalMux I__6768 (
            .O(N__33199),
            .I(N__33135));
    LocalMux I__6767 (
            .O(N__33196),
            .I(N__33135));
    InMux I__6766 (
            .O(N__33195),
            .I(N__33132));
    Span4Mux_v I__6765 (
            .O(N__33190),
            .I(N__33127));
    LocalMux I__6764 (
            .O(N__33187),
            .I(N__33127));
    InMux I__6763 (
            .O(N__33186),
            .I(N__33124));
    InMux I__6762 (
            .O(N__33185),
            .I(N__33121));
    InMux I__6761 (
            .O(N__33184),
            .I(N__33118));
    InMux I__6760 (
            .O(N__33183),
            .I(N__33115));
    InMux I__6759 (
            .O(N__33182),
            .I(N__33112));
    InMux I__6758 (
            .O(N__33181),
            .I(N__33109));
    Span4Mux_v I__6757 (
            .O(N__33168),
            .I(N__33102));
    LocalMux I__6756 (
            .O(N__33165),
            .I(N__33102));
    LocalMux I__6755 (
            .O(N__33162),
            .I(N__33102));
    InMux I__6754 (
            .O(N__33161),
            .I(N__33099));
    Span4Mux_v I__6753 (
            .O(N__33150),
            .I(N__33094));
    LocalMux I__6752 (
            .O(N__33147),
            .I(N__33091));
    LocalMux I__6751 (
            .O(N__33144),
            .I(N__33088));
    Span4Mux_h I__6750 (
            .O(N__33135),
            .I(N__33079));
    LocalMux I__6749 (
            .O(N__33132),
            .I(N__33079));
    Span4Mux_h I__6748 (
            .O(N__33127),
            .I(N__33079));
    LocalMux I__6747 (
            .O(N__33124),
            .I(N__33079));
    LocalMux I__6746 (
            .O(N__33121),
            .I(N__33076));
    LocalMux I__6745 (
            .O(N__33118),
            .I(N__33073));
    LocalMux I__6744 (
            .O(N__33115),
            .I(N__33068));
    LocalMux I__6743 (
            .O(N__33112),
            .I(N__33068));
    LocalMux I__6742 (
            .O(N__33109),
            .I(N__33065));
    Span4Mux_v I__6741 (
            .O(N__33102),
            .I(N__33060));
    LocalMux I__6740 (
            .O(N__33099),
            .I(N__33060));
    InMux I__6739 (
            .O(N__33098),
            .I(N__33057));
    CascadeMux I__6738 (
            .O(N__33097),
            .I(N__33054));
    Span4Mux_h I__6737 (
            .O(N__33094),
            .I(N__33048));
    Span4Mux_v I__6736 (
            .O(N__33091),
            .I(N__33048));
    Span12Mux_h I__6735 (
            .O(N__33088),
            .I(N__33045));
    Span4Mux_v I__6734 (
            .O(N__33079),
            .I(N__33040));
    Span4Mux_v I__6733 (
            .O(N__33076),
            .I(N__33040));
    Span4Mux_h I__6732 (
            .O(N__33073),
            .I(N__33037));
    Span4Mux_v I__6731 (
            .O(N__33068),
            .I(N__33030));
    Span4Mux_h I__6730 (
            .O(N__33065),
            .I(N__33030));
    Span4Mux_h I__6729 (
            .O(N__33060),
            .I(N__33030));
    LocalMux I__6728 (
            .O(N__33057),
            .I(N__33027));
    InMux I__6727 (
            .O(N__33054),
            .I(N__33022));
    InMux I__6726 (
            .O(N__33053),
            .I(N__33022));
    Odrv4 I__6725 (
            .O(N__33048),
            .I(n9452));
    Odrv12 I__6724 (
            .O(N__33045),
            .I(n9452));
    Odrv4 I__6723 (
            .O(N__33040),
            .I(n9452));
    Odrv4 I__6722 (
            .O(N__33037),
            .I(n9452));
    Odrv4 I__6721 (
            .O(N__33030),
            .I(n9452));
    Odrv12 I__6720 (
            .O(N__33027),
            .I(n9452));
    LocalMux I__6719 (
            .O(N__33022),
            .I(n9452));
    InMux I__6718 (
            .O(N__33007),
            .I(N__32993));
    InMux I__6717 (
            .O(N__33006),
            .I(N__32990));
    InMux I__6716 (
            .O(N__33005),
            .I(N__32985));
    InMux I__6715 (
            .O(N__33004),
            .I(N__32982));
    InMux I__6714 (
            .O(N__33003),
            .I(N__32979));
    InMux I__6713 (
            .O(N__33002),
            .I(N__32976));
    InMux I__6712 (
            .O(N__33001),
            .I(N__32973));
    InMux I__6711 (
            .O(N__33000),
            .I(N__32970));
    InMux I__6710 (
            .O(N__32999),
            .I(N__32967));
    InMux I__6709 (
            .O(N__32998),
            .I(N__32964));
    InMux I__6708 (
            .O(N__32997),
            .I(N__32961));
    InMux I__6707 (
            .O(N__32996),
            .I(N__32956));
    LocalMux I__6706 (
            .O(N__32993),
            .I(N__32951));
    LocalMux I__6705 (
            .O(N__32990),
            .I(N__32951));
    InMux I__6704 (
            .O(N__32989),
            .I(N__32948));
    InMux I__6703 (
            .O(N__32988),
            .I(N__32943));
    LocalMux I__6702 (
            .O(N__32985),
            .I(N__32938));
    LocalMux I__6701 (
            .O(N__32982),
            .I(N__32938));
    LocalMux I__6700 (
            .O(N__32979),
            .I(N__32935));
    LocalMux I__6699 (
            .O(N__32976),
            .I(N__32922));
    LocalMux I__6698 (
            .O(N__32973),
            .I(N__32922));
    LocalMux I__6697 (
            .O(N__32970),
            .I(N__32922));
    LocalMux I__6696 (
            .O(N__32967),
            .I(N__32922));
    LocalMux I__6695 (
            .O(N__32964),
            .I(N__32922));
    LocalMux I__6694 (
            .O(N__32961),
            .I(N__32922));
    InMux I__6693 (
            .O(N__32960),
            .I(N__32919));
    InMux I__6692 (
            .O(N__32959),
            .I(N__32915));
    LocalMux I__6691 (
            .O(N__32956),
            .I(N__32903));
    Span4Mux_v I__6690 (
            .O(N__32951),
            .I(N__32903));
    LocalMux I__6689 (
            .O(N__32948),
            .I(N__32903));
    InMux I__6688 (
            .O(N__32947),
            .I(N__32900));
    InMux I__6687 (
            .O(N__32946),
            .I(N__32897));
    LocalMux I__6686 (
            .O(N__32943),
            .I(N__32889));
    Span4Mux_v I__6685 (
            .O(N__32938),
            .I(N__32880));
    Span4Mux_s1_h I__6684 (
            .O(N__32935),
            .I(N__32880));
    Span4Mux_v I__6683 (
            .O(N__32922),
            .I(N__32880));
    LocalMux I__6682 (
            .O(N__32919),
            .I(N__32880));
    InMux I__6681 (
            .O(N__32918),
            .I(N__32877));
    LocalMux I__6680 (
            .O(N__32915),
            .I(N__32874));
    InMux I__6679 (
            .O(N__32914),
            .I(N__32871));
    InMux I__6678 (
            .O(N__32913),
            .I(N__32868));
    InMux I__6677 (
            .O(N__32912),
            .I(N__32865));
    InMux I__6676 (
            .O(N__32911),
            .I(N__32862));
    InMux I__6675 (
            .O(N__32910),
            .I(N__32859));
    Span4Mux_h I__6674 (
            .O(N__32903),
            .I(N__32852));
    LocalMux I__6673 (
            .O(N__32900),
            .I(N__32852));
    LocalMux I__6672 (
            .O(N__32897),
            .I(N__32852));
    InMux I__6671 (
            .O(N__32896),
            .I(N__32849));
    InMux I__6670 (
            .O(N__32895),
            .I(N__32842));
    InMux I__6669 (
            .O(N__32894),
            .I(N__32842));
    InMux I__6668 (
            .O(N__32893),
            .I(N__32839));
    InMux I__6667 (
            .O(N__32892),
            .I(N__32836));
    Span4Mux_v I__6666 (
            .O(N__32889),
            .I(N__32827));
    Span4Mux_h I__6665 (
            .O(N__32880),
            .I(N__32827));
    LocalMux I__6664 (
            .O(N__32877),
            .I(N__32827));
    Span4Mux_v I__6663 (
            .O(N__32874),
            .I(N__32823));
    LocalMux I__6662 (
            .O(N__32871),
            .I(N__32816));
    LocalMux I__6661 (
            .O(N__32868),
            .I(N__32816));
    LocalMux I__6660 (
            .O(N__32865),
            .I(N__32816));
    LocalMux I__6659 (
            .O(N__32862),
            .I(N__32807));
    LocalMux I__6658 (
            .O(N__32859),
            .I(N__32807));
    Span4Mux_v I__6657 (
            .O(N__32852),
            .I(N__32807));
    LocalMux I__6656 (
            .O(N__32849),
            .I(N__32807));
    InMux I__6655 (
            .O(N__32848),
            .I(N__32804));
    InMux I__6654 (
            .O(N__32847),
            .I(N__32799));
    LocalMux I__6653 (
            .O(N__32842),
            .I(N__32796));
    LocalMux I__6652 (
            .O(N__32839),
            .I(N__32791));
    LocalMux I__6651 (
            .O(N__32836),
            .I(N__32791));
    InMux I__6650 (
            .O(N__32835),
            .I(N__32787));
    InMux I__6649 (
            .O(N__32834),
            .I(N__32784));
    Span4Mux_h I__6648 (
            .O(N__32827),
            .I(N__32780));
    InMux I__6647 (
            .O(N__32826),
            .I(N__32777));
    Span4Mux_h I__6646 (
            .O(N__32823),
            .I(N__32768));
    Span4Mux_v I__6645 (
            .O(N__32816),
            .I(N__32768));
    Span4Mux_s3_h I__6644 (
            .O(N__32807),
            .I(N__32768));
    LocalMux I__6643 (
            .O(N__32804),
            .I(N__32768));
    InMux I__6642 (
            .O(N__32803),
            .I(N__32765));
    InMux I__6641 (
            .O(N__32802),
            .I(N__32762));
    LocalMux I__6640 (
            .O(N__32799),
            .I(N__32755));
    Span4Mux_v I__6639 (
            .O(N__32796),
            .I(N__32755));
    Span4Mux_h I__6638 (
            .O(N__32791),
            .I(N__32755));
    InMux I__6637 (
            .O(N__32790),
            .I(N__32752));
    LocalMux I__6636 (
            .O(N__32787),
            .I(N__32747));
    LocalMux I__6635 (
            .O(N__32784),
            .I(N__32747));
    InMux I__6634 (
            .O(N__32783),
            .I(N__32744));
    Odrv4 I__6633 (
            .O(N__32780),
            .I(n12933));
    LocalMux I__6632 (
            .O(N__32777),
            .I(n12933));
    Odrv4 I__6631 (
            .O(N__32768),
            .I(n12933));
    LocalMux I__6630 (
            .O(N__32765),
            .I(n12933));
    LocalMux I__6629 (
            .O(N__32762),
            .I(n12933));
    Odrv4 I__6628 (
            .O(N__32755),
            .I(n12933));
    LocalMux I__6627 (
            .O(N__32752),
            .I(n12933));
    Odrv12 I__6626 (
            .O(N__32747),
            .I(n12933));
    LocalMux I__6625 (
            .O(N__32744),
            .I(n12933));
    InMux I__6624 (
            .O(N__32725),
            .I(N__32722));
    LocalMux I__6623 (
            .O(N__32722),
            .I(N__32719));
    Span4Mux_h I__6622 (
            .O(N__32719),
            .I(N__32716));
    Span4Mux_h I__6621 (
            .O(N__32716),
            .I(N__32713));
    Odrv4 I__6620 (
            .O(N__32713),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_0 ));
    InMux I__6619 (
            .O(N__32710),
            .I(N__32706));
    CascadeMux I__6618 (
            .O(N__32709),
            .I(N__32701));
    LocalMux I__6617 (
            .O(N__32706),
            .I(N__32698));
    InMux I__6616 (
            .O(N__32705),
            .I(N__32695));
    InMux I__6615 (
            .O(N__32704),
            .I(N__32692));
    InMux I__6614 (
            .O(N__32701),
            .I(N__32687));
    Span4Mux_v I__6613 (
            .O(N__32698),
            .I(N__32682));
    LocalMux I__6612 (
            .O(N__32695),
            .I(N__32682));
    LocalMux I__6611 (
            .O(N__32692),
            .I(N__32679));
    InMux I__6610 (
            .O(N__32691),
            .I(N__32676));
    InMux I__6609 (
            .O(N__32690),
            .I(N__32673));
    LocalMux I__6608 (
            .O(N__32687),
            .I(N__32670));
    Span4Mux_v I__6607 (
            .O(N__32682),
            .I(N__32666));
    Span4Mux_v I__6606 (
            .O(N__32679),
            .I(N__32659));
    LocalMux I__6605 (
            .O(N__32676),
            .I(N__32659));
    LocalMux I__6604 (
            .O(N__32673),
            .I(N__32659));
    Span4Mux_v I__6603 (
            .O(N__32670),
            .I(N__32656));
    InMux I__6602 (
            .O(N__32669),
            .I(N__32653));
    Sp12to4 I__6601 (
            .O(N__32666),
            .I(N__32650));
    Span4Mux_v I__6600 (
            .O(N__32659),
            .I(N__32645));
    Span4Mux_h I__6599 (
            .O(N__32656),
            .I(N__32645));
    LocalMux I__6598 (
            .O(N__32653),
            .I(N__32642));
    Span12Mux_s10_h I__6597 (
            .O(N__32650),
            .I(N__32639));
    Span4Mux_h I__6596 (
            .O(N__32645),
            .I(N__32636));
    Span4Mux_h I__6595 (
            .O(N__32642),
            .I(N__32633));
    Odrv12 I__6594 (
            .O(N__32639),
            .I(\c0.FRAME_MATCHER_i_0 ));
    Odrv4 I__6593 (
            .O(N__32636),
            .I(\c0.FRAME_MATCHER_i_0 ));
    Odrv4 I__6592 (
            .O(N__32633),
            .I(\c0.FRAME_MATCHER_i_0 ));
    SRMux I__6591 (
            .O(N__32626),
            .I(N__32623));
    LocalMux I__6590 (
            .O(N__32623),
            .I(N__32620));
    Span4Mux_v I__6589 (
            .O(N__32620),
            .I(N__32617));
    Odrv4 I__6588 (
            .O(N__32617),
            .I(\c0.n3 ));
    InMux I__6587 (
            .O(N__32614),
            .I(N__32611));
    LocalMux I__6586 (
            .O(N__32611),
            .I(N__32606));
    InMux I__6585 (
            .O(N__32610),
            .I(N__32603));
    InMux I__6584 (
            .O(N__32609),
            .I(N__32600));
    Span4Mux_h I__6583 (
            .O(N__32606),
            .I(N__32597));
    LocalMux I__6582 (
            .O(N__32603),
            .I(\c0.FRAME_MATCHER_state_12 ));
    LocalMux I__6581 (
            .O(N__32600),
            .I(\c0.FRAME_MATCHER_state_12 ));
    Odrv4 I__6580 (
            .O(N__32597),
            .I(\c0.FRAME_MATCHER_state_12 ));
    InMux I__6579 (
            .O(N__32590),
            .I(N__32585));
    InMux I__6578 (
            .O(N__32589),
            .I(N__32578));
    InMux I__6577 (
            .O(N__32588),
            .I(N__32578));
    LocalMux I__6576 (
            .O(N__32585),
            .I(N__32575));
    CascadeMux I__6575 (
            .O(N__32584),
            .I(N__32572));
    CascadeMux I__6574 (
            .O(N__32583),
            .I(N__32568));
    LocalMux I__6573 (
            .O(N__32578),
            .I(N__32563));
    Span4Mux_h I__6572 (
            .O(N__32575),
            .I(N__32560));
    InMux I__6571 (
            .O(N__32572),
            .I(N__32549));
    InMux I__6570 (
            .O(N__32571),
            .I(N__32549));
    InMux I__6569 (
            .O(N__32568),
            .I(N__32549));
    InMux I__6568 (
            .O(N__32567),
            .I(N__32549));
    InMux I__6567 (
            .O(N__32566),
            .I(N__32549));
    Odrv12 I__6566 (
            .O(N__32563),
            .I(\c0.n4_adj_2360 ));
    Odrv4 I__6565 (
            .O(N__32560),
            .I(\c0.n4_adj_2360 ));
    LocalMux I__6564 (
            .O(N__32549),
            .I(\c0.n4_adj_2360 ));
    SRMux I__6563 (
            .O(N__32542),
            .I(N__32539));
    LocalMux I__6562 (
            .O(N__32539),
            .I(N__32536));
    Span4Mux_h I__6561 (
            .O(N__32536),
            .I(N__32533));
    Odrv4 I__6560 (
            .O(N__32533),
            .I(\c0.n16449 ));
    CascadeMux I__6559 (
            .O(N__32530),
            .I(N__32526));
    InMux I__6558 (
            .O(N__32529),
            .I(N__32523));
    InMux I__6557 (
            .O(N__32526),
            .I(N__32520));
    LocalMux I__6556 (
            .O(N__32523),
            .I(data_out_frame2_18_2));
    LocalMux I__6555 (
            .O(N__32520),
            .I(data_out_frame2_18_2));
    CascadeMux I__6554 (
            .O(N__32515),
            .I(\c0.n18119_cascade_ ));
    CascadeMux I__6553 (
            .O(N__32512),
            .I(\c0.n18122_cascade_ ));
    InMux I__6552 (
            .O(N__32509),
            .I(N__32506));
    LocalMux I__6551 (
            .O(N__32506),
            .I(N__32503));
    Span4Mux_v I__6550 (
            .O(N__32503),
            .I(N__32500));
    Span4Mux_v I__6549 (
            .O(N__32500),
            .I(N__32497));
    Odrv4 I__6548 (
            .O(N__32497),
            .I(\c0.tx2.r_Tx_Data_2 ));
    InMux I__6547 (
            .O(N__32494),
            .I(N__32491));
    LocalMux I__6546 (
            .O(N__32491),
            .I(N__32488));
    Odrv4 I__6545 (
            .O(N__32488),
            .I(\c0.n17340 ));
    InMux I__6544 (
            .O(N__32485),
            .I(N__32482));
    LocalMux I__6543 (
            .O(N__32482),
            .I(\c0.n2_adj_2137 ));
    InMux I__6542 (
            .O(N__32479),
            .I(N__32475));
    InMux I__6541 (
            .O(N__32478),
            .I(N__32472));
    LocalMux I__6540 (
            .O(N__32475),
            .I(\c0.data_out_1_4 ));
    LocalMux I__6539 (
            .O(N__32472),
            .I(\c0.data_out_1_4 ));
    InMux I__6538 (
            .O(N__32467),
            .I(N__32464));
    LocalMux I__6537 (
            .O(N__32464),
            .I(N__32461));
    Odrv12 I__6536 (
            .O(N__32461),
            .I(n16776));
    CascadeMux I__6535 (
            .O(N__32458),
            .I(N__32455));
    InMux I__6534 (
            .O(N__32455),
            .I(N__32451));
    InMux I__6533 (
            .O(N__32454),
            .I(N__32448));
    LocalMux I__6532 (
            .O(N__32451),
            .I(N__32444));
    LocalMux I__6531 (
            .O(N__32448),
            .I(N__32441));
    InMux I__6530 (
            .O(N__32447),
            .I(N__32438));
    Span4Mux_v I__6529 (
            .O(N__32444),
            .I(N__32435));
    Span4Mux_v I__6528 (
            .O(N__32441),
            .I(N__32432));
    LocalMux I__6527 (
            .O(N__32438),
            .I(N__32429));
    Span4Mux_h I__6526 (
            .O(N__32435),
            .I(N__32424));
    Span4Mux_s2_h I__6525 (
            .O(N__32432),
            .I(N__32424));
    Odrv4 I__6524 (
            .O(N__32429),
            .I(n17208));
    Odrv4 I__6523 (
            .O(N__32424),
            .I(n17208));
    InMux I__6522 (
            .O(N__32419),
            .I(N__32416));
    LocalMux I__6521 (
            .O(N__32416),
            .I(N__32413));
    Span4Mux_v I__6520 (
            .O(N__32413),
            .I(N__32410));
    Span4Mux_h I__6519 (
            .O(N__32410),
            .I(N__32407));
    Odrv4 I__6518 (
            .O(N__32407),
            .I(n8828));
    InMux I__6517 (
            .O(N__32404),
            .I(N__32398));
    InMux I__6516 (
            .O(N__32403),
            .I(N__32398));
    LocalMux I__6515 (
            .O(N__32398),
            .I(N__32393));
    InMux I__6514 (
            .O(N__32397),
            .I(N__32390));
    InMux I__6513 (
            .O(N__32396),
            .I(N__32386));
    Span4Mux_h I__6512 (
            .O(N__32393),
            .I(N__32383));
    LocalMux I__6511 (
            .O(N__32390),
            .I(N__32380));
    InMux I__6510 (
            .O(N__32389),
            .I(N__32377));
    LocalMux I__6509 (
            .O(N__32386),
            .I(\c0.FRAME_MATCHER_state_16 ));
    Odrv4 I__6508 (
            .O(N__32383),
            .I(\c0.FRAME_MATCHER_state_16 ));
    Odrv12 I__6507 (
            .O(N__32380),
            .I(\c0.FRAME_MATCHER_state_16 ));
    LocalMux I__6506 (
            .O(N__32377),
            .I(\c0.FRAME_MATCHER_state_16 ));
    InMux I__6505 (
            .O(N__32368),
            .I(N__32364));
    InMux I__6504 (
            .O(N__32367),
            .I(N__32361));
    LocalMux I__6503 (
            .O(N__32364),
            .I(N__32358));
    LocalMux I__6502 (
            .O(N__32361),
            .I(N__32355));
    Span4Mux_v I__6501 (
            .O(N__32358),
            .I(N__32352));
    Span4Mux_h I__6500 (
            .O(N__32355),
            .I(N__32349));
    Span4Mux_h I__6499 (
            .O(N__32352),
            .I(N__32344));
    Span4Mux_v I__6498 (
            .O(N__32349),
            .I(N__32344));
    Odrv4 I__6497 (
            .O(N__32344),
            .I(\c0.n47 ));
    CascadeMux I__6496 (
            .O(N__32341),
            .I(N__32338));
    InMux I__6495 (
            .O(N__32338),
            .I(N__32335));
    LocalMux I__6494 (
            .O(N__32335),
            .I(N__32332));
    Span12Mux_s10_h I__6493 (
            .O(N__32332),
            .I(N__32329));
    Odrv12 I__6492 (
            .O(N__32329),
            .I(\c0.n6_adj_2140 ));
    InMux I__6491 (
            .O(N__32326),
            .I(N__32319));
    InMux I__6490 (
            .O(N__32325),
            .I(N__32319));
    CascadeMux I__6489 (
            .O(N__32324),
            .I(N__32314));
    LocalMux I__6488 (
            .O(N__32319),
            .I(N__32311));
    InMux I__6487 (
            .O(N__32318),
            .I(N__32307));
    InMux I__6486 (
            .O(N__32317),
            .I(N__32303));
    InMux I__6485 (
            .O(N__32314),
            .I(N__32300));
    Span4Mux_v I__6484 (
            .O(N__32311),
            .I(N__32296));
    InMux I__6483 (
            .O(N__32310),
            .I(N__32293));
    LocalMux I__6482 (
            .O(N__32307),
            .I(N__32289));
    InMux I__6481 (
            .O(N__32306),
            .I(N__32286));
    LocalMux I__6480 (
            .O(N__32303),
            .I(N__32283));
    LocalMux I__6479 (
            .O(N__32300),
            .I(N__32280));
    InMux I__6478 (
            .O(N__32299),
            .I(N__32277));
    Span4Mux_h I__6477 (
            .O(N__32296),
            .I(N__32272));
    LocalMux I__6476 (
            .O(N__32293),
            .I(N__32272));
    InMux I__6475 (
            .O(N__32292),
            .I(N__32269));
    Span4Mux_v I__6474 (
            .O(N__32289),
            .I(N__32265));
    LocalMux I__6473 (
            .O(N__32286),
            .I(N__32262));
    Span4Mux_h I__6472 (
            .O(N__32283),
            .I(N__32253));
    Span4Mux_v I__6471 (
            .O(N__32280),
            .I(N__32253));
    LocalMux I__6470 (
            .O(N__32277),
            .I(N__32253));
    Span4Mux_v I__6469 (
            .O(N__32272),
            .I(N__32248));
    LocalMux I__6468 (
            .O(N__32269),
            .I(N__32248));
    InMux I__6467 (
            .O(N__32268),
            .I(N__32245));
    Span4Mux_h I__6466 (
            .O(N__32265),
            .I(N__32240));
    Span4Mux_v I__6465 (
            .O(N__32262),
            .I(N__32240));
    InMux I__6464 (
            .O(N__32261),
            .I(N__32235));
    InMux I__6463 (
            .O(N__32260),
            .I(N__32235));
    Span4Mux_h I__6462 (
            .O(N__32253),
            .I(N__32232));
    Span4Mux_h I__6461 (
            .O(N__32248),
            .I(N__32229));
    LocalMux I__6460 (
            .O(N__32245),
            .I(FRAME_MATCHER_state_1));
    Odrv4 I__6459 (
            .O(N__32240),
            .I(FRAME_MATCHER_state_1));
    LocalMux I__6458 (
            .O(N__32235),
            .I(FRAME_MATCHER_state_1));
    Odrv4 I__6457 (
            .O(N__32232),
            .I(FRAME_MATCHER_state_1));
    Odrv4 I__6456 (
            .O(N__32229),
            .I(FRAME_MATCHER_state_1));
    InMux I__6455 (
            .O(N__32218),
            .I(N__32215));
    LocalMux I__6454 (
            .O(N__32215),
            .I(N__32212));
    Span4Mux_v I__6453 (
            .O(N__32212),
            .I(N__32209));
    Odrv4 I__6452 (
            .O(N__32209),
            .I(\c0.n5_adj_2339 ));
    CascadeMux I__6451 (
            .O(N__32206),
            .I(\c0.n16814_cascade_ ));
    InMux I__6450 (
            .O(N__32203),
            .I(N__32200));
    LocalMux I__6449 (
            .O(N__32200),
            .I(N__32197));
    Odrv4 I__6448 (
            .O(N__32197),
            .I(\c0.tx2.n89 ));
    InMux I__6447 (
            .O(N__32194),
            .I(N__32187));
    InMux I__6446 (
            .O(N__32193),
            .I(N__32182));
    InMux I__6445 (
            .O(N__32192),
            .I(N__32182));
    InMux I__6444 (
            .O(N__32191),
            .I(N__32177));
    InMux I__6443 (
            .O(N__32190),
            .I(N__32177));
    LocalMux I__6442 (
            .O(N__32187),
            .I(\c0.FRAME_MATCHER_state_31 ));
    LocalMux I__6441 (
            .O(N__32182),
            .I(\c0.FRAME_MATCHER_state_31 ));
    LocalMux I__6440 (
            .O(N__32177),
            .I(\c0.FRAME_MATCHER_state_31 ));
    InMux I__6439 (
            .O(N__32170),
            .I(N__32166));
    InMux I__6438 (
            .O(N__32169),
            .I(N__32163));
    LocalMux I__6437 (
            .O(N__32166),
            .I(r_Tx_Data_7));
    LocalMux I__6436 (
            .O(N__32163),
            .I(r_Tx_Data_7));
    InMux I__6435 (
            .O(N__32158),
            .I(N__32155));
    LocalMux I__6434 (
            .O(N__32155),
            .I(\c0.n18014 ));
    CascadeMux I__6433 (
            .O(N__32152),
            .I(N__32149));
    InMux I__6432 (
            .O(N__32149),
            .I(N__32146));
    LocalMux I__6431 (
            .O(N__32146),
            .I(N__32143));
    Span4Mux_v I__6430 (
            .O(N__32143),
            .I(N__32140));
    Odrv4 I__6429 (
            .O(N__32140),
            .I(\c0.n17585 ));
    InMux I__6428 (
            .O(N__32137),
            .I(N__32134));
    LocalMux I__6427 (
            .O(N__32134),
            .I(n10_adj_2423));
    CascadeMux I__6426 (
            .O(N__32131),
            .I(n18044_cascade_));
    InMux I__6425 (
            .O(N__32128),
            .I(N__32125));
    LocalMux I__6424 (
            .O(N__32125),
            .I(n10_adj_2414));
    CascadeMux I__6423 (
            .O(N__32122),
            .I(N__32118));
    InMux I__6422 (
            .O(N__32121),
            .I(N__32115));
    InMux I__6421 (
            .O(N__32118),
            .I(N__32112));
    LocalMux I__6420 (
            .O(N__32115),
            .I(data_out_0_1));
    LocalMux I__6419 (
            .O(N__32112),
            .I(data_out_0_1));
    InMux I__6418 (
            .O(N__32107),
            .I(N__32104));
    LocalMux I__6417 (
            .O(N__32104),
            .I(N__32101));
    Odrv4 I__6416 (
            .O(N__32101),
            .I(\c0.n18080 ));
    InMux I__6415 (
            .O(N__32098),
            .I(N__32094));
    InMux I__6414 (
            .O(N__32097),
            .I(N__32091));
    LocalMux I__6413 (
            .O(N__32094),
            .I(data_out_3_7));
    LocalMux I__6412 (
            .O(N__32091),
            .I(data_out_3_7));
    CascadeMux I__6411 (
            .O(N__32086),
            .I(\c0.n29_cascade_ ));
    InMux I__6410 (
            .O(N__32083),
            .I(N__32079));
    InMux I__6409 (
            .O(N__32082),
            .I(N__32076));
    LocalMux I__6408 (
            .O(N__32079),
            .I(N__32073));
    LocalMux I__6407 (
            .O(N__32076),
            .I(r_Tx_Data_1));
    Odrv12 I__6406 (
            .O(N__32073),
            .I(r_Tx_Data_1));
    InMux I__6405 (
            .O(N__32068),
            .I(N__32062));
    InMux I__6404 (
            .O(N__32067),
            .I(N__32062));
    LocalMux I__6403 (
            .O(N__32062),
            .I(r_Tx_Data_5));
    InMux I__6402 (
            .O(N__32059),
            .I(N__32056));
    LocalMux I__6401 (
            .O(N__32056),
            .I(N__32052));
    InMux I__6400 (
            .O(N__32055),
            .I(N__32049));
    Span4Mux_h I__6399 (
            .O(N__32052),
            .I(N__32046));
    LocalMux I__6398 (
            .O(N__32049),
            .I(\c0.data_out_0_6 ));
    Odrv4 I__6397 (
            .O(N__32046),
            .I(\c0.data_out_0_6 ));
    CascadeMux I__6396 (
            .O(N__32041),
            .I(\c0.n9_adj_2143_cascade_ ));
    InMux I__6395 (
            .O(N__32038),
            .I(N__32035));
    LocalMux I__6394 (
            .O(N__32035),
            .I(\c0.n23 ));
    InMux I__6393 (
            .O(N__32032),
            .I(N__32029));
    LocalMux I__6392 (
            .O(N__32029),
            .I(N__32026));
    Span4Mux_h I__6391 (
            .O(N__32026),
            .I(N__32023));
    Odrv4 I__6390 (
            .O(N__32023),
            .I(\c0.n17547 ));
    CascadeMux I__6389 (
            .O(N__32020),
            .I(\c0.n5_adj_2326_cascade_ ));
    InMux I__6388 (
            .O(N__32017),
            .I(N__32014));
    LocalMux I__6387 (
            .O(N__32014),
            .I(N__32011));
    Odrv4 I__6386 (
            .O(N__32011),
            .I(\c0.n18023 ));
    InMux I__6385 (
            .O(N__32008),
            .I(N__32002));
    InMux I__6384 (
            .O(N__32007),
            .I(N__32002));
    LocalMux I__6383 (
            .O(N__32002),
            .I(N__31985));
    InMux I__6382 (
            .O(N__32001),
            .I(N__31976));
    InMux I__6381 (
            .O(N__32000),
            .I(N__31976));
    InMux I__6380 (
            .O(N__31999),
            .I(N__31976));
    InMux I__6379 (
            .O(N__31998),
            .I(N__31976));
    InMux I__6378 (
            .O(N__31997),
            .I(N__31967));
    InMux I__6377 (
            .O(N__31996),
            .I(N__31967));
    InMux I__6376 (
            .O(N__31995),
            .I(N__31967));
    InMux I__6375 (
            .O(N__31994),
            .I(N__31967));
    InMux I__6374 (
            .O(N__31993),
            .I(N__31964));
    InMux I__6373 (
            .O(N__31992),
            .I(N__31961));
    InMux I__6372 (
            .O(N__31991),
            .I(N__31956));
    InMux I__6371 (
            .O(N__31990),
            .I(N__31956));
    InMux I__6370 (
            .O(N__31989),
            .I(N__31951));
    InMux I__6369 (
            .O(N__31988),
            .I(N__31951));
    Odrv12 I__6368 (
            .O(N__31985),
            .I(\c0.n16891 ));
    LocalMux I__6367 (
            .O(N__31976),
            .I(\c0.n16891 ));
    LocalMux I__6366 (
            .O(N__31967),
            .I(\c0.n16891 ));
    LocalMux I__6365 (
            .O(N__31964),
            .I(\c0.n16891 ));
    LocalMux I__6364 (
            .O(N__31961),
            .I(\c0.n16891 ));
    LocalMux I__6363 (
            .O(N__31956),
            .I(\c0.n16891 ));
    LocalMux I__6362 (
            .O(N__31951),
            .I(\c0.n16891 ));
    InMux I__6361 (
            .O(N__31936),
            .I(N__31926));
    InMux I__6360 (
            .O(N__31935),
            .I(N__31926));
    InMux I__6359 (
            .O(N__31934),
            .I(N__31926));
    InMux I__6358 (
            .O(N__31933),
            .I(N__31914));
    LocalMux I__6357 (
            .O(N__31926),
            .I(N__31911));
    InMux I__6356 (
            .O(N__31925),
            .I(N__31908));
    InMux I__6355 (
            .O(N__31924),
            .I(N__31905));
    InMux I__6354 (
            .O(N__31923),
            .I(N__31896));
    InMux I__6353 (
            .O(N__31922),
            .I(N__31896));
    InMux I__6352 (
            .O(N__31921),
            .I(N__31896));
    InMux I__6351 (
            .O(N__31920),
            .I(N__31896));
    InMux I__6350 (
            .O(N__31919),
            .I(N__31893));
    InMux I__6349 (
            .O(N__31918),
            .I(N__31888));
    InMux I__6348 (
            .O(N__31917),
            .I(N__31888));
    LocalMux I__6347 (
            .O(N__31914),
            .I(N__31885));
    Span4Mux_h I__6346 (
            .O(N__31911),
            .I(N__31880));
    LocalMux I__6345 (
            .O(N__31908),
            .I(N__31880));
    LocalMux I__6344 (
            .O(N__31905),
            .I(N__31874));
    LocalMux I__6343 (
            .O(N__31896),
            .I(N__31867));
    LocalMux I__6342 (
            .O(N__31893),
            .I(N__31867));
    LocalMux I__6341 (
            .O(N__31888),
            .I(N__31867));
    Span4Mux_v I__6340 (
            .O(N__31885),
            .I(N__31864));
    Sp12to4 I__6339 (
            .O(N__31880),
            .I(N__31861));
    InMux I__6338 (
            .O(N__31879),
            .I(N__31856));
    InMux I__6337 (
            .O(N__31878),
            .I(N__31856));
    InMux I__6336 (
            .O(N__31877),
            .I(N__31853));
    Span4Mux_v I__6335 (
            .O(N__31874),
            .I(N__31848));
    Span4Mux_v I__6334 (
            .O(N__31867),
            .I(N__31848));
    Sp12to4 I__6333 (
            .O(N__31864),
            .I(N__31839));
    Span12Mux_v I__6332 (
            .O(N__31861),
            .I(N__31839));
    LocalMux I__6331 (
            .O(N__31856),
            .I(N__31839));
    LocalMux I__6330 (
            .O(N__31853),
            .I(N__31839));
    Odrv4 I__6329 (
            .O(N__31848),
            .I(\c0.n8 ));
    Odrv12 I__6328 (
            .O(N__31839),
            .I(\c0.n8 ));
    CascadeMux I__6327 (
            .O(N__31834),
            .I(N__31831));
    InMux I__6326 (
            .O(N__31831),
            .I(N__31827));
    CascadeMux I__6325 (
            .O(N__31830),
            .I(N__31823));
    LocalMux I__6324 (
            .O(N__31827),
            .I(N__31820));
    CascadeMux I__6323 (
            .O(N__31826),
            .I(N__31816));
    InMux I__6322 (
            .O(N__31823),
            .I(N__31813));
    Span4Mux_h I__6321 (
            .O(N__31820),
            .I(N__31809));
    InMux I__6320 (
            .O(N__31819),
            .I(N__31804));
    InMux I__6319 (
            .O(N__31816),
            .I(N__31804));
    LocalMux I__6318 (
            .O(N__31813),
            .I(N__31801));
    InMux I__6317 (
            .O(N__31812),
            .I(N__31798));
    Span4Mux_h I__6316 (
            .O(N__31809),
            .I(N__31789));
    LocalMux I__6315 (
            .O(N__31804),
            .I(N__31789));
    Sp12to4 I__6314 (
            .O(N__31801),
            .I(N__31784));
    LocalMux I__6313 (
            .O(N__31798),
            .I(N__31784));
    InMux I__6312 (
            .O(N__31797),
            .I(N__31781));
    InMux I__6311 (
            .O(N__31796),
            .I(N__31778));
    InMux I__6310 (
            .O(N__31795),
            .I(N__31775));
    InMux I__6309 (
            .O(N__31794),
            .I(N__31772));
    Odrv4 I__6308 (
            .O(N__31789),
            .I(rx_data_4));
    Odrv12 I__6307 (
            .O(N__31784),
            .I(rx_data_4));
    LocalMux I__6306 (
            .O(N__31781),
            .I(rx_data_4));
    LocalMux I__6305 (
            .O(N__31778),
            .I(rx_data_4));
    LocalMux I__6304 (
            .O(N__31775),
            .I(rx_data_4));
    LocalMux I__6303 (
            .O(N__31772),
            .I(rx_data_4));
    CascadeMux I__6302 (
            .O(N__31759),
            .I(N__31755));
    InMux I__6301 (
            .O(N__31758),
            .I(N__31752));
    InMux I__6300 (
            .O(N__31755),
            .I(N__31749));
    LocalMux I__6299 (
            .O(N__31752),
            .I(N__31744));
    LocalMux I__6298 (
            .O(N__31749),
            .I(N__31744));
    Odrv4 I__6297 (
            .O(N__31744),
            .I(\c0.data_in_frame_2_4 ));
    InMux I__6296 (
            .O(N__31741),
            .I(N__31738));
    LocalMux I__6295 (
            .O(N__31738),
            .I(N__31732));
    CascadeMux I__6294 (
            .O(N__31737),
            .I(N__31729));
    InMux I__6293 (
            .O(N__31736),
            .I(N__31725));
    InMux I__6292 (
            .O(N__31735),
            .I(N__31722));
    Span4Mux_v I__6291 (
            .O(N__31732),
            .I(N__31718));
    InMux I__6290 (
            .O(N__31729),
            .I(N__31715));
    InMux I__6289 (
            .O(N__31728),
            .I(N__31712));
    LocalMux I__6288 (
            .O(N__31725),
            .I(N__31707));
    LocalMux I__6287 (
            .O(N__31722),
            .I(N__31707));
    CascadeMux I__6286 (
            .O(N__31721),
            .I(N__31703));
    Span4Mux_h I__6285 (
            .O(N__31718),
            .I(N__31698));
    LocalMux I__6284 (
            .O(N__31715),
            .I(N__31698));
    LocalMux I__6283 (
            .O(N__31712),
            .I(N__31695));
    Span4Mux_h I__6282 (
            .O(N__31707),
            .I(N__31692));
    InMux I__6281 (
            .O(N__31706),
            .I(N__31687));
    InMux I__6280 (
            .O(N__31703),
            .I(N__31687));
    Span4Mux_h I__6279 (
            .O(N__31698),
            .I(N__31684));
    Span12Mux_v I__6278 (
            .O(N__31695),
            .I(N__31681));
    Odrv4 I__6277 (
            .O(N__31692),
            .I(\c0.r_SM_Main_2_N_2036_0 ));
    LocalMux I__6276 (
            .O(N__31687),
            .I(\c0.r_SM_Main_2_N_2036_0 ));
    Odrv4 I__6275 (
            .O(N__31684),
            .I(\c0.r_SM_Main_2_N_2036_0 ));
    Odrv12 I__6274 (
            .O(N__31681),
            .I(\c0.r_SM_Main_2_N_2036_0 ));
    InMux I__6273 (
            .O(N__31672),
            .I(N__31667));
    InMux I__6272 (
            .O(N__31671),
            .I(N__31664));
    InMux I__6271 (
            .O(N__31670),
            .I(N__31661));
    LocalMux I__6270 (
            .O(N__31667),
            .I(N__31657));
    LocalMux I__6269 (
            .O(N__31664),
            .I(N__31654));
    LocalMux I__6268 (
            .O(N__31661),
            .I(N__31651));
    InMux I__6267 (
            .O(N__31660),
            .I(N__31648));
    Span4Mux_v I__6266 (
            .O(N__31657),
            .I(N__31645));
    Span4Mux_h I__6265 (
            .O(N__31654),
            .I(N__31639));
    Span4Mux_h I__6264 (
            .O(N__31651),
            .I(N__31636));
    LocalMux I__6263 (
            .O(N__31648),
            .I(N__31633));
    Span4Mux_h I__6262 (
            .O(N__31645),
            .I(N__31630));
    InMux I__6261 (
            .O(N__31644),
            .I(N__31623));
    InMux I__6260 (
            .O(N__31643),
            .I(N__31623));
    InMux I__6259 (
            .O(N__31642),
            .I(N__31623));
    Odrv4 I__6258 (
            .O(N__31639),
            .I(tx_active));
    Odrv4 I__6257 (
            .O(N__31636),
            .I(tx_active));
    Odrv4 I__6256 (
            .O(N__31633),
            .I(tx_active));
    Odrv4 I__6255 (
            .O(N__31630),
            .I(tx_active));
    LocalMux I__6254 (
            .O(N__31623),
            .I(tx_active));
    CascadeMux I__6253 (
            .O(N__31612),
            .I(N__31609));
    InMux I__6252 (
            .O(N__31609),
            .I(N__31605));
    CascadeMux I__6251 (
            .O(N__31608),
            .I(N__31602));
    LocalMux I__6250 (
            .O(N__31605),
            .I(N__31598));
    InMux I__6249 (
            .O(N__31602),
            .I(N__31595));
    InMux I__6248 (
            .O(N__31601),
            .I(N__31592));
    Span4Mux_s2_v I__6247 (
            .O(N__31598),
            .I(N__31589));
    LocalMux I__6246 (
            .O(N__31595),
            .I(N__31584));
    LocalMux I__6245 (
            .O(N__31592),
            .I(N__31584));
    Span4Mux_h I__6244 (
            .O(N__31589),
            .I(N__31579));
    Span4Mux_s2_v I__6243 (
            .O(N__31584),
            .I(N__31579));
    Span4Mux_h I__6242 (
            .O(N__31579),
            .I(N__31576));
    Odrv4 I__6241 (
            .O(N__31576),
            .I(n17230));
    InMux I__6240 (
            .O(N__31573),
            .I(N__31567));
    InMux I__6239 (
            .O(N__31572),
            .I(N__31567));
    LocalMux I__6238 (
            .O(N__31567),
            .I(data_out_1_7));
    InMux I__6237 (
            .O(N__31564),
            .I(N__31561));
    LocalMux I__6236 (
            .O(N__31561),
            .I(N__31558));
    Span4Mux_h I__6235 (
            .O(N__31558),
            .I(N__31555));
    Odrv4 I__6234 (
            .O(N__31555),
            .I(\c0.n10 ));
    InMux I__6233 (
            .O(N__31552),
            .I(N__31547));
    InMux I__6232 (
            .O(N__31551),
            .I(N__31542));
    InMux I__6231 (
            .O(N__31550),
            .I(N__31539));
    LocalMux I__6230 (
            .O(N__31547),
            .I(N__31536));
    CascadeMux I__6229 (
            .O(N__31546),
            .I(N__31533));
    InMux I__6228 (
            .O(N__31545),
            .I(N__31529));
    LocalMux I__6227 (
            .O(N__31542),
            .I(N__31526));
    LocalMux I__6226 (
            .O(N__31539),
            .I(N__31521));
    Span4Mux_v I__6225 (
            .O(N__31536),
            .I(N__31518));
    InMux I__6224 (
            .O(N__31533),
            .I(N__31515));
    InMux I__6223 (
            .O(N__31532),
            .I(N__31510));
    LocalMux I__6222 (
            .O(N__31529),
            .I(N__31505));
    Span4Mux_v I__6221 (
            .O(N__31526),
            .I(N__31505));
    InMux I__6220 (
            .O(N__31525),
            .I(N__31500));
    InMux I__6219 (
            .O(N__31524),
            .I(N__31500));
    Span4Mux_v I__6218 (
            .O(N__31521),
            .I(N__31489));
    Span4Mux_h I__6217 (
            .O(N__31518),
            .I(N__31489));
    LocalMux I__6216 (
            .O(N__31515),
            .I(N__31489));
    CascadeMux I__6215 (
            .O(N__31514),
            .I(N__31482));
    InMux I__6214 (
            .O(N__31513),
            .I(N__31478));
    LocalMux I__6213 (
            .O(N__31510),
            .I(N__31475));
    Span4Mux_h I__6212 (
            .O(N__31505),
            .I(N__31470));
    LocalMux I__6211 (
            .O(N__31500),
            .I(N__31470));
    InMux I__6210 (
            .O(N__31499),
            .I(N__31467));
    InMux I__6209 (
            .O(N__31498),
            .I(N__31462));
    InMux I__6208 (
            .O(N__31497),
            .I(N__31462));
    InMux I__6207 (
            .O(N__31496),
            .I(N__31459));
    Span4Mux_h I__6206 (
            .O(N__31489),
            .I(N__31456));
    InMux I__6205 (
            .O(N__31488),
            .I(N__31449));
    InMux I__6204 (
            .O(N__31487),
            .I(N__31449));
    InMux I__6203 (
            .O(N__31486),
            .I(N__31449));
    InMux I__6202 (
            .O(N__31485),
            .I(N__31442));
    InMux I__6201 (
            .O(N__31482),
            .I(N__31442));
    InMux I__6200 (
            .O(N__31481),
            .I(N__31442));
    LocalMux I__6199 (
            .O(N__31478),
            .I(N__31435));
    Span4Mux_s1_h I__6198 (
            .O(N__31475),
            .I(N__31435));
    Span4Mux_h I__6197 (
            .O(N__31470),
            .I(N__31435));
    LocalMux I__6196 (
            .O(N__31467),
            .I(r_SM_Main_2_adj_2443));
    LocalMux I__6195 (
            .O(N__31462),
            .I(r_SM_Main_2_adj_2443));
    LocalMux I__6194 (
            .O(N__31459),
            .I(r_SM_Main_2_adj_2443));
    Odrv4 I__6193 (
            .O(N__31456),
            .I(r_SM_Main_2_adj_2443));
    LocalMux I__6192 (
            .O(N__31449),
            .I(r_SM_Main_2_adj_2443));
    LocalMux I__6191 (
            .O(N__31442),
            .I(r_SM_Main_2_adj_2443));
    Odrv4 I__6190 (
            .O(N__31435),
            .I(r_SM_Main_2_adj_2443));
    InMux I__6189 (
            .O(N__31420),
            .I(N__31417));
    LocalMux I__6188 (
            .O(N__31417),
            .I(N__31414));
    Span12Mux_h I__6187 (
            .O(N__31414),
            .I(N__31411));
    Odrv12 I__6186 (
            .O(N__31411),
            .I(n17544));
    CascadeMux I__6185 (
            .O(N__31408),
            .I(N__31404));
    InMux I__6184 (
            .O(N__31407),
            .I(N__31400));
    InMux I__6183 (
            .O(N__31404),
            .I(N__31397));
    InMux I__6182 (
            .O(N__31403),
            .I(N__31394));
    LocalMux I__6181 (
            .O(N__31400),
            .I(N__31389));
    LocalMux I__6180 (
            .O(N__31397),
            .I(N__31389));
    LocalMux I__6179 (
            .O(N__31394),
            .I(r_Clock_Count_0_adj_2454));
    Odrv12 I__6178 (
            .O(N__31389),
            .I(r_Clock_Count_0_adj_2454));
    CascadeMux I__6177 (
            .O(N__31384),
            .I(N__31380));
    InMux I__6176 (
            .O(N__31383),
            .I(N__31374));
    InMux I__6175 (
            .O(N__31380),
            .I(N__31371));
    InMux I__6174 (
            .O(N__31379),
            .I(N__31368));
    InMux I__6173 (
            .O(N__31378),
            .I(N__31365));
    InMux I__6172 (
            .O(N__31377),
            .I(N__31362));
    LocalMux I__6171 (
            .O(N__31374),
            .I(N__31356));
    LocalMux I__6170 (
            .O(N__31371),
            .I(N__31356));
    LocalMux I__6169 (
            .O(N__31368),
            .I(N__31353));
    LocalMux I__6168 (
            .O(N__31365),
            .I(N__31350));
    LocalMux I__6167 (
            .O(N__31362),
            .I(N__31347));
    CascadeMux I__6166 (
            .O(N__31361),
            .I(N__31344));
    Span4Mux_v I__6165 (
            .O(N__31356),
            .I(N__31338));
    Span4Mux_v I__6164 (
            .O(N__31353),
            .I(N__31338));
    Span4Mux_v I__6163 (
            .O(N__31350),
            .I(N__31333));
    Span4Mux_v I__6162 (
            .O(N__31347),
            .I(N__31333));
    InMux I__6161 (
            .O(N__31344),
            .I(N__31330));
    InMux I__6160 (
            .O(N__31343),
            .I(N__31327));
    Sp12to4 I__6159 (
            .O(N__31338),
            .I(N__31322));
    Sp12to4 I__6158 (
            .O(N__31333),
            .I(N__31322));
    LocalMux I__6157 (
            .O(N__31330),
            .I(r_Bit_Index_1));
    LocalMux I__6156 (
            .O(N__31327),
            .I(r_Bit_Index_1));
    Odrv12 I__6155 (
            .O(N__31322),
            .I(r_Bit_Index_1));
    InMux I__6154 (
            .O(N__31315),
            .I(N__31312));
    LocalMux I__6153 (
            .O(N__31312),
            .I(N__31309));
    Span4Mux_h I__6152 (
            .O(N__31309),
            .I(N__31306));
    Odrv4 I__6151 (
            .O(N__31306),
            .I(n17398));
    CascadeMux I__6150 (
            .O(N__31303),
            .I(\c0.n17918_cascade_ ));
    InMux I__6149 (
            .O(N__31300),
            .I(N__31297));
    LocalMux I__6148 (
            .O(N__31297),
            .I(\c0.n17343 ));
    InMux I__6147 (
            .O(N__31294),
            .I(N__31288));
    InMux I__6146 (
            .O(N__31293),
            .I(N__31288));
    LocalMux I__6145 (
            .O(N__31288),
            .I(N__31285));
    Span4Mux_h I__6144 (
            .O(N__31285),
            .I(N__31281));
    InMux I__6143 (
            .O(N__31284),
            .I(N__31278));
    Odrv4 I__6142 (
            .O(N__31281),
            .I(\c0.n17769 ));
    LocalMux I__6141 (
            .O(N__31278),
            .I(\c0.n17769 ));
    InMux I__6140 (
            .O(N__31273),
            .I(N__31270));
    LocalMux I__6139 (
            .O(N__31270),
            .I(N__31267));
    Span4Mux_h I__6138 (
            .O(N__31267),
            .I(N__31264));
    Odrv4 I__6137 (
            .O(N__31264),
            .I(\c0.n18 ));
    InMux I__6136 (
            .O(N__31261),
            .I(N__31258));
    LocalMux I__6135 (
            .O(N__31258),
            .I(N__31255));
    Span4Mux_h I__6134 (
            .O(N__31255),
            .I(N__31252));
    Odrv4 I__6133 (
            .O(N__31252),
            .I(\c0.n17 ));
    CascadeMux I__6132 (
            .O(N__31249),
            .I(N__31246));
    InMux I__6131 (
            .O(N__31246),
            .I(N__31243));
    LocalMux I__6130 (
            .O(N__31243),
            .I(\c0.n26_adj_2147 ));
    InMux I__6129 (
            .O(N__31240),
            .I(N__31237));
    LocalMux I__6128 (
            .O(N__31237),
            .I(N__31234));
    Odrv4 I__6127 (
            .O(N__31234),
            .I(\c0.n30_adj_2148 ));
    CascadeMux I__6126 (
            .O(N__31231),
            .I(N__31225));
    CascadeMux I__6125 (
            .O(N__31230),
            .I(N__31222));
    CascadeMux I__6124 (
            .O(N__31229),
            .I(N__31218));
    InMux I__6123 (
            .O(N__31228),
            .I(N__31213));
    InMux I__6122 (
            .O(N__31225),
            .I(N__31209));
    InMux I__6121 (
            .O(N__31222),
            .I(N__31206));
    InMux I__6120 (
            .O(N__31221),
            .I(N__31203));
    InMux I__6119 (
            .O(N__31218),
            .I(N__31199));
    InMux I__6118 (
            .O(N__31217),
            .I(N__31194));
    InMux I__6117 (
            .O(N__31216),
            .I(N__31194));
    LocalMux I__6116 (
            .O(N__31213),
            .I(N__31191));
    InMux I__6115 (
            .O(N__31212),
            .I(N__31188));
    LocalMux I__6114 (
            .O(N__31209),
            .I(N__31181));
    LocalMux I__6113 (
            .O(N__31206),
            .I(N__31181));
    LocalMux I__6112 (
            .O(N__31203),
            .I(N__31181));
    CascadeMux I__6111 (
            .O(N__31202),
            .I(N__31178));
    LocalMux I__6110 (
            .O(N__31199),
            .I(N__31175));
    LocalMux I__6109 (
            .O(N__31194),
            .I(N__31172));
    Span4Mux_v I__6108 (
            .O(N__31191),
            .I(N__31169));
    LocalMux I__6107 (
            .O(N__31188),
            .I(N__31164));
    Span4Mux_h I__6106 (
            .O(N__31181),
            .I(N__31164));
    InMux I__6105 (
            .O(N__31178),
            .I(N__31161));
    Span4Mux_v I__6104 (
            .O(N__31175),
            .I(N__31158));
    Span4Mux_h I__6103 (
            .O(N__31172),
            .I(N__31155));
    Span4Mux_v I__6102 (
            .O(N__31169),
            .I(N__31150));
    Span4Mux_h I__6101 (
            .O(N__31164),
            .I(N__31150));
    LocalMux I__6100 (
            .O(N__31161),
            .I(rx_data_5));
    Odrv4 I__6099 (
            .O(N__31158),
            .I(rx_data_5));
    Odrv4 I__6098 (
            .O(N__31155),
            .I(rx_data_5));
    Odrv4 I__6097 (
            .O(N__31150),
            .I(rx_data_5));
    InMux I__6096 (
            .O(N__31141),
            .I(N__31138));
    LocalMux I__6095 (
            .O(N__31138),
            .I(N__31130));
    InMux I__6094 (
            .O(N__31137),
            .I(N__31127));
    InMux I__6093 (
            .O(N__31136),
            .I(N__31124));
    InMux I__6092 (
            .O(N__31135),
            .I(N__31121));
    InMux I__6091 (
            .O(N__31134),
            .I(N__31116));
    InMux I__6090 (
            .O(N__31133),
            .I(N__31116));
    Span4Mux_h I__6089 (
            .O(N__31130),
            .I(N__31104));
    LocalMux I__6088 (
            .O(N__31127),
            .I(N__31095));
    LocalMux I__6087 (
            .O(N__31124),
            .I(N__31095));
    LocalMux I__6086 (
            .O(N__31121),
            .I(N__31095));
    LocalMux I__6085 (
            .O(N__31116),
            .I(N__31095));
    InMux I__6084 (
            .O(N__31115),
            .I(N__31092));
    InMux I__6083 (
            .O(N__31114),
            .I(N__31089));
    InMux I__6082 (
            .O(N__31113),
            .I(N__31086));
    InMux I__6081 (
            .O(N__31112),
            .I(N__31079));
    InMux I__6080 (
            .O(N__31111),
            .I(N__31079));
    InMux I__6079 (
            .O(N__31110),
            .I(N__31079));
    InMux I__6078 (
            .O(N__31109),
            .I(N__31072));
    InMux I__6077 (
            .O(N__31108),
            .I(N__31072));
    InMux I__6076 (
            .O(N__31107),
            .I(N__31072));
    Odrv4 I__6075 (
            .O(N__31104),
            .I(\c0.n16882 ));
    Odrv12 I__6074 (
            .O(N__31095),
            .I(\c0.n16882 ));
    LocalMux I__6073 (
            .O(N__31092),
            .I(\c0.n16882 ));
    LocalMux I__6072 (
            .O(N__31089),
            .I(\c0.n16882 ));
    LocalMux I__6071 (
            .O(N__31086),
            .I(\c0.n16882 ));
    LocalMux I__6070 (
            .O(N__31079),
            .I(\c0.n16882 ));
    LocalMux I__6069 (
            .O(N__31072),
            .I(\c0.n16882 ));
    CascadeMux I__6068 (
            .O(N__31057),
            .I(N__31054));
    InMux I__6067 (
            .O(N__31054),
            .I(N__31050));
    InMux I__6066 (
            .O(N__31053),
            .I(N__31047));
    LocalMux I__6065 (
            .O(N__31050),
            .I(N__31044));
    LocalMux I__6064 (
            .O(N__31047),
            .I(\c0.data_in_frame_10_5 ));
    Odrv4 I__6063 (
            .O(N__31044),
            .I(\c0.data_in_frame_10_5 ));
    InMux I__6062 (
            .O(N__31039),
            .I(N__31035));
    InMux I__6061 (
            .O(N__31038),
            .I(N__31032));
    LocalMux I__6060 (
            .O(N__31035),
            .I(N__31029));
    LocalMux I__6059 (
            .O(N__31032),
            .I(N__31023));
    Span4Mux_v I__6058 (
            .O(N__31029),
            .I(N__31018));
    InMux I__6057 (
            .O(N__31028),
            .I(N__31015));
    InMux I__6056 (
            .O(N__31027),
            .I(N__31010));
    InMux I__6055 (
            .O(N__31026),
            .I(N__31007));
    Span4Mux_v I__6054 (
            .O(N__31023),
            .I(N__31004));
    InMux I__6053 (
            .O(N__31022),
            .I(N__31001));
    CascadeMux I__6052 (
            .O(N__31021),
            .I(N__30998));
    Span4Mux_h I__6051 (
            .O(N__31018),
            .I(N__30989));
    LocalMux I__6050 (
            .O(N__31015),
            .I(N__30989));
    InMux I__6049 (
            .O(N__31014),
            .I(N__30986));
    InMux I__6048 (
            .O(N__31013),
            .I(N__30983));
    LocalMux I__6047 (
            .O(N__31010),
            .I(N__30974));
    LocalMux I__6046 (
            .O(N__31007),
            .I(N__30974));
    Sp12to4 I__6045 (
            .O(N__31004),
            .I(N__30974));
    LocalMux I__6044 (
            .O(N__31001),
            .I(N__30974));
    InMux I__6043 (
            .O(N__30998),
            .I(N__30969));
    InMux I__6042 (
            .O(N__30997),
            .I(N__30969));
    InMux I__6041 (
            .O(N__30996),
            .I(N__30964));
    InMux I__6040 (
            .O(N__30995),
            .I(N__30964));
    InMux I__6039 (
            .O(N__30994),
            .I(N__30961));
    Span4Mux_h I__6038 (
            .O(N__30989),
            .I(N__30958));
    LocalMux I__6037 (
            .O(N__30986),
            .I(r_SM_Main_1_adj_2444));
    LocalMux I__6036 (
            .O(N__30983),
            .I(r_SM_Main_1_adj_2444));
    Odrv12 I__6035 (
            .O(N__30974),
            .I(r_SM_Main_1_adj_2444));
    LocalMux I__6034 (
            .O(N__30969),
            .I(r_SM_Main_1_adj_2444));
    LocalMux I__6033 (
            .O(N__30964),
            .I(r_SM_Main_1_adj_2444));
    LocalMux I__6032 (
            .O(N__30961),
            .I(r_SM_Main_1_adj_2444));
    Odrv4 I__6031 (
            .O(N__30958),
            .I(r_SM_Main_1_adj_2444));
    CascadeMux I__6030 (
            .O(N__30943),
            .I(N__30940));
    InMux I__6029 (
            .O(N__30940),
            .I(N__30937));
    LocalMux I__6028 (
            .O(N__30937),
            .I(N__30934));
    Span4Mux_h I__6027 (
            .O(N__30934),
            .I(N__30931));
    Span4Mux_h I__6026 (
            .O(N__30931),
            .I(N__30928));
    Odrv4 I__6025 (
            .O(N__30928),
            .I(\c0.tx2.n6480 ));
    InMux I__6024 (
            .O(N__30925),
            .I(N__30922));
    LocalMux I__6023 (
            .O(N__30922),
            .I(N__30919));
    Span4Mux_h I__6022 (
            .O(N__30919),
            .I(N__30916));
    Span4Mux_h I__6021 (
            .O(N__30916),
            .I(N__30913));
    Odrv4 I__6020 (
            .O(N__30913),
            .I(\c0.tx2.n1 ));
    InMux I__6019 (
            .O(N__30910),
            .I(N__30907));
    LocalMux I__6018 (
            .O(N__30907),
            .I(N__30904));
    Odrv4 I__6017 (
            .O(N__30904),
            .I(\c0.tx2.n10101 ));
    InMux I__6016 (
            .O(N__30901),
            .I(N__30898));
    LocalMux I__6015 (
            .O(N__30898),
            .I(N__30894));
    InMux I__6014 (
            .O(N__30897),
            .I(N__30891));
    Span4Mux_h I__6013 (
            .O(N__30894),
            .I(N__30888));
    LocalMux I__6012 (
            .O(N__30891),
            .I(data_out_frame2_18_5));
    Odrv4 I__6011 (
            .O(N__30888),
            .I(data_out_frame2_18_5));
    InMux I__6010 (
            .O(N__30883),
            .I(N__30880));
    LocalMux I__6009 (
            .O(N__30880),
            .I(N__30877));
    Span4Mux_h I__6008 (
            .O(N__30877),
            .I(N__30871));
    InMux I__6007 (
            .O(N__30876),
            .I(N__30868));
    InMux I__6006 (
            .O(N__30875),
            .I(N__30865));
    InMux I__6005 (
            .O(N__30874),
            .I(N__30861));
    Span4Mux_h I__6004 (
            .O(N__30871),
            .I(N__30854));
    LocalMux I__6003 (
            .O(N__30868),
            .I(N__30854));
    LocalMux I__6002 (
            .O(N__30865),
            .I(N__30854));
    InMux I__6001 (
            .O(N__30864),
            .I(N__30849));
    LocalMux I__6000 (
            .O(N__30861),
            .I(N__30845));
    Span4Mux_h I__5999 (
            .O(N__30854),
            .I(N__30842));
    InMux I__5998 (
            .O(N__30853),
            .I(N__30837));
    InMux I__5997 (
            .O(N__30852),
            .I(N__30837));
    LocalMux I__5996 (
            .O(N__30849),
            .I(N__30834));
    InMux I__5995 (
            .O(N__30848),
            .I(N__30831));
    Span4Mux_v I__5994 (
            .O(N__30845),
            .I(N__30827));
    Span4Mux_v I__5993 (
            .O(N__30842),
            .I(N__30824));
    LocalMux I__5992 (
            .O(N__30837),
            .I(N__30821));
    Span4Mux_h I__5991 (
            .O(N__30834),
            .I(N__30816));
    LocalMux I__5990 (
            .O(N__30831),
            .I(N__30816));
    InMux I__5989 (
            .O(N__30830),
            .I(N__30813));
    Odrv4 I__5988 (
            .O(N__30827),
            .I(r_SM_Main_2_adj_2439));
    Odrv4 I__5987 (
            .O(N__30824),
            .I(r_SM_Main_2_adj_2439));
    Odrv12 I__5986 (
            .O(N__30821),
            .I(r_SM_Main_2_adj_2439));
    Odrv4 I__5985 (
            .O(N__30816),
            .I(r_SM_Main_2_adj_2439));
    LocalMux I__5984 (
            .O(N__30813),
            .I(r_SM_Main_2_adj_2439));
    InMux I__5983 (
            .O(N__30802),
            .I(N__30799));
    LocalMux I__5982 (
            .O(N__30799),
            .I(N__30796));
    Span4Mux_v I__5981 (
            .O(N__30796),
            .I(N__30793));
    Span4Mux_h I__5980 (
            .O(N__30793),
            .I(N__30790));
    Odrv4 I__5979 (
            .O(N__30790),
            .I(n13440));
    CascadeMux I__5978 (
            .O(N__30787),
            .I(N__30784));
    InMux I__5977 (
            .O(N__30784),
            .I(N__30781));
    LocalMux I__5976 (
            .O(N__30781),
            .I(N__30776));
    InMux I__5975 (
            .O(N__30780),
            .I(N__30771));
    InMux I__5974 (
            .O(N__30779),
            .I(N__30771));
    Span4Mux_v I__5973 (
            .O(N__30776),
            .I(N__30765));
    LocalMux I__5972 (
            .O(N__30771),
            .I(N__30762));
    InMux I__5971 (
            .O(N__30770),
            .I(N__30756));
    InMux I__5970 (
            .O(N__30769),
            .I(N__30753));
    CascadeMux I__5969 (
            .O(N__30768),
            .I(N__30750));
    Span4Mux_h I__5968 (
            .O(N__30765),
            .I(N__30744));
    Span4Mux_v I__5967 (
            .O(N__30762),
            .I(N__30744));
    InMux I__5966 (
            .O(N__30761),
            .I(N__30739));
    InMux I__5965 (
            .O(N__30760),
            .I(N__30739));
    InMux I__5964 (
            .O(N__30759),
            .I(N__30736));
    LocalMux I__5963 (
            .O(N__30756),
            .I(N__30730));
    LocalMux I__5962 (
            .O(N__30753),
            .I(N__30730));
    InMux I__5961 (
            .O(N__30750),
            .I(N__30727));
    InMux I__5960 (
            .O(N__30749),
            .I(N__30724));
    Sp12to4 I__5959 (
            .O(N__30744),
            .I(N__30721));
    LocalMux I__5958 (
            .O(N__30739),
            .I(N__30716));
    LocalMux I__5957 (
            .O(N__30736),
            .I(N__30716));
    InMux I__5956 (
            .O(N__30735),
            .I(N__30713));
    Span4Mux_s2_h I__5955 (
            .O(N__30730),
            .I(N__30710));
    LocalMux I__5954 (
            .O(N__30727),
            .I(r_SM_Main_1_adj_2440));
    LocalMux I__5953 (
            .O(N__30724),
            .I(r_SM_Main_1_adj_2440));
    Odrv12 I__5952 (
            .O(N__30721),
            .I(r_SM_Main_1_adj_2440));
    Odrv4 I__5951 (
            .O(N__30716),
            .I(r_SM_Main_1_adj_2440));
    LocalMux I__5950 (
            .O(N__30713),
            .I(r_SM_Main_1_adj_2440));
    Odrv4 I__5949 (
            .O(N__30710),
            .I(r_SM_Main_1_adj_2440));
    InMux I__5948 (
            .O(N__30697),
            .I(N__30690));
    InMux I__5947 (
            .O(N__30696),
            .I(N__30687));
    InMux I__5946 (
            .O(N__30695),
            .I(N__30684));
    CascadeMux I__5945 (
            .O(N__30694),
            .I(N__30680));
    CascadeMux I__5944 (
            .O(N__30693),
            .I(N__30676));
    LocalMux I__5943 (
            .O(N__30690),
            .I(N__30669));
    LocalMux I__5942 (
            .O(N__30687),
            .I(N__30669));
    LocalMux I__5941 (
            .O(N__30684),
            .I(N__30669));
    InMux I__5940 (
            .O(N__30683),
            .I(N__30666));
    InMux I__5939 (
            .O(N__30680),
            .I(N__30662));
    InMux I__5938 (
            .O(N__30679),
            .I(N__30659));
    InMux I__5937 (
            .O(N__30676),
            .I(N__30656));
    Span4Mux_v I__5936 (
            .O(N__30669),
            .I(N__30653));
    LocalMux I__5935 (
            .O(N__30666),
            .I(N__30650));
    CascadeMux I__5934 (
            .O(N__30665),
            .I(N__30646));
    LocalMux I__5933 (
            .O(N__30662),
            .I(N__30639));
    LocalMux I__5932 (
            .O(N__30659),
            .I(N__30639));
    LocalMux I__5931 (
            .O(N__30656),
            .I(N__30639));
    Span4Mux_h I__5930 (
            .O(N__30653),
            .I(N__30636));
    Span4Mux_v I__5929 (
            .O(N__30650),
            .I(N__30633));
    InMux I__5928 (
            .O(N__30649),
            .I(N__30628));
    InMux I__5927 (
            .O(N__30646),
            .I(N__30628));
    Odrv12 I__5926 (
            .O(N__30639),
            .I(rx_data_1));
    Odrv4 I__5925 (
            .O(N__30636),
            .I(rx_data_1));
    Odrv4 I__5924 (
            .O(N__30633),
            .I(rx_data_1));
    LocalMux I__5923 (
            .O(N__30628),
            .I(rx_data_1));
    InMux I__5922 (
            .O(N__30619),
            .I(N__30615));
    InMux I__5921 (
            .O(N__30618),
            .I(N__30612));
    LocalMux I__5920 (
            .O(N__30615),
            .I(N__30609));
    LocalMux I__5919 (
            .O(N__30612),
            .I(\c0.data_in_frame_2_1 ));
    Odrv4 I__5918 (
            .O(N__30609),
            .I(\c0.data_in_frame_2_1 ));
    InMux I__5917 (
            .O(N__30604),
            .I(N__30598));
    InMux I__5916 (
            .O(N__30603),
            .I(N__30598));
    LocalMux I__5915 (
            .O(N__30598),
            .I(N__30594));
    InMux I__5914 (
            .O(N__30597),
            .I(N__30591));
    Sp12to4 I__5913 (
            .O(N__30594),
            .I(N__30588));
    LocalMux I__5912 (
            .O(N__30591),
            .I(\c0.tx2.tx2_active ));
    Odrv12 I__5911 (
            .O(N__30588),
            .I(\c0.tx2.tx2_active ));
    CascadeMux I__5910 (
            .O(N__30583),
            .I(\c0.n17334_cascade_ ));
    InMux I__5909 (
            .O(N__30580),
            .I(N__30576));
    InMux I__5908 (
            .O(N__30579),
            .I(N__30572));
    LocalMux I__5907 (
            .O(N__30576),
            .I(N__30569));
    InMux I__5906 (
            .O(N__30575),
            .I(N__30566));
    LocalMux I__5905 (
            .O(N__30572),
            .I(N__30563));
    Odrv12 I__5904 (
            .O(N__30569),
            .I(\c0.n2334 ));
    LocalMux I__5903 (
            .O(N__30566),
            .I(\c0.n2334 ));
    Odrv4 I__5902 (
            .O(N__30563),
            .I(\c0.n2334 ));
    InMux I__5901 (
            .O(N__30556),
            .I(N__30552));
    InMux I__5900 (
            .O(N__30555),
            .I(N__30549));
    LocalMux I__5899 (
            .O(N__30552),
            .I(N__30546));
    LocalMux I__5898 (
            .O(N__30549),
            .I(N__30543));
    Odrv4 I__5897 (
            .O(N__30546),
            .I(\c0.n2351 ));
    Odrv4 I__5896 (
            .O(N__30543),
            .I(\c0.n2351 ));
    InMux I__5895 (
            .O(N__30538),
            .I(N__30535));
    LocalMux I__5894 (
            .O(N__30535),
            .I(\c0.n18_adj_2343 ));
    CascadeMux I__5893 (
            .O(N__30532),
            .I(N__30528));
    CascadeMux I__5892 (
            .O(N__30531),
            .I(N__30525));
    InMux I__5891 (
            .O(N__30528),
            .I(N__30519));
    InMux I__5890 (
            .O(N__30525),
            .I(N__30516));
    InMux I__5889 (
            .O(N__30524),
            .I(N__30513));
    InMux I__5888 (
            .O(N__30523),
            .I(N__30509));
    InMux I__5887 (
            .O(N__30522),
            .I(N__30506));
    LocalMux I__5886 (
            .O(N__30519),
            .I(N__30500));
    LocalMux I__5885 (
            .O(N__30516),
            .I(N__30500));
    LocalMux I__5884 (
            .O(N__30513),
            .I(N__30497));
    InMux I__5883 (
            .O(N__30512),
            .I(N__30494));
    LocalMux I__5882 (
            .O(N__30509),
            .I(N__30489));
    LocalMux I__5881 (
            .O(N__30506),
            .I(N__30489));
    InMux I__5880 (
            .O(N__30505),
            .I(N__30484));
    Span4Mux_v I__5879 (
            .O(N__30500),
            .I(N__30479));
    Span4Mux_h I__5878 (
            .O(N__30497),
            .I(N__30479));
    LocalMux I__5877 (
            .O(N__30494),
            .I(N__30476));
    Span4Mux_v I__5876 (
            .O(N__30489),
            .I(N__30473));
    InMux I__5875 (
            .O(N__30488),
            .I(N__30470));
    CascadeMux I__5874 (
            .O(N__30487),
            .I(N__30467));
    LocalMux I__5873 (
            .O(N__30484),
            .I(N__30464));
    Span4Mux_h I__5872 (
            .O(N__30479),
            .I(N__30461));
    Span4Mux_v I__5871 (
            .O(N__30476),
            .I(N__30454));
    Span4Mux_s3_h I__5870 (
            .O(N__30473),
            .I(N__30454));
    LocalMux I__5869 (
            .O(N__30470),
            .I(N__30454));
    InMux I__5868 (
            .O(N__30467),
            .I(N__30451));
    Odrv12 I__5867 (
            .O(N__30464),
            .I(rx_data_3));
    Odrv4 I__5866 (
            .O(N__30461),
            .I(rx_data_3));
    Odrv4 I__5865 (
            .O(N__30454),
            .I(rx_data_3));
    LocalMux I__5864 (
            .O(N__30451),
            .I(rx_data_3));
    InMux I__5863 (
            .O(N__30442),
            .I(N__30438));
    InMux I__5862 (
            .O(N__30441),
            .I(N__30431));
    LocalMux I__5861 (
            .O(N__30438),
            .I(N__30428));
    InMux I__5860 (
            .O(N__30437),
            .I(N__30423));
    InMux I__5859 (
            .O(N__30436),
            .I(N__30423));
    InMux I__5858 (
            .O(N__30435),
            .I(N__30418));
    InMux I__5857 (
            .O(N__30434),
            .I(N__30415));
    LocalMux I__5856 (
            .O(N__30431),
            .I(N__30412));
    Span4Mux_h I__5855 (
            .O(N__30428),
            .I(N__30407));
    LocalMux I__5854 (
            .O(N__30423),
            .I(N__30407));
    InMux I__5853 (
            .O(N__30422),
            .I(N__30402));
    InMux I__5852 (
            .O(N__30421),
            .I(N__30402));
    LocalMux I__5851 (
            .O(N__30418),
            .I(N__30397));
    LocalMux I__5850 (
            .O(N__30415),
            .I(N__30397));
    Span4Mux_v I__5849 (
            .O(N__30412),
            .I(N__30390));
    Span4Mux_h I__5848 (
            .O(N__30407),
            .I(N__30390));
    LocalMux I__5847 (
            .O(N__30402),
            .I(N__30390));
    Span12Mux_s11_v I__5846 (
            .O(N__30397),
            .I(N__30387));
    Span4Mux_v I__5845 (
            .O(N__30390),
            .I(N__30384));
    Odrv12 I__5844 (
            .O(N__30387),
            .I(n16897));
    Odrv4 I__5843 (
            .O(N__30384),
            .I(n16897));
    InMux I__5842 (
            .O(N__30379),
            .I(N__30372));
    InMux I__5841 (
            .O(N__30378),
            .I(N__30372));
    InMux I__5840 (
            .O(N__30377),
            .I(N__30368));
    LocalMux I__5839 (
            .O(N__30372),
            .I(N__30365));
    InMux I__5838 (
            .O(N__30371),
            .I(N__30362));
    LocalMux I__5837 (
            .O(N__30368),
            .I(N__30359));
    Span4Mux_h I__5836 (
            .O(N__30365),
            .I(N__30356));
    LocalMux I__5835 (
            .O(N__30362),
            .I(data_in_frame_0_3));
    Odrv4 I__5834 (
            .O(N__30359),
            .I(data_in_frame_0_3));
    Odrv4 I__5833 (
            .O(N__30356),
            .I(data_in_frame_0_3));
    CascadeMux I__5832 (
            .O(N__30349),
            .I(\c0.n17337_cascade_ ));
    InMux I__5831 (
            .O(N__30346),
            .I(N__30343));
    LocalMux I__5830 (
            .O(N__30343),
            .I(N__30340));
    Span4Mux_v I__5829 (
            .O(N__30340),
            .I(N__30336));
    InMux I__5828 (
            .O(N__30339),
            .I(N__30331));
    Span4Mux_h I__5827 (
            .O(N__30336),
            .I(N__30328));
    InMux I__5826 (
            .O(N__30335),
            .I(N__30323));
    InMux I__5825 (
            .O(N__30334),
            .I(N__30323));
    LocalMux I__5824 (
            .O(N__30331),
            .I(data_in_frame_0_4));
    Odrv4 I__5823 (
            .O(N__30328),
            .I(data_in_frame_0_4));
    LocalMux I__5822 (
            .O(N__30323),
            .I(data_in_frame_0_4));
    InMux I__5821 (
            .O(N__30316),
            .I(N__30312));
    InMux I__5820 (
            .O(N__30315),
            .I(N__30309));
    LocalMux I__5819 (
            .O(N__30312),
            .I(N__30306));
    LocalMux I__5818 (
            .O(N__30309),
            .I(N__30301));
    Span4Mux_h I__5817 (
            .O(N__30306),
            .I(N__30296));
    InMux I__5816 (
            .O(N__30305),
            .I(N__30291));
    InMux I__5815 (
            .O(N__30304),
            .I(N__30291));
    Span4Mux_h I__5814 (
            .O(N__30301),
            .I(N__30288));
    InMux I__5813 (
            .O(N__30300),
            .I(N__30285));
    InMux I__5812 (
            .O(N__30299),
            .I(N__30282));
    Odrv4 I__5811 (
            .O(N__30296),
            .I(data_in_frame_0_5));
    LocalMux I__5810 (
            .O(N__30291),
            .I(data_in_frame_0_5));
    Odrv4 I__5809 (
            .O(N__30288),
            .I(data_in_frame_0_5));
    LocalMux I__5808 (
            .O(N__30285),
            .I(data_in_frame_0_5));
    LocalMux I__5807 (
            .O(N__30282),
            .I(data_in_frame_0_5));
    InMux I__5806 (
            .O(N__30271),
            .I(N__30268));
    LocalMux I__5805 (
            .O(N__30268),
            .I(N__30264));
    InMux I__5804 (
            .O(N__30267),
            .I(N__30261));
    Span4Mux_v I__5803 (
            .O(N__30264),
            .I(N__30258));
    LocalMux I__5802 (
            .O(N__30261),
            .I(N__30255));
    Span4Mux_h I__5801 (
            .O(N__30258),
            .I(N__30252));
    Span4Mux_v I__5800 (
            .O(N__30255),
            .I(N__30249));
    Odrv4 I__5799 (
            .O(N__30252),
            .I(\c0.n2338 ));
    Odrv4 I__5798 (
            .O(N__30249),
            .I(\c0.n2338 ));
    InMux I__5797 (
            .O(N__30244),
            .I(N__30241));
    LocalMux I__5796 (
            .O(N__30241),
            .I(N__30238));
    Span4Mux_h I__5795 (
            .O(N__30238),
            .I(N__30234));
    InMux I__5794 (
            .O(N__30237),
            .I(N__30231));
    Span4Mux_h I__5793 (
            .O(N__30234),
            .I(N__30228));
    LocalMux I__5792 (
            .O(N__30231),
            .I(\c0.data_in_frame_2_6 ));
    Odrv4 I__5791 (
            .O(N__30228),
            .I(\c0.data_in_frame_2_6 ));
    InMux I__5790 (
            .O(N__30223),
            .I(N__30220));
    LocalMux I__5789 (
            .O(N__30220),
            .I(N__30216));
    InMux I__5788 (
            .O(N__30219),
            .I(N__30213));
    Span4Mux_h I__5787 (
            .O(N__30216),
            .I(N__30210));
    LocalMux I__5786 (
            .O(N__30213),
            .I(N__30207));
    Span4Mux_h I__5785 (
            .O(N__30210),
            .I(N__30204));
    Odrv4 I__5784 (
            .O(N__30207),
            .I(\c0.data_in_frame_2_0 ));
    Odrv4 I__5783 (
            .O(N__30204),
            .I(\c0.data_in_frame_2_0 ));
    CascadeMux I__5782 (
            .O(N__30199),
            .I(\c0.n2338_cascade_ ));
    InMux I__5781 (
            .O(N__30196),
            .I(N__30193));
    LocalMux I__5780 (
            .O(N__30193),
            .I(N__30188));
    InMux I__5779 (
            .O(N__30192),
            .I(N__30185));
    InMux I__5778 (
            .O(N__30191),
            .I(N__30182));
    Span4Mux_v I__5777 (
            .O(N__30188),
            .I(N__30177));
    LocalMux I__5776 (
            .O(N__30185),
            .I(N__30177));
    LocalMux I__5775 (
            .O(N__30182),
            .I(\c0.n2352 ));
    Odrv4 I__5774 (
            .O(N__30177),
            .I(\c0.n2352 ));
    InMux I__5773 (
            .O(N__30172),
            .I(N__30169));
    LocalMux I__5772 (
            .O(N__30169),
            .I(N__30166));
    Span4Mux_h I__5771 (
            .O(N__30166),
            .I(N__30163));
    Odrv4 I__5770 (
            .O(N__30163),
            .I(\c0.n26_adj_2344 ));
    CascadeMux I__5769 (
            .O(N__30160),
            .I(\c0.n17_adj_2346_cascade_ ));
    InMux I__5768 (
            .O(N__30157),
            .I(N__30154));
    LocalMux I__5767 (
            .O(N__30154),
            .I(\c0.n30_adj_2345 ));
    CascadeMux I__5766 (
            .O(N__30151),
            .I(n31_cascade_));
    InMux I__5765 (
            .O(N__30148),
            .I(N__30145));
    LocalMux I__5764 (
            .O(N__30145),
            .I(N__30142));
    Odrv4 I__5763 (
            .O(N__30142),
            .I(\c0.n5_adj_2322 ));
    CascadeMux I__5762 (
            .O(N__30139),
            .I(\c0.n5_cascade_ ));
    CascadeMux I__5761 (
            .O(N__30136),
            .I(\c0.n17328_cascade_ ));
    InMux I__5760 (
            .O(N__30133),
            .I(N__30130));
    LocalMux I__5759 (
            .O(N__30130),
            .I(N__30126));
    InMux I__5758 (
            .O(N__30129),
            .I(N__30123));
    Span4Mux_v I__5757 (
            .O(N__30126),
            .I(N__30118));
    LocalMux I__5756 (
            .O(N__30123),
            .I(N__30118));
    Span4Mux_h I__5755 (
            .O(N__30118),
            .I(N__30114));
    InMux I__5754 (
            .O(N__30117),
            .I(N__30111));
    Span4Mux_h I__5753 (
            .O(N__30114),
            .I(N__30104));
    LocalMux I__5752 (
            .O(N__30111),
            .I(N__30104));
    InMux I__5751 (
            .O(N__30110),
            .I(N__30101));
    InMux I__5750 (
            .O(N__30109),
            .I(N__30098));
    Span4Mux_v I__5749 (
            .O(N__30104),
            .I(N__30095));
    LocalMux I__5748 (
            .O(N__30101),
            .I(\c0.FRAME_MATCHER_state_8 ));
    LocalMux I__5747 (
            .O(N__30098),
            .I(\c0.FRAME_MATCHER_state_8 ));
    Odrv4 I__5746 (
            .O(N__30095),
            .I(\c0.FRAME_MATCHER_state_8 ));
    CascadeMux I__5745 (
            .O(N__30088),
            .I(N__30085));
    InMux I__5744 (
            .O(N__30085),
            .I(N__30081));
    InMux I__5743 (
            .O(N__30084),
            .I(N__30078));
    LocalMux I__5742 (
            .O(N__30081),
            .I(N__30073));
    LocalMux I__5741 (
            .O(N__30078),
            .I(N__30073));
    Span4Mux_h I__5740 (
            .O(N__30073),
            .I(N__30070));
    Span4Mux_h I__5739 (
            .O(N__30070),
            .I(N__30067));
    Odrv4 I__5738 (
            .O(N__30067),
            .I(\c0.n16905 ));
    CascadeMux I__5737 (
            .O(N__30064),
            .I(N__30061));
    InMux I__5736 (
            .O(N__30061),
            .I(N__30058));
    LocalMux I__5735 (
            .O(N__30058),
            .I(N__30052));
    InMux I__5734 (
            .O(N__30057),
            .I(N__30049));
    InMux I__5733 (
            .O(N__30056),
            .I(N__30044));
    InMux I__5732 (
            .O(N__30055),
            .I(N__30044));
    Span4Mux_v I__5731 (
            .O(N__30052),
            .I(N__30041));
    LocalMux I__5730 (
            .O(N__30049),
            .I(\c0.FRAME_MATCHER_state_17 ));
    LocalMux I__5729 (
            .O(N__30044),
            .I(\c0.FRAME_MATCHER_state_17 ));
    Odrv4 I__5728 (
            .O(N__30041),
            .I(\c0.FRAME_MATCHER_state_17 ));
    SRMux I__5727 (
            .O(N__30034),
            .I(N__30031));
    LocalMux I__5726 (
            .O(N__30031),
            .I(\c0.n16345 ));
    InMux I__5725 (
            .O(N__30028),
            .I(N__30022));
    InMux I__5724 (
            .O(N__30027),
            .I(N__30019));
    InMux I__5723 (
            .O(N__30026),
            .I(N__30015));
    InMux I__5722 (
            .O(N__30025),
            .I(N__30012));
    LocalMux I__5721 (
            .O(N__30022),
            .I(N__30009));
    LocalMux I__5720 (
            .O(N__30019),
            .I(N__30006));
    InMux I__5719 (
            .O(N__30018),
            .I(N__30003));
    LocalMux I__5718 (
            .O(N__30015),
            .I(N__30000));
    LocalMux I__5717 (
            .O(N__30012),
            .I(N__29995));
    Span4Mux_h I__5716 (
            .O(N__30009),
            .I(N__29995));
    Span4Mux_v I__5715 (
            .O(N__30006),
            .I(N__29992));
    LocalMux I__5714 (
            .O(N__30003),
            .I(\c0.FRAME_MATCHER_state_4 ));
    Odrv12 I__5713 (
            .O(N__30000),
            .I(\c0.FRAME_MATCHER_state_4 ));
    Odrv4 I__5712 (
            .O(N__29995),
            .I(\c0.FRAME_MATCHER_state_4 ));
    Odrv4 I__5711 (
            .O(N__29992),
            .I(\c0.FRAME_MATCHER_state_4 ));
    CascadeMux I__5710 (
            .O(N__29983),
            .I(N__29978));
    CascadeMux I__5709 (
            .O(N__29982),
            .I(N__29975));
    CascadeMux I__5708 (
            .O(N__29981),
            .I(N__29969));
    InMux I__5707 (
            .O(N__29978),
            .I(N__29955));
    InMux I__5706 (
            .O(N__29975),
            .I(N__29955));
    InMux I__5705 (
            .O(N__29974),
            .I(N__29955));
    InMux I__5704 (
            .O(N__29973),
            .I(N__29955));
    InMux I__5703 (
            .O(N__29972),
            .I(N__29955));
    InMux I__5702 (
            .O(N__29969),
            .I(N__29949));
    InMux I__5701 (
            .O(N__29968),
            .I(N__29949));
    InMux I__5700 (
            .O(N__29967),
            .I(N__29946));
    InMux I__5699 (
            .O(N__29966),
            .I(N__29942));
    LocalMux I__5698 (
            .O(N__29955),
            .I(N__29938));
    InMux I__5697 (
            .O(N__29954),
            .I(N__29935));
    LocalMux I__5696 (
            .O(N__29949),
            .I(N__29930));
    LocalMux I__5695 (
            .O(N__29946),
            .I(N__29930));
    InMux I__5694 (
            .O(N__29945),
            .I(N__29927));
    LocalMux I__5693 (
            .O(N__29942),
            .I(N__29924));
    InMux I__5692 (
            .O(N__29941),
            .I(N__29921));
    Span4Mux_v I__5691 (
            .O(N__29938),
            .I(N__29912));
    LocalMux I__5690 (
            .O(N__29935),
            .I(N__29912));
    Span4Mux_v I__5689 (
            .O(N__29930),
            .I(N__29907));
    LocalMux I__5688 (
            .O(N__29927),
            .I(N__29907));
    Span4Mux_h I__5687 (
            .O(N__29924),
            .I(N__29904));
    LocalMux I__5686 (
            .O(N__29921),
            .I(N__29901));
    InMux I__5685 (
            .O(N__29920),
            .I(N__29898));
    InMux I__5684 (
            .O(N__29919),
            .I(N__29895));
    CascadeMux I__5683 (
            .O(N__29918),
            .I(N__29890));
    CascadeMux I__5682 (
            .O(N__29917),
            .I(N__29886));
    Span4Mux_h I__5681 (
            .O(N__29912),
            .I(N__29881));
    Span4Mux_v I__5680 (
            .O(N__29907),
            .I(N__29878));
    Span4Mux_v I__5679 (
            .O(N__29904),
            .I(N__29873));
    Span4Mux_h I__5678 (
            .O(N__29901),
            .I(N__29873));
    LocalMux I__5677 (
            .O(N__29898),
            .I(N__29868));
    LocalMux I__5676 (
            .O(N__29895),
            .I(N__29868));
    InMux I__5675 (
            .O(N__29894),
            .I(N__29865));
    InMux I__5674 (
            .O(N__29893),
            .I(N__29862));
    InMux I__5673 (
            .O(N__29890),
            .I(N__29851));
    InMux I__5672 (
            .O(N__29889),
            .I(N__29851));
    InMux I__5671 (
            .O(N__29886),
            .I(N__29851));
    InMux I__5670 (
            .O(N__29885),
            .I(N__29851));
    InMux I__5669 (
            .O(N__29884),
            .I(N__29851));
    Odrv4 I__5668 (
            .O(N__29881),
            .I(\c0.n4 ));
    Odrv4 I__5667 (
            .O(N__29878),
            .I(\c0.n4 ));
    Odrv4 I__5666 (
            .O(N__29873),
            .I(\c0.n4 ));
    Odrv12 I__5665 (
            .O(N__29868),
            .I(\c0.n4 ));
    LocalMux I__5664 (
            .O(N__29865),
            .I(\c0.n4 ));
    LocalMux I__5663 (
            .O(N__29862),
            .I(\c0.n4 ));
    LocalMux I__5662 (
            .O(N__29851),
            .I(\c0.n4 ));
    SRMux I__5661 (
            .O(N__29836),
            .I(N__29833));
    LocalMux I__5660 (
            .O(N__29833),
            .I(N__29830));
    Span4Mux_h I__5659 (
            .O(N__29830),
            .I(N__29827));
    Odrv4 I__5658 (
            .O(N__29827),
            .I(\c0.n16339 ));
    InMux I__5657 (
            .O(N__29824),
            .I(N__29820));
    InMux I__5656 (
            .O(N__29823),
            .I(N__29817));
    LocalMux I__5655 (
            .O(N__29820),
            .I(N__29813));
    LocalMux I__5654 (
            .O(N__29817),
            .I(N__29810));
    InMux I__5653 (
            .O(N__29816),
            .I(N__29806));
    Span4Mux_v I__5652 (
            .O(N__29813),
            .I(N__29803));
    Span4Mux_v I__5651 (
            .O(N__29810),
            .I(N__29800));
    InMux I__5650 (
            .O(N__29809),
            .I(N__29797));
    LocalMux I__5649 (
            .O(N__29806),
            .I(\c0.FRAME_MATCHER_state_14 ));
    Odrv4 I__5648 (
            .O(N__29803),
            .I(\c0.FRAME_MATCHER_state_14 ));
    Odrv4 I__5647 (
            .O(N__29800),
            .I(\c0.FRAME_MATCHER_state_14 ));
    LocalMux I__5646 (
            .O(N__29797),
            .I(\c0.FRAME_MATCHER_state_14 ));
    CascadeMux I__5645 (
            .O(N__29788),
            .I(N__29785));
    InMux I__5644 (
            .O(N__29785),
            .I(N__29782));
    LocalMux I__5643 (
            .O(N__29782),
            .I(N__29779));
    Odrv4 I__5642 (
            .O(N__29779),
            .I(\c0.n16871 ));
    InMux I__5641 (
            .O(N__29776),
            .I(N__29772));
    InMux I__5640 (
            .O(N__29775),
            .I(N__29769));
    LocalMux I__5639 (
            .O(N__29772),
            .I(N__29766));
    LocalMux I__5638 (
            .O(N__29769),
            .I(N__29763));
    Span12Mux_v I__5637 (
            .O(N__29766),
            .I(N__29760));
    Span4Mux_h I__5636 (
            .O(N__29763),
            .I(N__29757));
    Odrv12 I__5635 (
            .O(N__29760),
            .I(\c0.n16772 ));
    Odrv4 I__5634 (
            .O(N__29757),
            .I(\c0.n16772 ));
    CascadeMux I__5633 (
            .O(N__29752),
            .I(\c0.n17349_cascade_ ));
    CascadeMux I__5632 (
            .O(N__29749),
            .I(N__29746));
    InMux I__5631 (
            .O(N__29746),
            .I(N__29736));
    InMux I__5630 (
            .O(N__29745),
            .I(N__29736));
    InMux I__5629 (
            .O(N__29744),
            .I(N__29736));
    InMux I__5628 (
            .O(N__29743),
            .I(N__29729));
    LocalMux I__5627 (
            .O(N__29736),
            .I(N__29723));
    InMux I__5626 (
            .O(N__29735),
            .I(N__29716));
    InMux I__5625 (
            .O(N__29734),
            .I(N__29716));
    InMux I__5624 (
            .O(N__29733),
            .I(N__29716));
    CascadeMux I__5623 (
            .O(N__29732),
            .I(N__29713));
    LocalMux I__5622 (
            .O(N__29729),
            .I(N__29702));
    InMux I__5621 (
            .O(N__29728),
            .I(N__29695));
    InMux I__5620 (
            .O(N__29727),
            .I(N__29695));
    InMux I__5619 (
            .O(N__29726),
            .I(N__29695));
    Span4Mux_h I__5618 (
            .O(N__29723),
            .I(N__29690));
    LocalMux I__5617 (
            .O(N__29716),
            .I(N__29690));
    InMux I__5616 (
            .O(N__29713),
            .I(N__29685));
    InMux I__5615 (
            .O(N__29712),
            .I(N__29685));
    CascadeMux I__5614 (
            .O(N__29711),
            .I(N__29681));
    InMux I__5613 (
            .O(N__29710),
            .I(N__29672));
    InMux I__5612 (
            .O(N__29709),
            .I(N__29672));
    InMux I__5611 (
            .O(N__29708),
            .I(N__29672));
    CascadeMux I__5610 (
            .O(N__29707),
            .I(N__29669));
    CascadeMux I__5609 (
            .O(N__29706),
            .I(N__29666));
    CascadeMux I__5608 (
            .O(N__29705),
            .I(N__29662));
    Span4Mux_h I__5607 (
            .O(N__29702),
            .I(N__29653));
    LocalMux I__5606 (
            .O(N__29695),
            .I(N__29650));
    Span4Mux_v I__5605 (
            .O(N__29690),
            .I(N__29645));
    LocalMux I__5604 (
            .O(N__29685),
            .I(N__29642));
    InMux I__5603 (
            .O(N__29684),
            .I(N__29633));
    InMux I__5602 (
            .O(N__29681),
            .I(N__29633));
    InMux I__5601 (
            .O(N__29680),
            .I(N__29633));
    InMux I__5600 (
            .O(N__29679),
            .I(N__29633));
    LocalMux I__5599 (
            .O(N__29672),
            .I(N__29630));
    InMux I__5598 (
            .O(N__29669),
            .I(N__29619));
    InMux I__5597 (
            .O(N__29666),
            .I(N__29619));
    InMux I__5596 (
            .O(N__29665),
            .I(N__29619));
    InMux I__5595 (
            .O(N__29662),
            .I(N__29619));
    InMux I__5594 (
            .O(N__29661),
            .I(N__29619));
    InMux I__5593 (
            .O(N__29660),
            .I(N__29608));
    InMux I__5592 (
            .O(N__29659),
            .I(N__29608));
    InMux I__5591 (
            .O(N__29658),
            .I(N__29608));
    InMux I__5590 (
            .O(N__29657),
            .I(N__29608));
    InMux I__5589 (
            .O(N__29656),
            .I(N__29608));
    Span4Mux_h I__5588 (
            .O(N__29653),
            .I(N__29603));
    Span4Mux_h I__5587 (
            .O(N__29650),
            .I(N__29603));
    InMux I__5586 (
            .O(N__29649),
            .I(N__29598));
    InMux I__5585 (
            .O(N__29648),
            .I(N__29598));
    Odrv4 I__5584 (
            .O(N__29645),
            .I(\c0.n1439 ));
    Odrv12 I__5583 (
            .O(N__29642),
            .I(\c0.n1439 ));
    LocalMux I__5582 (
            .O(N__29633),
            .I(\c0.n1439 ));
    Odrv4 I__5581 (
            .O(N__29630),
            .I(\c0.n1439 ));
    LocalMux I__5580 (
            .O(N__29619),
            .I(\c0.n1439 ));
    LocalMux I__5579 (
            .O(N__29608),
            .I(\c0.n1439 ));
    Odrv4 I__5578 (
            .O(N__29603),
            .I(\c0.n1439 ));
    LocalMux I__5577 (
            .O(N__29598),
            .I(\c0.n1439 ));
    InMux I__5576 (
            .O(N__29581),
            .I(N__29578));
    LocalMux I__5575 (
            .O(N__29578),
            .I(N__29575));
    Span4Mux_h I__5574 (
            .O(N__29575),
            .I(N__29571));
    InMux I__5573 (
            .O(N__29574),
            .I(N__29568));
    Span4Mux_h I__5572 (
            .O(N__29571),
            .I(N__29565));
    LocalMux I__5571 (
            .O(N__29568),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_0 ));
    Odrv4 I__5570 (
            .O(N__29565),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_0 ));
    CascadeMux I__5569 (
            .O(N__29560),
            .I(\c0.n17590_cascade_ ));
    InMux I__5568 (
            .O(N__29557),
            .I(N__29554));
    LocalMux I__5567 (
            .O(N__29554),
            .I(n18026));
    SRMux I__5566 (
            .O(N__29551),
            .I(N__29548));
    LocalMux I__5565 (
            .O(N__29548),
            .I(N__29545));
    Span4Mux_h I__5564 (
            .O(N__29545),
            .I(N__29542));
    Span4Mux_h I__5563 (
            .O(N__29542),
            .I(N__29539));
    Odrv4 I__5562 (
            .O(N__29539),
            .I(\c0.n16347 ));
    CascadeMux I__5561 (
            .O(N__29536),
            .I(N__29533));
    InMux I__5560 (
            .O(N__29533),
            .I(N__29529));
    InMux I__5559 (
            .O(N__29532),
            .I(N__29526));
    LocalMux I__5558 (
            .O(N__29529),
            .I(N__29523));
    LocalMux I__5557 (
            .O(N__29526),
            .I(N__29520));
    Span4Mux_h I__5556 (
            .O(N__29523),
            .I(N__29517));
    Span4Mux_h I__5555 (
            .O(N__29520),
            .I(N__29514));
    Odrv4 I__5554 (
            .O(N__29517),
            .I(\c0.n16761 ));
    Odrv4 I__5553 (
            .O(N__29514),
            .I(\c0.n16761 ));
    InMux I__5552 (
            .O(N__29509),
            .I(N__29506));
    LocalMux I__5551 (
            .O(N__29506),
            .I(N__29500));
    InMux I__5550 (
            .O(N__29505),
            .I(N__29493));
    InMux I__5549 (
            .O(N__29504),
            .I(N__29493));
    InMux I__5548 (
            .O(N__29503),
            .I(N__29493));
    Span4Mux_h I__5547 (
            .O(N__29500),
            .I(N__29490));
    LocalMux I__5546 (
            .O(N__29493),
            .I(\c0.FRAME_MATCHER_state_28 ));
    Odrv4 I__5545 (
            .O(N__29490),
            .I(\c0.FRAME_MATCHER_state_28 ));
    SRMux I__5544 (
            .O(N__29485),
            .I(N__29482));
    LocalMux I__5543 (
            .O(N__29482),
            .I(N__29479));
    Odrv4 I__5542 (
            .O(N__29479),
            .I(\c0.n16353 ));
    CascadeMux I__5541 (
            .O(N__29476),
            .I(N__29469));
    InMux I__5540 (
            .O(N__29475),
            .I(N__29466));
    InMux I__5539 (
            .O(N__29474),
            .I(N__29463));
    InMux I__5538 (
            .O(N__29473),
            .I(N__29460));
    InMux I__5537 (
            .O(N__29472),
            .I(N__29455));
    InMux I__5536 (
            .O(N__29469),
            .I(N__29455));
    LocalMux I__5535 (
            .O(N__29466),
            .I(N__29452));
    LocalMux I__5534 (
            .O(N__29463),
            .I(N__29449));
    LocalMux I__5533 (
            .O(N__29460),
            .I(N__29444));
    LocalMux I__5532 (
            .O(N__29455),
            .I(N__29444));
    Span4Mux_h I__5531 (
            .O(N__29452),
            .I(N__29439));
    Span4Mux_h I__5530 (
            .O(N__29449),
            .I(N__29439));
    Odrv4 I__5529 (
            .O(N__29444),
            .I(\c0.FRAME_MATCHER_state_24 ));
    Odrv4 I__5528 (
            .O(N__29439),
            .I(\c0.FRAME_MATCHER_state_24 ));
    SRMux I__5527 (
            .O(N__29434),
            .I(N__29431));
    LocalMux I__5526 (
            .O(N__29431),
            .I(\c0.n16361 ));
    InMux I__5525 (
            .O(N__29428),
            .I(N__29422));
    InMux I__5524 (
            .O(N__29427),
            .I(N__29422));
    LocalMux I__5523 (
            .O(N__29422),
            .I(r_Tx_Data_0));
    InMux I__5522 (
            .O(N__29419),
            .I(N__29416));
    LocalMux I__5521 (
            .O(N__29416),
            .I(N__29413));
    Span4Mux_h I__5520 (
            .O(N__29413),
            .I(N__29410));
    Odrv4 I__5519 (
            .O(N__29410),
            .I(n17394));
    InMux I__5518 (
            .O(N__29407),
            .I(N__29404));
    LocalMux I__5517 (
            .O(N__29404),
            .I(N__29401));
    Odrv4 I__5516 (
            .O(N__29401),
            .I(\c0.n8_adj_2160 ));
    CascadeMux I__5515 (
            .O(N__29398),
            .I(\c0.n15_cascade_ ));
    CascadeMux I__5514 (
            .O(N__29395),
            .I(\c0.n12_adj_2150_cascade_ ));
    InMux I__5513 (
            .O(N__29392),
            .I(N__29388));
    InMux I__5512 (
            .O(N__29391),
            .I(N__29385));
    LocalMux I__5511 (
            .O(N__29388),
            .I(r_Tx_Data_2));
    LocalMux I__5510 (
            .O(N__29385),
            .I(r_Tx_Data_2));
    CascadeMux I__5509 (
            .O(N__29380),
            .I(N__29377));
    InMux I__5508 (
            .O(N__29377),
            .I(N__29374));
    LocalMux I__5507 (
            .O(N__29374),
            .I(n10_adj_2426));
    CascadeMux I__5506 (
            .O(N__29371),
            .I(n10_adj_2407_cascade_));
    InMux I__5505 (
            .O(N__29368),
            .I(N__29365));
    LocalMux I__5504 (
            .O(N__29365),
            .I(N__29362));
    Span4Mux_h I__5503 (
            .O(N__29362),
            .I(N__29358));
    InMux I__5502 (
            .O(N__29361),
            .I(N__29355));
    Span4Mux_h I__5501 (
            .O(N__29358),
            .I(N__29352));
    LocalMux I__5500 (
            .O(N__29355),
            .I(r_Tx_Data_4));
    Odrv4 I__5499 (
            .O(N__29352),
            .I(r_Tx_Data_4));
    CascadeMux I__5498 (
            .O(N__29347),
            .I(\c0.tx2.o_Tx_Serial_N_2064_cascade_ ));
    CascadeMux I__5497 (
            .O(N__29344),
            .I(N__29337));
    CascadeMux I__5496 (
            .O(N__29343),
            .I(N__29334));
    InMux I__5495 (
            .O(N__29342),
            .I(N__29331));
    InMux I__5494 (
            .O(N__29341),
            .I(N__29328));
    InMux I__5493 (
            .O(N__29340),
            .I(N__29322));
    InMux I__5492 (
            .O(N__29337),
            .I(N__29315));
    InMux I__5491 (
            .O(N__29334),
            .I(N__29315));
    LocalMux I__5490 (
            .O(N__29331),
            .I(N__29310));
    LocalMux I__5489 (
            .O(N__29328),
            .I(N__29310));
    InMux I__5488 (
            .O(N__29327),
            .I(N__29307));
    InMux I__5487 (
            .O(N__29326),
            .I(N__29302));
    InMux I__5486 (
            .O(N__29325),
            .I(N__29302));
    LocalMux I__5485 (
            .O(N__29322),
            .I(N__29299));
    InMux I__5484 (
            .O(N__29321),
            .I(N__29296));
    InMux I__5483 (
            .O(N__29320),
            .I(N__29293));
    LocalMux I__5482 (
            .O(N__29315),
            .I(N__29288));
    Span4Mux_h I__5481 (
            .O(N__29310),
            .I(N__29288));
    LocalMux I__5480 (
            .O(N__29307),
            .I(r_SM_Main_0_adj_2445));
    LocalMux I__5479 (
            .O(N__29302),
            .I(r_SM_Main_0_adj_2445));
    Odrv12 I__5478 (
            .O(N__29299),
            .I(r_SM_Main_0_adj_2445));
    LocalMux I__5477 (
            .O(N__29296),
            .I(r_SM_Main_0_adj_2445));
    LocalMux I__5476 (
            .O(N__29293),
            .I(r_SM_Main_0_adj_2445));
    Odrv4 I__5475 (
            .O(N__29288),
            .I(r_SM_Main_0_adj_2445));
    InMux I__5474 (
            .O(N__29275),
            .I(N__29272));
    LocalMux I__5473 (
            .O(N__29272),
            .I(N__29269));
    Odrv4 I__5472 (
            .O(N__29269),
            .I(n3));
    CascadeMux I__5471 (
            .O(N__29266),
            .I(N__29263));
    InMux I__5470 (
            .O(N__29263),
            .I(N__29260));
    LocalMux I__5469 (
            .O(N__29260),
            .I(n5029));
    CascadeMux I__5468 (
            .O(N__29257),
            .I(N__29252));
    InMux I__5467 (
            .O(N__29256),
            .I(N__29249));
    InMux I__5466 (
            .O(N__29255),
            .I(N__29244));
    InMux I__5465 (
            .O(N__29252),
            .I(N__29244));
    LocalMux I__5464 (
            .O(N__29249),
            .I(r_Bit_Index_2_adj_2455));
    LocalMux I__5463 (
            .O(N__29244),
            .I(r_Bit_Index_2_adj_2455));
    CascadeMux I__5462 (
            .O(N__29239),
            .I(N__29236));
    InMux I__5461 (
            .O(N__29236),
            .I(N__29233));
    LocalMux I__5460 (
            .O(N__29233),
            .I(N__29229));
    InMux I__5459 (
            .O(N__29232),
            .I(N__29226));
    Odrv12 I__5458 (
            .O(N__29229),
            .I(\c0.tx2.n13281 ));
    LocalMux I__5457 (
            .O(N__29226),
            .I(\c0.tx2.n13281 ));
    CascadeMux I__5456 (
            .O(N__29221),
            .I(\c0.n2_adj_2266_cascade_ ));
    CascadeMux I__5455 (
            .O(N__29218),
            .I(\c0.n18098_cascade_ ));
    CascadeMux I__5454 (
            .O(N__29215),
            .I(\c0.n10_adj_2139_cascade_ ));
    InMux I__5453 (
            .O(N__29212),
            .I(N__29209));
    LocalMux I__5452 (
            .O(N__29209),
            .I(N__29206));
    Span4Mux_h I__5451 (
            .O(N__29206),
            .I(N__29203));
    IoSpan4Mux I__5450 (
            .O(N__29203),
            .I(N__29200));
    Odrv4 I__5449 (
            .O(N__29200),
            .I(\c0.rx.r_Rx_Data_R ));
    CascadeMux I__5448 (
            .O(N__29197),
            .I(\c0.tx2.n18113_cascade_ ));
    InMux I__5447 (
            .O(N__29194),
            .I(N__29188));
    InMux I__5446 (
            .O(N__29193),
            .I(N__29188));
    LocalMux I__5445 (
            .O(N__29188),
            .I(n10398));
    InMux I__5444 (
            .O(N__29185),
            .I(N__29177));
    InMux I__5443 (
            .O(N__29184),
            .I(N__29177));
    InMux I__5442 (
            .O(N__29183),
            .I(N__29172));
    InMux I__5441 (
            .O(N__29182),
            .I(N__29172));
    LocalMux I__5440 (
            .O(N__29177),
            .I(N__29169));
    LocalMux I__5439 (
            .O(N__29172),
            .I(N__29166));
    Span12Mux_h I__5438 (
            .O(N__29169),
            .I(N__29163));
    Span4Mux_h I__5437 (
            .O(N__29166),
            .I(N__29160));
    Odrv12 I__5436 (
            .O(N__29163),
            .I(n17194));
    Odrv4 I__5435 (
            .O(N__29160),
            .I(n17194));
    CascadeMux I__5434 (
            .O(N__29155),
            .I(n10398_cascade_));
    InMux I__5433 (
            .O(N__29152),
            .I(N__29149));
    LocalMux I__5432 (
            .O(N__29149),
            .I(\c0.tx2.n17906 ));
    InMux I__5431 (
            .O(N__29146),
            .I(N__29143));
    LocalMux I__5430 (
            .O(N__29143),
            .I(N__29140));
    Odrv4 I__5429 (
            .O(N__29140),
            .I(\c0.tx2.n18116 ));
    InMux I__5428 (
            .O(N__29137),
            .I(N__29134));
    LocalMux I__5427 (
            .O(N__29134),
            .I(N__29129));
    InMux I__5426 (
            .O(N__29133),
            .I(N__29126));
    InMux I__5425 (
            .O(N__29132),
            .I(N__29123));
    Span4Mux_v I__5424 (
            .O(N__29129),
            .I(N__29116));
    LocalMux I__5423 (
            .O(N__29126),
            .I(N__29116));
    LocalMux I__5422 (
            .O(N__29123),
            .I(N__29116));
    Span4Mux_h I__5421 (
            .O(N__29116),
            .I(N__29111));
    InMux I__5420 (
            .O(N__29115),
            .I(N__29106));
    InMux I__5419 (
            .O(N__29114),
            .I(N__29106));
    Odrv4 I__5418 (
            .O(N__29111),
            .I(\c0.data_in_frame_1_1 ));
    LocalMux I__5417 (
            .O(N__29106),
            .I(\c0.data_in_frame_1_1 ));
    InMux I__5416 (
            .O(N__29101),
            .I(N__29098));
    LocalMux I__5415 (
            .O(N__29098),
            .I(N__29095));
    Span4Mux_v I__5414 (
            .O(N__29095),
            .I(N__29092));
    Odrv4 I__5413 (
            .O(N__29092),
            .I(\c0.n17014 ));
    CascadeMux I__5412 (
            .O(N__29089),
            .I(\c0.n23_adj_2156_cascade_ ));
    InMux I__5411 (
            .O(N__29086),
            .I(N__29082));
    InMux I__5410 (
            .O(N__29085),
            .I(N__29079));
    LocalMux I__5409 (
            .O(N__29082),
            .I(N__29076));
    LocalMux I__5408 (
            .O(N__29079),
            .I(N__29073));
    Span4Mux_h I__5407 (
            .O(N__29076),
            .I(N__29070));
    Span4Mux_h I__5406 (
            .O(N__29073),
            .I(N__29067));
    Odrv4 I__5405 (
            .O(N__29070),
            .I(\c0.n17001 ));
    Odrv4 I__5404 (
            .O(N__29067),
            .I(\c0.n17001 ));
    InMux I__5403 (
            .O(N__29062),
            .I(N__29059));
    LocalMux I__5402 (
            .O(N__29059),
            .I(\c0.n28_adj_2183 ));
    InMux I__5401 (
            .O(N__29056),
            .I(N__29052));
    InMux I__5400 (
            .O(N__29055),
            .I(N__29046));
    LocalMux I__5399 (
            .O(N__29052),
            .I(N__29042));
    InMux I__5398 (
            .O(N__29051),
            .I(N__29037));
    InMux I__5397 (
            .O(N__29050),
            .I(N__29037));
    InMux I__5396 (
            .O(N__29049),
            .I(N__29033));
    LocalMux I__5395 (
            .O(N__29046),
            .I(N__29030));
    InMux I__5394 (
            .O(N__29045),
            .I(N__29027));
    Span4Mux_h I__5393 (
            .O(N__29042),
            .I(N__29022));
    LocalMux I__5392 (
            .O(N__29037),
            .I(N__29022));
    InMux I__5391 (
            .O(N__29036),
            .I(N__29019));
    LocalMux I__5390 (
            .O(N__29033),
            .I(N__29014));
    Span4Mux_h I__5389 (
            .O(N__29030),
            .I(N__29014));
    LocalMux I__5388 (
            .O(N__29027),
            .I(data_in_frame_0_6));
    Odrv4 I__5387 (
            .O(N__29022),
            .I(data_in_frame_0_6));
    LocalMux I__5386 (
            .O(N__29019),
            .I(data_in_frame_0_6));
    Odrv4 I__5385 (
            .O(N__29014),
            .I(data_in_frame_0_6));
    InMux I__5384 (
            .O(N__29005),
            .I(N__29002));
    LocalMux I__5383 (
            .O(N__29002),
            .I(N__28999));
    Odrv4 I__5382 (
            .O(N__28999),
            .I(\c0.n2340 ));
    CascadeMux I__5381 (
            .O(N__28996),
            .I(N__28993));
    InMux I__5380 (
            .O(N__28993),
            .I(N__28989));
    InMux I__5379 (
            .O(N__28992),
            .I(N__28986));
    LocalMux I__5378 (
            .O(N__28989),
            .I(N__28983));
    LocalMux I__5377 (
            .O(N__28986),
            .I(\c0.data_in_frame_9_0 ));
    Odrv12 I__5376 (
            .O(N__28983),
            .I(\c0.data_in_frame_9_0 ));
    InMux I__5375 (
            .O(N__28978),
            .I(N__28974));
    InMux I__5374 (
            .O(N__28977),
            .I(N__28971));
    LocalMux I__5373 (
            .O(N__28974),
            .I(N__28968));
    LocalMux I__5372 (
            .O(N__28971),
            .I(N__28965));
    Odrv12 I__5371 (
            .O(N__28968),
            .I(\c0.n17004 ));
    Odrv4 I__5370 (
            .O(N__28965),
            .I(\c0.n17004 ));
    InMux I__5369 (
            .O(N__28960),
            .I(N__28957));
    LocalMux I__5368 (
            .O(N__28957),
            .I(\c0.n19 ));
    InMux I__5367 (
            .O(N__28954),
            .I(N__28950));
    InMux I__5366 (
            .O(N__28953),
            .I(N__28947));
    LocalMux I__5365 (
            .O(N__28950),
            .I(N__28944));
    LocalMux I__5364 (
            .O(N__28947),
            .I(data_in_frame_7_3));
    Odrv12 I__5363 (
            .O(N__28944),
            .I(data_in_frame_7_3));
    InMux I__5362 (
            .O(N__28939),
            .I(N__28935));
    InMux I__5361 (
            .O(N__28938),
            .I(N__28932));
    LocalMux I__5360 (
            .O(N__28935),
            .I(N__28929));
    LocalMux I__5359 (
            .O(N__28932),
            .I(N__28926));
    Span4Mux_v I__5358 (
            .O(N__28929),
            .I(N__28923));
    Odrv4 I__5357 (
            .O(N__28926),
            .I(\c0.n2336 ));
    Odrv4 I__5356 (
            .O(N__28923),
            .I(\c0.n2336 ));
    CascadeMux I__5355 (
            .O(N__28918),
            .I(N__28915));
    InMux I__5354 (
            .O(N__28915),
            .I(N__28912));
    LocalMux I__5353 (
            .O(N__28912),
            .I(N__28909));
    Span4Mux_h I__5352 (
            .O(N__28909),
            .I(N__28905));
    InMux I__5351 (
            .O(N__28908),
            .I(N__28902));
    Span4Mux_h I__5350 (
            .O(N__28905),
            .I(N__28899));
    LocalMux I__5349 (
            .O(N__28902),
            .I(data_in_frame_7_5));
    Odrv4 I__5348 (
            .O(N__28899),
            .I(data_in_frame_7_5));
    InMux I__5347 (
            .O(N__28894),
            .I(N__28891));
    LocalMux I__5346 (
            .O(N__28891),
            .I(N__28888));
    Span4Mux_h I__5345 (
            .O(N__28888),
            .I(N__28884));
    InMux I__5344 (
            .O(N__28887),
            .I(N__28881));
    Odrv4 I__5343 (
            .O(N__28884),
            .I(\c0.n9541 ));
    LocalMux I__5342 (
            .O(N__28881),
            .I(\c0.n9541 ));
    InMux I__5341 (
            .O(N__28876),
            .I(N__28873));
    LocalMux I__5340 (
            .O(N__28873),
            .I(N__28869));
    InMux I__5339 (
            .O(N__28872),
            .I(N__28866));
    Span4Mux_h I__5338 (
            .O(N__28869),
            .I(N__28863));
    LocalMux I__5337 (
            .O(N__28866),
            .I(data_in_frame_6_0));
    Odrv4 I__5336 (
            .O(N__28863),
            .I(data_in_frame_6_0));
    InMux I__5335 (
            .O(N__28858),
            .I(N__28855));
    LocalMux I__5334 (
            .O(N__28855),
            .I(N__28852));
    Span4Mux_h I__5333 (
            .O(N__28852),
            .I(N__28848));
    InMux I__5332 (
            .O(N__28851),
            .I(N__28845));
    Span4Mux_h I__5331 (
            .O(N__28848),
            .I(N__28842));
    LocalMux I__5330 (
            .O(N__28845),
            .I(data_in_frame_6_5));
    Odrv4 I__5329 (
            .O(N__28842),
            .I(data_in_frame_6_5));
    CascadeMux I__5328 (
            .O(N__28837),
            .I(\c0.n20_cascade_ ));
    InMux I__5327 (
            .O(N__28834),
            .I(N__28828));
    InMux I__5326 (
            .O(N__28833),
            .I(N__28828));
    LocalMux I__5325 (
            .O(N__28828),
            .I(N__28824));
    InMux I__5324 (
            .O(N__28827),
            .I(N__28821));
    Odrv4 I__5323 (
            .O(N__28824),
            .I(\c0.n2342 ));
    LocalMux I__5322 (
            .O(N__28821),
            .I(\c0.n2342 ));
    InMux I__5321 (
            .O(N__28816),
            .I(N__28812));
    InMux I__5320 (
            .O(N__28815),
            .I(N__28809));
    LocalMux I__5319 (
            .O(N__28812),
            .I(\c0.data_in_frame_9_1 ));
    LocalMux I__5318 (
            .O(N__28809),
            .I(\c0.data_in_frame_9_1 ));
    CascadeMux I__5317 (
            .O(N__28804),
            .I(N__28792));
    InMux I__5316 (
            .O(N__28803),
            .I(N__28789));
    InMux I__5315 (
            .O(N__28802),
            .I(N__28786));
    InMux I__5314 (
            .O(N__28801),
            .I(N__28782));
    InMux I__5313 (
            .O(N__28800),
            .I(N__28779));
    InMux I__5312 (
            .O(N__28799),
            .I(N__28770));
    InMux I__5311 (
            .O(N__28798),
            .I(N__28770));
    InMux I__5310 (
            .O(N__28797),
            .I(N__28770));
    InMux I__5309 (
            .O(N__28796),
            .I(N__28770));
    InMux I__5308 (
            .O(N__28795),
            .I(N__28765));
    InMux I__5307 (
            .O(N__28792),
            .I(N__28765));
    LocalMux I__5306 (
            .O(N__28789),
            .I(N__28755));
    LocalMux I__5305 (
            .O(N__28786),
            .I(N__28755));
    InMux I__5304 (
            .O(N__28785),
            .I(N__28752));
    LocalMux I__5303 (
            .O(N__28782),
            .I(N__28747));
    LocalMux I__5302 (
            .O(N__28779),
            .I(N__28747));
    LocalMux I__5301 (
            .O(N__28770),
            .I(N__28742));
    LocalMux I__5300 (
            .O(N__28765),
            .I(N__28742));
    InMux I__5299 (
            .O(N__28764),
            .I(N__28739));
    InMux I__5298 (
            .O(N__28763),
            .I(N__28736));
    InMux I__5297 (
            .O(N__28762),
            .I(N__28729));
    InMux I__5296 (
            .O(N__28761),
            .I(N__28729));
    InMux I__5295 (
            .O(N__28760),
            .I(N__28729));
    Span4Mux_v I__5294 (
            .O(N__28755),
            .I(N__28726));
    LocalMux I__5293 (
            .O(N__28752),
            .I(N__28723));
    Span4Mux_v I__5292 (
            .O(N__28747),
            .I(N__28718));
    Span4Mux_h I__5291 (
            .O(N__28742),
            .I(N__28718));
    LocalMux I__5290 (
            .O(N__28739),
            .I(\c0.n8_adj_2310 ));
    LocalMux I__5289 (
            .O(N__28736),
            .I(\c0.n8_adj_2310 ));
    LocalMux I__5288 (
            .O(N__28729),
            .I(\c0.n8_adj_2310 ));
    Odrv4 I__5287 (
            .O(N__28726),
            .I(\c0.n8_adj_2310 ));
    Odrv12 I__5286 (
            .O(N__28723),
            .I(\c0.n8_adj_2310 ));
    Odrv4 I__5285 (
            .O(N__28718),
            .I(\c0.n8_adj_2310 ));
    InMux I__5284 (
            .O(N__28705),
            .I(N__28699));
    InMux I__5283 (
            .O(N__28704),
            .I(N__28699));
    LocalMux I__5282 (
            .O(N__28699),
            .I(\c0.data_in_frame_9_5 ));
    IoInMux I__5281 (
            .O(N__28696),
            .I(N__28693));
    LocalMux I__5280 (
            .O(N__28693),
            .I(N__28690));
    IoSpan4Mux I__5279 (
            .O(N__28690),
            .I(N__28686));
    InMux I__5278 (
            .O(N__28689),
            .I(N__28683));
    Sp12to4 I__5277 (
            .O(N__28686),
            .I(N__28678));
    LocalMux I__5276 (
            .O(N__28683),
            .I(N__28678));
    Span12Mux_s6_h I__5275 (
            .O(N__28678),
            .I(N__28674));
    InMux I__5274 (
            .O(N__28677),
            .I(N__28671));
    Odrv12 I__5273 (
            .O(N__28674),
            .I(tx2_o));
    LocalMux I__5272 (
            .O(N__28671),
            .I(tx2_o));
    SRMux I__5271 (
            .O(N__28666),
            .I(N__28663));
    LocalMux I__5270 (
            .O(N__28663),
            .I(N__28660));
    Span4Mux_h I__5269 (
            .O(N__28660),
            .I(N__28657));
    Odrv4 I__5268 (
            .O(N__28657),
            .I(\c0.n3_adj_2240 ));
    InMux I__5267 (
            .O(N__28654),
            .I(N__28651));
    LocalMux I__5266 (
            .O(N__28651),
            .I(N__28646));
    InMux I__5265 (
            .O(N__28650),
            .I(N__28638));
    InMux I__5264 (
            .O(N__28649),
            .I(N__28638));
    Span4Mux_h I__5263 (
            .O(N__28646),
            .I(N__28635));
    InMux I__5262 (
            .O(N__28645),
            .I(N__28632));
    InMux I__5261 (
            .O(N__28644),
            .I(N__28627));
    InMux I__5260 (
            .O(N__28643),
            .I(N__28627));
    LocalMux I__5259 (
            .O(N__28638),
            .I(N__28624));
    Odrv4 I__5258 (
            .O(N__28635),
            .I(data_in_frame_0_7));
    LocalMux I__5257 (
            .O(N__28632),
            .I(data_in_frame_0_7));
    LocalMux I__5256 (
            .O(N__28627),
            .I(data_in_frame_0_7));
    Odrv4 I__5255 (
            .O(N__28624),
            .I(data_in_frame_0_7));
    CascadeMux I__5254 (
            .O(N__28615),
            .I(N__28612));
    InMux I__5253 (
            .O(N__28612),
            .I(N__28607));
    CascadeMux I__5252 (
            .O(N__28611),
            .I(N__28604));
    InMux I__5251 (
            .O(N__28610),
            .I(N__28600));
    LocalMux I__5250 (
            .O(N__28607),
            .I(N__28597));
    InMux I__5249 (
            .O(N__28604),
            .I(N__28594));
    InMux I__5248 (
            .O(N__28603),
            .I(N__28591));
    LocalMux I__5247 (
            .O(N__28600),
            .I(N__28586));
    Span4Mux_v I__5246 (
            .O(N__28597),
            .I(N__28586));
    LocalMux I__5245 (
            .O(N__28594),
            .I(\c0.data_in_frame_1_7 ));
    LocalMux I__5244 (
            .O(N__28591),
            .I(\c0.data_in_frame_1_7 ));
    Odrv4 I__5243 (
            .O(N__28586),
            .I(\c0.data_in_frame_1_7 ));
    InMux I__5242 (
            .O(N__28579),
            .I(N__28576));
    LocalMux I__5241 (
            .O(N__28576),
            .I(N__28572));
    InMux I__5240 (
            .O(N__28575),
            .I(N__28569));
    Span4Mux_v I__5239 (
            .O(N__28572),
            .I(N__28565));
    LocalMux I__5238 (
            .O(N__28569),
            .I(N__28562));
    InMux I__5237 (
            .O(N__28568),
            .I(N__28558));
    Span4Mux_h I__5236 (
            .O(N__28565),
            .I(N__28555));
    Span4Mux_h I__5235 (
            .O(N__28562),
            .I(N__28552));
    InMux I__5234 (
            .O(N__28561),
            .I(N__28549));
    LocalMux I__5233 (
            .O(N__28558),
            .I(\c0.data_in_frame_1_4 ));
    Odrv4 I__5232 (
            .O(N__28555),
            .I(\c0.data_in_frame_1_4 ));
    Odrv4 I__5231 (
            .O(N__28552),
            .I(\c0.data_in_frame_1_4 ));
    LocalMux I__5230 (
            .O(N__28549),
            .I(\c0.data_in_frame_1_4 ));
    InMux I__5229 (
            .O(N__28540),
            .I(N__28537));
    LocalMux I__5228 (
            .O(N__28537),
            .I(N__28534));
    Span4Mux_v I__5227 (
            .O(N__28534),
            .I(N__28531));
    Odrv4 I__5226 (
            .O(N__28531),
            .I(\c0.n27_adj_2342 ));
    CascadeMux I__5225 (
            .O(N__28528),
            .I(\c0.n23_adj_2341_cascade_ ));
    InMux I__5224 (
            .O(N__28525),
            .I(N__28521));
    CascadeMux I__5223 (
            .O(N__28524),
            .I(N__28518));
    LocalMux I__5222 (
            .O(N__28521),
            .I(N__28515));
    InMux I__5221 (
            .O(N__28518),
            .I(N__28510));
    Span4Mux_h I__5220 (
            .O(N__28515),
            .I(N__28507));
    InMux I__5219 (
            .O(N__28514),
            .I(N__28502));
    InMux I__5218 (
            .O(N__28513),
            .I(N__28502));
    LocalMux I__5217 (
            .O(N__28510),
            .I(\c0.data_in_frame_1_3 ));
    Odrv4 I__5216 (
            .O(N__28507),
            .I(\c0.data_in_frame_1_3 ));
    LocalMux I__5215 (
            .O(N__28502),
            .I(\c0.data_in_frame_1_3 ));
    InMux I__5214 (
            .O(N__28495),
            .I(N__28492));
    LocalMux I__5213 (
            .O(N__28492),
            .I(N__28489));
    Odrv12 I__5212 (
            .O(N__28489),
            .I(\c0.n21_adj_2171 ));
    CascadeMux I__5211 (
            .O(N__28486),
            .I(N__28483));
    InMux I__5210 (
            .O(N__28483),
            .I(N__28480));
    LocalMux I__5209 (
            .O(N__28480),
            .I(N__28477));
    Span4Mux_h I__5208 (
            .O(N__28477),
            .I(N__28474));
    Odrv4 I__5207 (
            .O(N__28474),
            .I(\c0.n15930 ));
    InMux I__5206 (
            .O(N__28471),
            .I(N__28468));
    LocalMux I__5205 (
            .O(N__28468),
            .I(N__28464));
    InMux I__5204 (
            .O(N__28467),
            .I(N__28461));
    Span4Mux_h I__5203 (
            .O(N__28464),
            .I(N__28458));
    LocalMux I__5202 (
            .O(N__28461),
            .I(\c0.data_in_frame_10_7 ));
    Odrv4 I__5201 (
            .O(N__28458),
            .I(\c0.data_in_frame_10_7 ));
    CascadeMux I__5200 (
            .O(N__28453),
            .I(\c0.n17352_cascade_ ));
    CascadeMux I__5199 (
            .O(N__28450),
            .I(N__28447));
    InMux I__5198 (
            .O(N__28447),
            .I(N__28444));
    LocalMux I__5197 (
            .O(N__28444),
            .I(\c0.n27_adj_2196 ));
    InMux I__5196 (
            .O(N__28441),
            .I(N__28438));
    LocalMux I__5195 (
            .O(N__28438),
            .I(N__28435));
    Odrv12 I__5194 (
            .O(N__28435),
            .I(\c0.n25 ));
    CascadeMux I__5193 (
            .O(N__28432),
            .I(\c0.n15846_cascade_ ));
    InMux I__5192 (
            .O(N__28429),
            .I(N__28426));
    LocalMux I__5191 (
            .O(N__28426),
            .I(N__28423));
    Odrv4 I__5190 (
            .O(N__28423),
            .I(\c0.n15929 ));
    InMux I__5189 (
            .O(N__28420),
            .I(N__28417));
    LocalMux I__5188 (
            .O(N__28417),
            .I(\c0.n26_adj_2184 ));
    InMux I__5187 (
            .O(N__28414),
            .I(N__28411));
    LocalMux I__5186 (
            .O(N__28411),
            .I(N__28408));
    Span4Mux_h I__5185 (
            .O(N__28408),
            .I(N__28405));
    Odrv4 I__5184 (
            .O(N__28405),
            .I(\c0.n15938 ));
    InMux I__5183 (
            .O(N__28402),
            .I(N__28399));
    LocalMux I__5182 (
            .O(N__28399),
            .I(N__28394));
    InMux I__5181 (
            .O(N__28398),
            .I(N__28389));
    InMux I__5180 (
            .O(N__28397),
            .I(N__28386));
    Span4Mux_v I__5179 (
            .O(N__28394),
            .I(N__28383));
    InMux I__5178 (
            .O(N__28393),
            .I(N__28380));
    InMux I__5177 (
            .O(N__28392),
            .I(N__28377));
    LocalMux I__5176 (
            .O(N__28389),
            .I(N__28374));
    LocalMux I__5175 (
            .O(N__28386),
            .I(\c0.data_in_frame_1_2 ));
    Odrv4 I__5174 (
            .O(N__28383),
            .I(\c0.data_in_frame_1_2 ));
    LocalMux I__5173 (
            .O(N__28380),
            .I(\c0.data_in_frame_1_2 ));
    LocalMux I__5172 (
            .O(N__28377),
            .I(\c0.data_in_frame_1_2 ));
    Odrv4 I__5171 (
            .O(N__28374),
            .I(\c0.data_in_frame_1_2 ));
    CascadeMux I__5170 (
            .O(N__28363),
            .I(N__28360));
    InMux I__5169 (
            .O(N__28360),
            .I(N__28357));
    LocalMux I__5168 (
            .O(N__28357),
            .I(N__28353));
    InMux I__5167 (
            .O(N__28356),
            .I(N__28350));
    Span4Mux_v I__5166 (
            .O(N__28353),
            .I(N__28347));
    LocalMux I__5165 (
            .O(N__28350),
            .I(\c0.data_in_frame_9_3 ));
    Odrv4 I__5164 (
            .O(N__28347),
            .I(\c0.data_in_frame_9_3 ));
    CascadeMux I__5163 (
            .O(N__28342),
            .I(N__28339));
    InMux I__5162 (
            .O(N__28339),
            .I(N__28336));
    LocalMux I__5161 (
            .O(N__28336),
            .I(N__28333));
    Span4Mux_v I__5160 (
            .O(N__28333),
            .I(N__28330));
    Span4Mux_h I__5159 (
            .O(N__28330),
            .I(N__28327));
    Odrv4 I__5158 (
            .O(N__28327),
            .I(\c0.n8603 ));
    CascadeMux I__5157 (
            .O(N__28324),
            .I(N__28318));
    CascadeMux I__5156 (
            .O(N__28323),
            .I(N__28315));
    CascadeMux I__5155 (
            .O(N__28322),
            .I(N__28312));
    InMux I__5154 (
            .O(N__28321),
            .I(N__28309));
    InMux I__5153 (
            .O(N__28318),
            .I(N__28304));
    InMux I__5152 (
            .O(N__28315),
            .I(N__28304));
    InMux I__5151 (
            .O(N__28312),
            .I(N__28301));
    LocalMux I__5150 (
            .O(N__28309),
            .I(N__28298));
    LocalMux I__5149 (
            .O(N__28304),
            .I(\c0.FRAME_MATCHER_i_11 ));
    LocalMux I__5148 (
            .O(N__28301),
            .I(\c0.FRAME_MATCHER_i_11 ));
    Odrv12 I__5147 (
            .O(N__28298),
            .I(\c0.FRAME_MATCHER_i_11 ));
    InMux I__5146 (
            .O(N__28291),
            .I(N__28287));
    CascadeMux I__5145 (
            .O(N__28290),
            .I(N__28284));
    LocalMux I__5144 (
            .O(N__28287),
            .I(N__28279));
    InMux I__5143 (
            .O(N__28284),
            .I(N__28274));
    InMux I__5142 (
            .O(N__28283),
            .I(N__28274));
    InMux I__5141 (
            .O(N__28282),
            .I(N__28271));
    Span4Mux_v I__5140 (
            .O(N__28279),
            .I(N__28268));
    LocalMux I__5139 (
            .O(N__28274),
            .I(N__28261));
    LocalMux I__5138 (
            .O(N__28271),
            .I(N__28261));
    Span4Mux_h I__5137 (
            .O(N__28268),
            .I(N__28261));
    Odrv4 I__5136 (
            .O(N__28261),
            .I(\c0.FRAME_MATCHER_i_14 ));
    CascadeMux I__5135 (
            .O(N__28258),
            .I(N__28255));
    InMux I__5134 (
            .O(N__28255),
            .I(N__28251));
    CascadeMux I__5133 (
            .O(N__28254),
            .I(N__28246));
    LocalMux I__5132 (
            .O(N__28251),
            .I(N__28243));
    CascadeMux I__5131 (
            .O(N__28250),
            .I(N__28240));
    CascadeMux I__5130 (
            .O(N__28249),
            .I(N__28237));
    InMux I__5129 (
            .O(N__28246),
            .I(N__28234));
    Span4Mux_v I__5128 (
            .O(N__28243),
            .I(N__28231));
    InMux I__5127 (
            .O(N__28240),
            .I(N__28226));
    InMux I__5126 (
            .O(N__28237),
            .I(N__28226));
    LocalMux I__5125 (
            .O(N__28234),
            .I(N__28223));
    Span4Mux_h I__5124 (
            .O(N__28231),
            .I(N__28220));
    LocalMux I__5123 (
            .O(N__28226),
            .I(\c0.FRAME_MATCHER_i_15 ));
    Odrv4 I__5122 (
            .O(N__28223),
            .I(\c0.FRAME_MATCHER_i_15 ));
    Odrv4 I__5121 (
            .O(N__28220),
            .I(\c0.FRAME_MATCHER_i_15 ));
    InMux I__5120 (
            .O(N__28213),
            .I(N__28210));
    LocalMux I__5119 (
            .O(N__28210),
            .I(N__28207));
    Odrv4 I__5118 (
            .O(N__28207),
            .I(\c0.n48 ));
    InMux I__5117 (
            .O(N__28204),
            .I(N__28201));
    LocalMux I__5116 (
            .O(N__28201),
            .I(N__28198));
    Span4Mux_h I__5115 (
            .O(N__28198),
            .I(N__28195));
    Span4Mux_h I__5114 (
            .O(N__28195),
            .I(N__28192));
    Odrv4 I__5113 (
            .O(N__28192),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_10 ));
    CascadeMux I__5112 (
            .O(N__28189),
            .I(N__28186));
    InMux I__5111 (
            .O(N__28186),
            .I(N__28179));
    InMux I__5110 (
            .O(N__28185),
            .I(N__28179));
    InMux I__5109 (
            .O(N__28184),
            .I(N__28176));
    LocalMux I__5108 (
            .O(N__28179),
            .I(N__28173));
    LocalMux I__5107 (
            .O(N__28176),
            .I(N__28170));
    Sp12to4 I__5106 (
            .O(N__28173),
            .I(N__28164));
    Span12Mux_s10_v I__5105 (
            .O(N__28170),
            .I(N__28164));
    InMux I__5104 (
            .O(N__28169),
            .I(N__28161));
    Odrv12 I__5103 (
            .O(N__28164),
            .I(\c0.FRAME_MATCHER_i_10 ));
    LocalMux I__5102 (
            .O(N__28161),
            .I(\c0.FRAME_MATCHER_i_10 ));
    SRMux I__5101 (
            .O(N__28156),
            .I(N__28153));
    LocalMux I__5100 (
            .O(N__28153),
            .I(N__28150));
    Span4Mux_h I__5099 (
            .O(N__28150),
            .I(N__28147));
    Odrv4 I__5098 (
            .O(N__28147),
            .I(\c0.n3_adj_2247 ));
    CascadeMux I__5097 (
            .O(N__28144),
            .I(\c0.n9819_cascade_ ));
    InMux I__5096 (
            .O(N__28141),
            .I(N__28136));
    InMux I__5095 (
            .O(N__28140),
            .I(N__28133));
    InMux I__5094 (
            .O(N__28139),
            .I(N__28129));
    LocalMux I__5093 (
            .O(N__28136),
            .I(N__28126));
    LocalMux I__5092 (
            .O(N__28133),
            .I(N__28123));
    InMux I__5091 (
            .O(N__28132),
            .I(N__28120));
    LocalMux I__5090 (
            .O(N__28129),
            .I(N__28117));
    Span4Mux_h I__5089 (
            .O(N__28126),
            .I(N__28114));
    Span4Mux_h I__5088 (
            .O(N__28123),
            .I(N__28111));
    LocalMux I__5087 (
            .O(N__28120),
            .I(\c0.FRAME_MATCHER_state_25 ));
    Odrv4 I__5086 (
            .O(N__28117),
            .I(\c0.FRAME_MATCHER_state_25 ));
    Odrv4 I__5085 (
            .O(N__28114),
            .I(\c0.FRAME_MATCHER_state_25 ));
    Odrv4 I__5084 (
            .O(N__28111),
            .I(\c0.FRAME_MATCHER_state_25 ));
    SRMux I__5083 (
            .O(N__28102),
            .I(N__28099));
    LocalMux I__5082 (
            .O(N__28099),
            .I(N__28096));
    Odrv12 I__5081 (
            .O(N__28096),
            .I(\c0.n16359 ));
    InMux I__5080 (
            .O(N__28093),
            .I(N__28090));
    LocalMux I__5079 (
            .O(N__28090),
            .I(N__28087));
    Odrv12 I__5078 (
            .O(N__28087),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_17 ));
    CascadeMux I__5077 (
            .O(N__28084),
            .I(N__28078));
    CascadeMux I__5076 (
            .O(N__28083),
            .I(N__28075));
    CascadeMux I__5075 (
            .O(N__28082),
            .I(N__28072));
    InMux I__5074 (
            .O(N__28081),
            .I(N__28069));
    InMux I__5073 (
            .O(N__28078),
            .I(N__28066));
    InMux I__5072 (
            .O(N__28075),
            .I(N__28063));
    InMux I__5071 (
            .O(N__28072),
            .I(N__28060));
    LocalMux I__5070 (
            .O(N__28069),
            .I(N__28057));
    LocalMux I__5069 (
            .O(N__28066),
            .I(N__28054));
    LocalMux I__5068 (
            .O(N__28063),
            .I(N__28049));
    LocalMux I__5067 (
            .O(N__28060),
            .I(N__28049));
    Span4Mux_h I__5066 (
            .O(N__28057),
            .I(N__28046));
    Span4Mux_h I__5065 (
            .O(N__28054),
            .I(N__28043));
    Odrv12 I__5064 (
            .O(N__28049),
            .I(\c0.FRAME_MATCHER_i_17 ));
    Odrv4 I__5063 (
            .O(N__28046),
            .I(\c0.FRAME_MATCHER_i_17 ));
    Odrv4 I__5062 (
            .O(N__28043),
            .I(\c0.FRAME_MATCHER_i_17 ));
    InMux I__5061 (
            .O(N__28036),
            .I(N__28033));
    LocalMux I__5060 (
            .O(N__28033),
            .I(N__28030));
    Span4Mux_h I__5059 (
            .O(N__28030),
            .I(N__28026));
    InMux I__5058 (
            .O(N__28029),
            .I(N__28023));
    Span4Mux_h I__5057 (
            .O(N__28026),
            .I(N__28020));
    LocalMux I__5056 (
            .O(N__28023),
            .I(N__28017));
    Odrv4 I__5055 (
            .O(N__28020),
            .I(n17));
    Odrv4 I__5054 (
            .O(N__28017),
            .I(n17));
    SRMux I__5053 (
            .O(N__28012),
            .I(N__28009));
    LocalMux I__5052 (
            .O(N__28009),
            .I(N__28006));
    Span4Mux_h I__5051 (
            .O(N__28006),
            .I(N__28003));
    Odrv4 I__5050 (
            .O(N__28003),
            .I(\c0.n16369 ));
    InMux I__5049 (
            .O(N__28000),
            .I(N__27997));
    LocalMux I__5048 (
            .O(N__27997),
            .I(N__27994));
    Odrv4 I__5047 (
            .O(N__27994),
            .I(\c0.n12_adj_2189 ));
    InMux I__5046 (
            .O(N__27991),
            .I(N__27987));
    InMux I__5045 (
            .O(N__27990),
            .I(N__27984));
    LocalMux I__5044 (
            .O(N__27987),
            .I(N__27978));
    LocalMux I__5043 (
            .O(N__27984),
            .I(N__27975));
    InMux I__5042 (
            .O(N__27983),
            .I(N__27972));
    InMux I__5041 (
            .O(N__27982),
            .I(N__27969));
    InMux I__5040 (
            .O(N__27981),
            .I(N__27966));
    Span4Mux_v I__5039 (
            .O(N__27978),
            .I(N__27963));
    Span4Mux_h I__5038 (
            .O(N__27975),
            .I(N__27958));
    LocalMux I__5037 (
            .O(N__27972),
            .I(N__27958));
    LocalMux I__5036 (
            .O(N__27969),
            .I(N__27955));
    LocalMux I__5035 (
            .O(N__27966),
            .I(N__27948));
    Span4Mux_h I__5034 (
            .O(N__27963),
            .I(N__27948));
    Span4Mux_v I__5033 (
            .O(N__27958),
            .I(N__27948));
    Odrv12 I__5032 (
            .O(N__27955),
            .I(\c0.FRAME_MATCHER_state_20 ));
    Odrv4 I__5031 (
            .O(N__27948),
            .I(\c0.FRAME_MATCHER_state_20 ));
    InMux I__5030 (
            .O(N__27943),
            .I(N__27940));
    LocalMux I__5029 (
            .O(N__27940),
            .I(N__27934));
    InMux I__5028 (
            .O(N__27939),
            .I(N__27931));
    InMux I__5027 (
            .O(N__27938),
            .I(N__27926));
    InMux I__5026 (
            .O(N__27937),
            .I(N__27926));
    Span4Mux_h I__5025 (
            .O(N__27934),
            .I(N__27923));
    LocalMux I__5024 (
            .O(N__27931),
            .I(N__27920));
    LocalMux I__5023 (
            .O(N__27926),
            .I(N__27917));
    Odrv4 I__5022 (
            .O(N__27923),
            .I(n9460));
    Odrv12 I__5021 (
            .O(N__27920),
            .I(n9460));
    Odrv12 I__5020 (
            .O(N__27917),
            .I(n9460));
    CascadeMux I__5019 (
            .O(N__27910),
            .I(n9460_cascade_));
    InMux I__5018 (
            .O(N__27907),
            .I(N__27903));
    InMux I__5017 (
            .O(N__27906),
            .I(N__27900));
    LocalMux I__5016 (
            .O(N__27903),
            .I(N__27897));
    LocalMux I__5015 (
            .O(N__27900),
            .I(N__27894));
    Span4Mux_h I__5014 (
            .O(N__27897),
            .I(N__27891));
    Span4Mux_h I__5013 (
            .O(N__27894),
            .I(N__27888));
    Span4Mux_h I__5012 (
            .O(N__27891),
            .I(N__27885));
    Odrv4 I__5011 (
            .O(N__27888),
            .I(n9462));
    Odrv4 I__5010 (
            .O(N__27885),
            .I(n9462));
    InMux I__5009 (
            .O(N__27880),
            .I(N__27875));
    InMux I__5008 (
            .O(N__27879),
            .I(N__27872));
    InMux I__5007 (
            .O(N__27878),
            .I(N__27869));
    LocalMux I__5006 (
            .O(N__27875),
            .I(N__27866));
    LocalMux I__5005 (
            .O(N__27872),
            .I(N__27861));
    LocalMux I__5004 (
            .O(N__27869),
            .I(N__27856));
    Span4Mux_v I__5003 (
            .O(N__27866),
            .I(N__27856));
    InMux I__5002 (
            .O(N__27865),
            .I(N__27851));
    InMux I__5001 (
            .O(N__27864),
            .I(N__27851));
    Span4Mux_h I__5000 (
            .O(N__27861),
            .I(N__27848));
    Odrv4 I__4999 (
            .O(N__27856),
            .I(\c0.FRAME_MATCHER_state_18 ));
    LocalMux I__4998 (
            .O(N__27851),
            .I(\c0.FRAME_MATCHER_state_18 ));
    Odrv4 I__4997 (
            .O(N__27848),
            .I(\c0.FRAME_MATCHER_state_18 ));
    SRMux I__4996 (
            .O(N__27841),
            .I(N__27838));
    LocalMux I__4995 (
            .O(N__27838),
            .I(\c0.n16343 ));
    InMux I__4994 (
            .O(N__27835),
            .I(N__27832));
    LocalMux I__4993 (
            .O(N__27832),
            .I(N__27829));
    Span4Mux_v I__4992 (
            .O(N__27829),
            .I(N__27825));
    InMux I__4991 (
            .O(N__27828),
            .I(N__27821));
    Span4Mux_h I__4990 (
            .O(N__27825),
            .I(N__27818));
    InMux I__4989 (
            .O(N__27824),
            .I(N__27815));
    LocalMux I__4988 (
            .O(N__27821),
            .I(data_in_2_6));
    Odrv4 I__4987 (
            .O(N__27818),
            .I(data_in_2_6));
    LocalMux I__4986 (
            .O(N__27815),
            .I(data_in_2_6));
    CascadeMux I__4985 (
            .O(N__27808),
            .I(N__27805));
    InMux I__4984 (
            .O(N__27805),
            .I(N__27791));
    InMux I__4983 (
            .O(N__27804),
            .I(N__27791));
    InMux I__4982 (
            .O(N__27803),
            .I(N__27791));
    InMux I__4981 (
            .O(N__27802),
            .I(N__27791));
    InMux I__4980 (
            .O(N__27801),
            .I(N__27787));
    InMux I__4979 (
            .O(N__27800),
            .I(N__27784));
    LocalMux I__4978 (
            .O(N__27791),
            .I(N__27779));
    InMux I__4977 (
            .O(N__27790),
            .I(N__27776));
    LocalMux I__4976 (
            .O(N__27787),
            .I(N__27771));
    LocalMux I__4975 (
            .O(N__27784),
            .I(N__27771));
    CascadeMux I__4974 (
            .O(N__27783),
            .I(N__27765));
    InMux I__4973 (
            .O(N__27782),
            .I(N__27758));
    Span4Mux_v I__4972 (
            .O(N__27779),
            .I(N__27753));
    LocalMux I__4971 (
            .O(N__27776),
            .I(N__27753));
    Span4Mux_h I__4970 (
            .O(N__27771),
            .I(N__27750));
    InMux I__4969 (
            .O(N__27770),
            .I(N__27747));
    InMux I__4968 (
            .O(N__27769),
            .I(N__27736));
    InMux I__4967 (
            .O(N__27768),
            .I(N__27736));
    InMux I__4966 (
            .O(N__27765),
            .I(N__27731));
    InMux I__4965 (
            .O(N__27764),
            .I(N__27731));
    InMux I__4964 (
            .O(N__27763),
            .I(N__27724));
    InMux I__4963 (
            .O(N__27762),
            .I(N__27724));
    InMux I__4962 (
            .O(N__27761),
            .I(N__27724));
    LocalMux I__4961 (
            .O(N__27758),
            .I(N__27721));
    Span4Mux_h I__4960 (
            .O(N__27753),
            .I(N__27714));
    Span4Mux_v I__4959 (
            .O(N__27750),
            .I(N__27714));
    LocalMux I__4958 (
            .O(N__27747),
            .I(N__27714));
    InMux I__4957 (
            .O(N__27746),
            .I(N__27695));
    InMux I__4956 (
            .O(N__27745),
            .I(N__27695));
    InMux I__4955 (
            .O(N__27744),
            .I(N__27695));
    InMux I__4954 (
            .O(N__27743),
            .I(N__27695));
    InMux I__4953 (
            .O(N__27742),
            .I(N__27690));
    InMux I__4952 (
            .O(N__27741),
            .I(N__27690));
    LocalMux I__4951 (
            .O(N__27736),
            .I(N__27687));
    LocalMux I__4950 (
            .O(N__27731),
            .I(N__27680));
    LocalMux I__4949 (
            .O(N__27724),
            .I(N__27680));
    Span4Mux_v I__4948 (
            .O(N__27721),
            .I(N__27680));
    Span4Mux_h I__4947 (
            .O(N__27714),
            .I(N__27677));
    CascadeMux I__4946 (
            .O(N__27713),
            .I(N__27674));
    InMux I__4945 (
            .O(N__27712),
            .I(N__27666));
    InMux I__4944 (
            .O(N__27711),
            .I(N__27666));
    InMux I__4943 (
            .O(N__27710),
            .I(N__27657));
    InMux I__4942 (
            .O(N__27709),
            .I(N__27657));
    InMux I__4941 (
            .O(N__27708),
            .I(N__27657));
    InMux I__4940 (
            .O(N__27707),
            .I(N__27657));
    InMux I__4939 (
            .O(N__27706),
            .I(N__27650));
    InMux I__4938 (
            .O(N__27705),
            .I(N__27650));
    InMux I__4937 (
            .O(N__27704),
            .I(N__27650));
    LocalMux I__4936 (
            .O(N__27695),
            .I(N__27647));
    LocalMux I__4935 (
            .O(N__27690),
            .I(N__27644));
    Span4Mux_h I__4934 (
            .O(N__27687),
            .I(N__27641));
    Span4Mux_h I__4933 (
            .O(N__27680),
            .I(N__27636));
    Span4Mux_v I__4932 (
            .O(N__27677),
            .I(N__27636));
    InMux I__4931 (
            .O(N__27674),
            .I(N__27627));
    InMux I__4930 (
            .O(N__27673),
            .I(N__27627));
    InMux I__4929 (
            .O(N__27672),
            .I(N__27627));
    InMux I__4928 (
            .O(N__27671),
            .I(N__27627));
    LocalMux I__4927 (
            .O(N__27666),
            .I(rx_data_ready));
    LocalMux I__4926 (
            .O(N__27657),
            .I(rx_data_ready));
    LocalMux I__4925 (
            .O(N__27650),
            .I(rx_data_ready));
    Odrv4 I__4924 (
            .O(N__27647),
            .I(rx_data_ready));
    Odrv12 I__4923 (
            .O(N__27644),
            .I(rx_data_ready));
    Odrv4 I__4922 (
            .O(N__27641),
            .I(rx_data_ready));
    Odrv4 I__4921 (
            .O(N__27636),
            .I(rx_data_ready));
    LocalMux I__4920 (
            .O(N__27627),
            .I(rx_data_ready));
    InMux I__4919 (
            .O(N__27610),
            .I(N__27605));
    InMux I__4918 (
            .O(N__27609),
            .I(N__27600));
    InMux I__4917 (
            .O(N__27608),
            .I(N__27600));
    LocalMux I__4916 (
            .O(N__27605),
            .I(N__27597));
    LocalMux I__4915 (
            .O(N__27600),
            .I(N__27593));
    Span12Mux_s8_h I__4914 (
            .O(N__27597),
            .I(N__27590));
    InMux I__4913 (
            .O(N__27596),
            .I(N__27587));
    Span4Mux_h I__4912 (
            .O(N__27593),
            .I(N__27584));
    Odrv12 I__4911 (
            .O(N__27590),
            .I(data_in_1_6));
    LocalMux I__4910 (
            .O(N__27587),
            .I(data_in_1_6));
    Odrv4 I__4909 (
            .O(N__27584),
            .I(data_in_1_6));
    InMux I__4908 (
            .O(N__27577),
            .I(N__27570));
    InMux I__4907 (
            .O(N__27576),
            .I(N__27565));
    InMux I__4906 (
            .O(N__27575),
            .I(N__27560));
    InMux I__4905 (
            .O(N__27574),
            .I(N__27560));
    CascadeMux I__4904 (
            .O(N__27573),
            .I(N__27553));
    LocalMux I__4903 (
            .O(N__27570),
            .I(N__27545));
    InMux I__4902 (
            .O(N__27569),
            .I(N__27540));
    InMux I__4901 (
            .O(N__27568),
            .I(N__27540));
    LocalMux I__4900 (
            .O(N__27565),
            .I(N__27535));
    LocalMux I__4899 (
            .O(N__27560),
            .I(N__27535));
    InMux I__4898 (
            .O(N__27559),
            .I(N__27529));
    InMux I__4897 (
            .O(N__27558),
            .I(N__27520));
    InMux I__4896 (
            .O(N__27557),
            .I(N__27520));
    InMux I__4895 (
            .O(N__27556),
            .I(N__27520));
    InMux I__4894 (
            .O(N__27553),
            .I(N__27520));
    InMux I__4893 (
            .O(N__27552),
            .I(N__27515));
    InMux I__4892 (
            .O(N__27551),
            .I(N__27515));
    InMux I__4891 (
            .O(N__27550),
            .I(N__27510));
    InMux I__4890 (
            .O(N__27549),
            .I(N__27510));
    InMux I__4889 (
            .O(N__27548),
            .I(N__27507));
    Span4Mux_v I__4888 (
            .O(N__27545),
            .I(N__27500));
    LocalMux I__4887 (
            .O(N__27540),
            .I(N__27500));
    Span4Mux_s1_v I__4886 (
            .O(N__27535),
            .I(N__27500));
    InMux I__4885 (
            .O(N__27534),
            .I(N__27495));
    InMux I__4884 (
            .O(N__27533),
            .I(N__27495));
    InMux I__4883 (
            .O(N__27532),
            .I(N__27492));
    LocalMux I__4882 (
            .O(N__27529),
            .I(n29));
    LocalMux I__4881 (
            .O(N__27520),
            .I(n29));
    LocalMux I__4880 (
            .O(N__27515),
            .I(n29));
    LocalMux I__4879 (
            .O(N__27510),
            .I(n29));
    LocalMux I__4878 (
            .O(N__27507),
            .I(n29));
    Odrv4 I__4877 (
            .O(N__27500),
            .I(n29));
    LocalMux I__4876 (
            .O(N__27495),
            .I(n29));
    LocalMux I__4875 (
            .O(N__27492),
            .I(n29));
    CascadeMux I__4874 (
            .O(N__27475),
            .I(N__27472));
    InMux I__4873 (
            .O(N__27472),
            .I(N__27468));
    InMux I__4872 (
            .O(N__27471),
            .I(N__27465));
    LocalMux I__4871 (
            .O(N__27468),
            .I(N__27461));
    LocalMux I__4870 (
            .O(N__27465),
            .I(N__27458));
    CascadeMux I__4869 (
            .O(N__27464),
            .I(N__27455));
    Span4Mux_s3_v I__4868 (
            .O(N__27461),
            .I(N__27452));
    Span4Mux_h I__4867 (
            .O(N__27458),
            .I(N__27449));
    InMux I__4866 (
            .O(N__27455),
            .I(N__27446));
    Span4Mux_h I__4865 (
            .O(N__27452),
            .I(N__27443));
    Sp12to4 I__4864 (
            .O(N__27449),
            .I(N__27438));
    LocalMux I__4863 (
            .O(N__27446),
            .I(N__27438));
    Span4Mux_v I__4862 (
            .O(N__27443),
            .I(N__27435));
    Span12Mux_s10_v I__4861 (
            .O(N__27438),
            .I(N__27432));
    Odrv4 I__4860 (
            .O(N__27435),
            .I(n445));
    Odrv12 I__4859 (
            .O(N__27432),
            .I(n445));
    InMux I__4858 (
            .O(N__27427),
            .I(N__27422));
    InMux I__4857 (
            .O(N__27426),
            .I(N__27417));
    InMux I__4856 (
            .O(N__27425),
            .I(N__27417));
    LocalMux I__4855 (
            .O(N__27422),
            .I(n10031));
    LocalMux I__4854 (
            .O(N__27417),
            .I(n10031));
    CascadeMux I__4853 (
            .O(N__27412),
            .I(n17479_cascade_));
    InMux I__4852 (
            .O(N__27409),
            .I(N__27406));
    LocalMux I__4851 (
            .O(N__27406),
            .I(N__27403));
    Span4Mux_h I__4850 (
            .O(N__27403),
            .I(N__27399));
    InMux I__4849 (
            .O(N__27402),
            .I(N__27396));
    Odrv4 I__4848 (
            .O(N__27399),
            .I(n16886));
    LocalMux I__4847 (
            .O(N__27396),
            .I(n16886));
    InMux I__4846 (
            .O(N__27391),
            .I(N__27388));
    LocalMux I__4845 (
            .O(N__27388),
            .I(n38));
    InMux I__4844 (
            .O(N__27385),
            .I(N__27382));
    LocalMux I__4843 (
            .O(N__27382),
            .I(\c0.n44_adj_2163 ));
    InMux I__4842 (
            .O(N__27379),
            .I(N__27366));
    InMux I__4841 (
            .O(N__27378),
            .I(N__27366));
    InMux I__4840 (
            .O(N__27377),
            .I(N__27366));
    InMux I__4839 (
            .O(N__27376),
            .I(N__27366));
    InMux I__4838 (
            .O(N__27375),
            .I(N__27363));
    LocalMux I__4837 (
            .O(N__27366),
            .I(n9357));
    LocalMux I__4836 (
            .O(N__27363),
            .I(n9357));
    CascadeMux I__4835 (
            .O(N__27358),
            .I(N__27354));
    InMux I__4834 (
            .O(N__27357),
            .I(N__27349));
    InMux I__4833 (
            .O(N__27354),
            .I(N__27344));
    InMux I__4832 (
            .O(N__27353),
            .I(N__27339));
    InMux I__4831 (
            .O(N__27352),
            .I(N__27339));
    LocalMux I__4830 (
            .O(N__27349),
            .I(N__27335));
    InMux I__4829 (
            .O(N__27348),
            .I(N__27330));
    InMux I__4828 (
            .O(N__27347),
            .I(N__27330));
    LocalMux I__4827 (
            .O(N__27344),
            .I(N__27325));
    LocalMux I__4826 (
            .O(N__27339),
            .I(N__27325));
    InMux I__4825 (
            .O(N__27338),
            .I(N__27322));
    Odrv4 I__4824 (
            .O(N__27335),
            .I(\c0.tx_transmit_N_1949_2 ));
    LocalMux I__4823 (
            .O(N__27330),
            .I(\c0.tx_transmit_N_1949_2 ));
    Odrv4 I__4822 (
            .O(N__27325),
            .I(\c0.tx_transmit_N_1949_2 ));
    LocalMux I__4821 (
            .O(N__27322),
            .I(\c0.tx_transmit_N_1949_2 ));
    InMux I__4820 (
            .O(N__27313),
            .I(N__27303));
    InMux I__4819 (
            .O(N__27312),
            .I(N__27303));
    InMux I__4818 (
            .O(N__27311),
            .I(N__27300));
    InMux I__4817 (
            .O(N__27310),
            .I(N__27297));
    InMux I__4816 (
            .O(N__27309),
            .I(N__27294));
    InMux I__4815 (
            .O(N__27308),
            .I(N__27291));
    LocalMux I__4814 (
            .O(N__27303),
            .I(\c0.n4_adj_2311 ));
    LocalMux I__4813 (
            .O(N__27300),
            .I(\c0.n4_adj_2311 ));
    LocalMux I__4812 (
            .O(N__27297),
            .I(\c0.n4_adj_2311 ));
    LocalMux I__4811 (
            .O(N__27294),
            .I(\c0.n4_adj_2311 ));
    LocalMux I__4810 (
            .O(N__27291),
            .I(\c0.n4_adj_2311 ));
    InMux I__4809 (
            .O(N__27280),
            .I(N__27277));
    LocalMux I__4808 (
            .O(N__27277),
            .I(N__27274));
    Odrv12 I__4807 (
            .O(N__27274),
            .I(\c0.n17475 ));
    CascadeMux I__4806 (
            .O(N__27271),
            .I(\c0.tx2_transmit_N_1997_cascade_ ));
    InMux I__4805 (
            .O(N__27268),
            .I(N__27265));
    LocalMux I__4804 (
            .O(N__27265),
            .I(\c0.tx2.n113 ));
    CascadeMux I__4803 (
            .O(N__27262),
            .I(\c0.tx2.n113_cascade_ ));
    CascadeMux I__4802 (
            .O(N__27259),
            .I(N__27256));
    InMux I__4801 (
            .O(N__27256),
            .I(N__27253));
    LocalMux I__4800 (
            .O(N__27253),
            .I(N__27250));
    Span4Mux_v I__4799 (
            .O(N__27250),
            .I(N__27245));
    InMux I__4798 (
            .O(N__27249),
            .I(N__27242));
    InMux I__4797 (
            .O(N__27248),
            .I(N__27239));
    Span4Mux_h I__4796 (
            .O(N__27245),
            .I(N__27236));
    LocalMux I__4795 (
            .O(N__27242),
            .I(N__27231));
    LocalMux I__4794 (
            .O(N__27239),
            .I(N__27231));
    Span4Mux_h I__4793 (
            .O(N__27236),
            .I(N__27226));
    Span12Mux_v I__4792 (
            .O(N__27231),
            .I(N__27223));
    InMux I__4791 (
            .O(N__27230),
            .I(N__27218));
    InMux I__4790 (
            .O(N__27229),
            .I(N__27218));
    Span4Mux_v I__4789 (
            .O(N__27226),
            .I(N__27215));
    Odrv12 I__4788 (
            .O(N__27223),
            .I(\c0.r_SM_Main_2_N_2036_0_adj_2261 ));
    LocalMux I__4787 (
            .O(N__27218),
            .I(\c0.r_SM_Main_2_N_2036_0_adj_2261 ));
    Odrv4 I__4786 (
            .O(N__27215),
            .I(\c0.r_SM_Main_2_N_2036_0_adj_2261 ));
    InMux I__4785 (
            .O(N__27208),
            .I(N__27205));
    LocalMux I__4784 (
            .O(N__27205),
            .I(N__27202));
    Span4Mux_h I__4783 (
            .O(N__27202),
            .I(N__27199));
    Odrv4 I__4782 (
            .O(N__27199),
            .I(n491));
    CascadeMux I__4781 (
            .O(N__27196),
            .I(n491_cascade_));
    InMux I__4780 (
            .O(N__27193),
            .I(N__27190));
    LocalMux I__4779 (
            .O(N__27190),
            .I(N__27185));
    InMux I__4778 (
            .O(N__27189),
            .I(N__27182));
    InMux I__4777 (
            .O(N__27188),
            .I(N__27179));
    Odrv4 I__4776 (
            .O(N__27185),
            .I(\c0.n8938 ));
    LocalMux I__4775 (
            .O(N__27182),
            .I(\c0.n8938 ));
    LocalMux I__4774 (
            .O(N__27179),
            .I(\c0.n8938 ));
    InMux I__4773 (
            .O(N__27172),
            .I(N__27165));
    InMux I__4772 (
            .O(N__27171),
            .I(N__27160));
    InMux I__4771 (
            .O(N__27170),
            .I(N__27160));
    InMux I__4770 (
            .O(N__27169),
            .I(N__27155));
    InMux I__4769 (
            .O(N__27168),
            .I(N__27155));
    LocalMux I__4768 (
            .O(N__27165),
            .I(\c0.tx_transmit_N_1949_3 ));
    LocalMux I__4767 (
            .O(N__27160),
            .I(\c0.tx_transmit_N_1949_3 ));
    LocalMux I__4766 (
            .O(N__27155),
            .I(\c0.tx_transmit_N_1949_3 ));
    InMux I__4765 (
            .O(N__27148),
            .I(N__27135));
    InMux I__4764 (
            .O(N__27147),
            .I(N__27135));
    InMux I__4763 (
            .O(N__27146),
            .I(N__27135));
    InMux I__4762 (
            .O(N__27145),
            .I(N__27132));
    InMux I__4761 (
            .O(N__27144),
            .I(N__27125));
    InMux I__4760 (
            .O(N__27143),
            .I(N__27125));
    InMux I__4759 (
            .O(N__27142),
            .I(N__27125));
    LocalMux I__4758 (
            .O(N__27135),
            .I(\c0.n16839 ));
    LocalMux I__4757 (
            .O(N__27132),
            .I(\c0.n16839 ));
    LocalMux I__4756 (
            .O(N__27125),
            .I(\c0.n16839 ));
    InMux I__4755 (
            .O(N__27118),
            .I(N__27114));
    InMux I__4754 (
            .O(N__27117),
            .I(N__27111));
    LocalMux I__4753 (
            .O(N__27114),
            .I(\c0.tx_transmit_N_1949_7 ));
    LocalMux I__4752 (
            .O(N__27111),
            .I(\c0.tx_transmit_N_1949_7 ));
    InMux I__4751 (
            .O(N__27106),
            .I(N__27102));
    InMux I__4750 (
            .O(N__27105),
            .I(N__27099));
    LocalMux I__4749 (
            .O(N__27102),
            .I(\c0.byte_transmit_counter_7 ));
    LocalMux I__4748 (
            .O(N__27099),
            .I(\c0.byte_transmit_counter_7 ));
    CascadeMux I__4747 (
            .O(N__27094),
            .I(n17834_cascade_));
    InMux I__4746 (
            .O(N__27091),
            .I(N__27088));
    LocalMux I__4745 (
            .O(N__27088),
            .I(n17162));
    CascadeMux I__4744 (
            .O(N__27085),
            .I(n9358_cascade_));
    CascadeMux I__4743 (
            .O(N__27082),
            .I(n41_cascade_));
    InMux I__4742 (
            .O(N__27079),
            .I(N__27076));
    LocalMux I__4741 (
            .O(N__27076),
            .I(n35));
    InMux I__4740 (
            .O(N__27073),
            .I(N__27070));
    LocalMux I__4739 (
            .O(N__27070),
            .I(\c0.n17254 ));
    CascadeMux I__4738 (
            .O(N__27067),
            .I(\c0.n17254_cascade_ ));
    InMux I__4737 (
            .O(N__27064),
            .I(N__27061));
    LocalMux I__4736 (
            .O(N__27061),
            .I(N__27058));
    Span4Mux_s2_v I__4735 (
            .O(N__27058),
            .I(N__27055));
    Odrv4 I__4734 (
            .O(N__27055),
            .I(\c0.n17290 ));
    CascadeMux I__4733 (
            .O(N__27052),
            .I(N__27049));
    InMux I__4732 (
            .O(N__27049),
            .I(N__27043));
    InMux I__4731 (
            .O(N__27048),
            .I(N__27043));
    LocalMux I__4730 (
            .O(N__27043),
            .I(\c0.tx_transmit_N_1949_5 ));
    InMux I__4729 (
            .O(N__27040),
            .I(N__27036));
    InMux I__4728 (
            .O(N__27039),
            .I(N__27033));
    LocalMux I__4727 (
            .O(N__27036),
            .I(\c0.n5_adj_2319 ));
    LocalMux I__4726 (
            .O(N__27033),
            .I(\c0.n5_adj_2319 ));
    InMux I__4725 (
            .O(N__27028),
            .I(N__27021));
    InMux I__4724 (
            .O(N__27027),
            .I(N__27021));
    InMux I__4723 (
            .O(N__27026),
            .I(N__27018));
    LocalMux I__4722 (
            .O(N__27021),
            .I(\c0.tx_transmit_N_1949_6 ));
    LocalMux I__4721 (
            .O(N__27018),
            .I(\c0.tx_transmit_N_1949_6 ));
    InMux I__4720 (
            .O(N__27013),
            .I(N__27009));
    InMux I__4719 (
            .O(N__27012),
            .I(N__27006));
    LocalMux I__4718 (
            .O(N__27009),
            .I(\c0.byte_transmit_counter_6 ));
    LocalMux I__4717 (
            .O(N__27006),
            .I(\c0.byte_transmit_counter_6 ));
    InMux I__4716 (
            .O(N__27001),
            .I(N__26998));
    LocalMux I__4715 (
            .O(N__26998),
            .I(\c0.n23_adj_2309 ));
    InMux I__4714 (
            .O(N__26995),
            .I(N__26992));
    LocalMux I__4713 (
            .O(N__26992),
            .I(N__26989));
    Odrv12 I__4712 (
            .O(N__26989),
            .I(\c0.n17278 ));
    InMux I__4711 (
            .O(N__26986),
            .I(N__26983));
    LocalMux I__4710 (
            .O(N__26983),
            .I(N__26980));
    Span4Mux_s2_v I__4709 (
            .O(N__26980),
            .I(N__26977));
    Odrv4 I__4708 (
            .O(N__26977),
            .I(\c0.n17276 ));
    InMux I__4707 (
            .O(N__26974),
            .I(N__26970));
    InMux I__4706 (
            .O(N__26973),
            .I(N__26967));
    LocalMux I__4705 (
            .O(N__26970),
            .I(\c0.tx_transmit_N_1949_0 ));
    LocalMux I__4704 (
            .O(N__26967),
            .I(\c0.tx_transmit_N_1949_0 ));
    CascadeMux I__4703 (
            .O(N__26962),
            .I(\c0.n16839_cascade_ ));
    InMux I__4702 (
            .O(N__26959),
            .I(N__26954));
    InMux I__4701 (
            .O(N__26958),
            .I(N__26951));
    InMux I__4700 (
            .O(N__26957),
            .I(N__26948));
    LocalMux I__4699 (
            .O(N__26954),
            .I(\c0.tx_transmit_N_1949_4 ));
    LocalMux I__4698 (
            .O(N__26951),
            .I(\c0.tx_transmit_N_1949_4 ));
    LocalMux I__4697 (
            .O(N__26948),
            .I(\c0.tx_transmit_N_1949_4 ));
    CascadeMux I__4696 (
            .O(N__26941),
            .I(N__26937));
    CascadeMux I__4695 (
            .O(N__26940),
            .I(N__26933));
    InMux I__4694 (
            .O(N__26937),
            .I(N__26929));
    InMux I__4693 (
            .O(N__26936),
            .I(N__26926));
    InMux I__4692 (
            .O(N__26933),
            .I(N__26923));
    CascadeMux I__4691 (
            .O(N__26932),
            .I(N__26920));
    LocalMux I__4690 (
            .O(N__26929),
            .I(N__26915));
    LocalMux I__4689 (
            .O(N__26926),
            .I(N__26912));
    LocalMux I__4688 (
            .O(N__26923),
            .I(N__26907));
    InMux I__4687 (
            .O(N__26920),
            .I(N__26902));
    InMux I__4686 (
            .O(N__26919),
            .I(N__26902));
    CascadeMux I__4685 (
            .O(N__26918),
            .I(N__26898));
    Span4Mux_v I__4684 (
            .O(N__26915),
            .I(N__26895));
    Span4Mux_h I__4683 (
            .O(N__26912),
            .I(N__26892));
    InMux I__4682 (
            .O(N__26911),
            .I(N__26889));
    InMux I__4681 (
            .O(N__26910),
            .I(N__26886));
    Span4Mux_h I__4680 (
            .O(N__26907),
            .I(N__26881));
    LocalMux I__4679 (
            .O(N__26902),
            .I(N__26881));
    InMux I__4678 (
            .O(N__26901),
            .I(N__26878));
    InMux I__4677 (
            .O(N__26898),
            .I(N__26875));
    Odrv4 I__4676 (
            .O(N__26895),
            .I(rx_data_2));
    Odrv4 I__4675 (
            .O(N__26892),
            .I(rx_data_2));
    LocalMux I__4674 (
            .O(N__26889),
            .I(rx_data_2));
    LocalMux I__4673 (
            .O(N__26886),
            .I(rx_data_2));
    Odrv4 I__4672 (
            .O(N__26881),
            .I(rx_data_2));
    LocalMux I__4671 (
            .O(N__26878),
            .I(rx_data_2));
    LocalMux I__4670 (
            .O(N__26875),
            .I(rx_data_2));
    InMux I__4669 (
            .O(N__26860),
            .I(N__26853));
    InMux I__4668 (
            .O(N__26859),
            .I(N__26853));
    InMux I__4667 (
            .O(N__26858),
            .I(N__26848));
    LocalMux I__4666 (
            .O(N__26853),
            .I(N__26845));
    InMux I__4665 (
            .O(N__26852),
            .I(N__26840));
    InMux I__4664 (
            .O(N__26851),
            .I(N__26840));
    LocalMux I__4663 (
            .O(N__26848),
            .I(data_in_frame_0_0));
    Odrv4 I__4662 (
            .O(N__26845),
            .I(data_in_frame_0_0));
    LocalMux I__4661 (
            .O(N__26840),
            .I(data_in_frame_0_0));
    CascadeMux I__4660 (
            .O(N__26833),
            .I(N__26828));
    InMux I__4659 (
            .O(N__26832),
            .I(N__26825));
    InMux I__4658 (
            .O(N__26831),
            .I(N__26821));
    InMux I__4657 (
            .O(N__26828),
            .I(N__26817));
    LocalMux I__4656 (
            .O(N__26825),
            .I(N__26814));
    InMux I__4655 (
            .O(N__26824),
            .I(N__26811));
    LocalMux I__4654 (
            .O(N__26821),
            .I(N__26808));
    InMux I__4653 (
            .O(N__26820),
            .I(N__26805));
    LocalMux I__4652 (
            .O(N__26817),
            .I(\c0.data_in_frame_1_6 ));
    Odrv4 I__4651 (
            .O(N__26814),
            .I(\c0.data_in_frame_1_6 ));
    LocalMux I__4650 (
            .O(N__26811),
            .I(\c0.data_in_frame_1_6 ));
    Odrv4 I__4649 (
            .O(N__26808),
            .I(\c0.data_in_frame_1_6 ));
    LocalMux I__4648 (
            .O(N__26805),
            .I(\c0.data_in_frame_1_6 ));
    CascadeMux I__4647 (
            .O(N__26794),
            .I(N__26790));
    InMux I__4646 (
            .O(N__26793),
            .I(N__26785));
    InMux I__4645 (
            .O(N__26790),
            .I(N__26785));
    LocalMux I__4644 (
            .O(N__26785),
            .I(\c0.data_in_frame_10_2 ));
    InMux I__4643 (
            .O(N__26782),
            .I(N__26775));
    InMux I__4642 (
            .O(N__26781),
            .I(N__26775));
    InMux I__4641 (
            .O(N__26780),
            .I(N__26770));
    LocalMux I__4640 (
            .O(N__26775),
            .I(N__26767));
    InMux I__4639 (
            .O(N__26774),
            .I(N__26762));
    InMux I__4638 (
            .O(N__26773),
            .I(N__26762));
    LocalMux I__4637 (
            .O(N__26770),
            .I(data_in_frame_0_1));
    Odrv4 I__4636 (
            .O(N__26767),
            .I(data_in_frame_0_1));
    LocalMux I__4635 (
            .O(N__26762),
            .I(data_in_frame_0_1));
    InMux I__4634 (
            .O(N__26755),
            .I(N__26752));
    LocalMux I__4633 (
            .O(N__26752),
            .I(\c0.n17460 ));
    InMux I__4632 (
            .O(N__26749),
            .I(N__26746));
    LocalMux I__4631 (
            .O(N__26746),
            .I(N__26742));
    InMux I__4630 (
            .O(N__26745),
            .I(N__26739));
    Odrv4 I__4629 (
            .O(N__26742),
            .I(r_Tx_Data_3));
    LocalMux I__4628 (
            .O(N__26739),
            .I(r_Tx_Data_3));
    InMux I__4627 (
            .O(N__26734),
            .I(N__26729));
    InMux I__4626 (
            .O(N__26733),
            .I(N__26726));
    InMux I__4625 (
            .O(N__26732),
            .I(N__26722));
    LocalMux I__4624 (
            .O(N__26729),
            .I(N__26719));
    LocalMux I__4623 (
            .O(N__26726),
            .I(N__26716));
    InMux I__4622 (
            .O(N__26725),
            .I(N__26713));
    LocalMux I__4621 (
            .O(N__26722),
            .I(\c0.delay_counter_13 ));
    Odrv12 I__4620 (
            .O(N__26719),
            .I(\c0.delay_counter_13 ));
    Odrv4 I__4619 (
            .O(N__26716),
            .I(\c0.delay_counter_13 ));
    LocalMux I__4618 (
            .O(N__26713),
            .I(\c0.delay_counter_13 ));
    InMux I__4617 (
            .O(N__26704),
            .I(N__26700));
    InMux I__4616 (
            .O(N__26703),
            .I(N__26695));
    LocalMux I__4615 (
            .O(N__26700),
            .I(N__26692));
    InMux I__4614 (
            .O(N__26699),
            .I(N__26689));
    InMux I__4613 (
            .O(N__26698),
            .I(N__26686));
    LocalMux I__4612 (
            .O(N__26695),
            .I(N__26679));
    Span4Mux_h I__4611 (
            .O(N__26692),
            .I(N__26679));
    LocalMux I__4610 (
            .O(N__26689),
            .I(N__26679));
    LocalMux I__4609 (
            .O(N__26686),
            .I(\c0.delay_counter_8 ));
    Odrv4 I__4608 (
            .O(N__26679),
            .I(\c0.delay_counter_8 ));
    InMux I__4607 (
            .O(N__26674),
            .I(N__26671));
    LocalMux I__4606 (
            .O(N__26671),
            .I(N__26665));
    InMux I__4605 (
            .O(N__26670),
            .I(N__26662));
    InMux I__4604 (
            .O(N__26669),
            .I(N__26657));
    InMux I__4603 (
            .O(N__26668),
            .I(N__26657));
    Odrv12 I__4602 (
            .O(N__26665),
            .I(\c0.delay_counter_4 ));
    LocalMux I__4601 (
            .O(N__26662),
            .I(\c0.delay_counter_4 ));
    LocalMux I__4600 (
            .O(N__26657),
            .I(\c0.delay_counter_4 ));
    CascadeMux I__4599 (
            .O(N__26650),
            .I(N__26646));
    InMux I__4598 (
            .O(N__26649),
            .I(N__26642));
    InMux I__4597 (
            .O(N__26646),
            .I(N__26639));
    InMux I__4596 (
            .O(N__26645),
            .I(N__26636));
    LocalMux I__4595 (
            .O(N__26642),
            .I(N__26632));
    LocalMux I__4594 (
            .O(N__26639),
            .I(N__26627));
    LocalMux I__4593 (
            .O(N__26636),
            .I(N__26627));
    InMux I__4592 (
            .O(N__26635),
            .I(N__26624));
    Span4Mux_s1_v I__4591 (
            .O(N__26632),
            .I(N__26621));
    Odrv4 I__4590 (
            .O(N__26627),
            .I(\c0.delay_counter_2 ));
    LocalMux I__4589 (
            .O(N__26624),
            .I(\c0.delay_counter_2 ));
    Odrv4 I__4588 (
            .O(N__26621),
            .I(\c0.delay_counter_2 ));
    CascadeMux I__4587 (
            .O(N__26614),
            .I(N__26611));
    InMux I__4586 (
            .O(N__26611),
            .I(N__26608));
    LocalMux I__4585 (
            .O(N__26608),
            .I(N__26605));
    Odrv4 I__4584 (
            .O(N__26605),
            .I(\c0.n17236 ));
    InMux I__4583 (
            .O(N__26602),
            .I(N__26599));
    LocalMux I__4582 (
            .O(N__26599),
            .I(\c0.n42_adj_2165 ));
    CascadeMux I__4581 (
            .O(N__26596),
            .I(N__26592));
    InMux I__4580 (
            .O(N__26595),
            .I(N__26589));
    InMux I__4579 (
            .O(N__26592),
            .I(N__26586));
    LocalMux I__4578 (
            .O(N__26589),
            .I(\c0.byte_transmit_counter_5 ));
    LocalMux I__4577 (
            .O(N__26586),
            .I(\c0.byte_transmit_counter_5 ));
    InMux I__4576 (
            .O(N__26581),
            .I(N__26578));
    LocalMux I__4575 (
            .O(N__26578),
            .I(N__26574));
    InMux I__4574 (
            .O(N__26577),
            .I(N__26571));
    Span4Mux_v I__4573 (
            .O(N__26574),
            .I(N__26568));
    LocalMux I__4572 (
            .O(N__26571),
            .I(data_in_frame_7_2));
    Odrv4 I__4571 (
            .O(N__26568),
            .I(data_in_frame_7_2));
    InMux I__4570 (
            .O(N__26563),
            .I(N__26559));
    InMux I__4569 (
            .O(N__26562),
            .I(N__26556));
    LocalMux I__4568 (
            .O(N__26559),
            .I(N__26553));
    LocalMux I__4567 (
            .O(N__26556),
            .I(data_in_frame_6_2));
    Odrv4 I__4566 (
            .O(N__26553),
            .I(data_in_frame_6_2));
    CascadeMux I__4565 (
            .O(N__26548),
            .I(\c0.n22_cascade_ ));
    InMux I__4564 (
            .O(N__26545),
            .I(N__26542));
    LocalMux I__4563 (
            .O(N__26542),
            .I(\c0.n27 ));
    CascadeMux I__4562 (
            .O(N__26539),
            .I(N__26533));
    CascadeMux I__4561 (
            .O(N__26538),
            .I(N__26529));
    CascadeMux I__4560 (
            .O(N__26537),
            .I(N__26526));
    CascadeMux I__4559 (
            .O(N__26536),
            .I(N__26522));
    InMux I__4558 (
            .O(N__26533),
            .I(N__26517));
    InMux I__4557 (
            .O(N__26532),
            .I(N__26514));
    InMux I__4556 (
            .O(N__26529),
            .I(N__26511));
    InMux I__4555 (
            .O(N__26526),
            .I(N__26508));
    InMux I__4554 (
            .O(N__26525),
            .I(N__26505));
    InMux I__4553 (
            .O(N__26522),
            .I(N__26502));
    InMux I__4552 (
            .O(N__26521),
            .I(N__26499));
    InMux I__4551 (
            .O(N__26520),
            .I(N__26496));
    LocalMux I__4550 (
            .O(N__26517),
            .I(N__26491));
    LocalMux I__4549 (
            .O(N__26514),
            .I(N__26491));
    LocalMux I__4548 (
            .O(N__26511),
            .I(N__26485));
    LocalMux I__4547 (
            .O(N__26508),
            .I(N__26485));
    LocalMux I__4546 (
            .O(N__26505),
            .I(N__26482));
    LocalMux I__4545 (
            .O(N__26502),
            .I(N__26477));
    LocalMux I__4544 (
            .O(N__26499),
            .I(N__26477));
    LocalMux I__4543 (
            .O(N__26496),
            .I(N__26474));
    Span4Mux_v I__4542 (
            .O(N__26491),
            .I(N__26471));
    CascadeMux I__4541 (
            .O(N__26490),
            .I(N__26468));
    Span4Mux_v I__4540 (
            .O(N__26485),
            .I(N__26465));
    Span4Mux_h I__4539 (
            .O(N__26482),
            .I(N__26462));
    Span12Mux_h I__4538 (
            .O(N__26477),
            .I(N__26459));
    Span4Mux_v I__4537 (
            .O(N__26474),
            .I(N__26456));
    Span4Mux_s3_h I__4536 (
            .O(N__26471),
            .I(N__26453));
    InMux I__4535 (
            .O(N__26468),
            .I(N__26450));
    Odrv4 I__4534 (
            .O(N__26465),
            .I(rx_data_7));
    Odrv4 I__4533 (
            .O(N__26462),
            .I(rx_data_7));
    Odrv12 I__4532 (
            .O(N__26459),
            .I(rx_data_7));
    Odrv4 I__4531 (
            .O(N__26456),
            .I(rx_data_7));
    Odrv4 I__4530 (
            .O(N__26453),
            .I(rx_data_7));
    LocalMux I__4529 (
            .O(N__26450),
            .I(rx_data_7));
    InMux I__4528 (
            .O(N__26437),
            .I(N__26432));
    CascadeMux I__4527 (
            .O(N__26436),
            .I(N__26429));
    InMux I__4526 (
            .O(N__26435),
            .I(N__26425));
    LocalMux I__4525 (
            .O(N__26432),
            .I(N__26422));
    InMux I__4524 (
            .O(N__26429),
            .I(N__26419));
    InMux I__4523 (
            .O(N__26428),
            .I(N__26416));
    LocalMux I__4522 (
            .O(N__26425),
            .I(N__26413));
    Span4Mux_h I__4521 (
            .O(N__26422),
            .I(N__26410));
    LocalMux I__4520 (
            .O(N__26419),
            .I(\c0.data_in_frame_1_0 ));
    LocalMux I__4519 (
            .O(N__26416),
            .I(\c0.data_in_frame_1_0 ));
    Odrv4 I__4518 (
            .O(N__26413),
            .I(\c0.data_in_frame_1_0 ));
    Odrv4 I__4517 (
            .O(N__26410),
            .I(\c0.data_in_frame_1_0 ));
    InMux I__4516 (
            .O(N__26401),
            .I(N__26398));
    LocalMux I__4515 (
            .O(N__26398),
            .I(N__26395));
    Odrv12 I__4514 (
            .O(N__26395),
            .I(n17634));
    InMux I__4513 (
            .O(N__26392),
            .I(N__26383));
    InMux I__4512 (
            .O(N__26391),
            .I(N__26383));
    InMux I__4511 (
            .O(N__26390),
            .I(N__26383));
    LocalMux I__4510 (
            .O(N__26383),
            .I(N__26379));
    InMux I__4509 (
            .O(N__26382),
            .I(N__26375));
    Span4Mux_s3_h I__4508 (
            .O(N__26379),
            .I(N__26372));
    InMux I__4507 (
            .O(N__26378),
            .I(N__26369));
    LocalMux I__4506 (
            .O(N__26375),
            .I(N__26366));
    Span4Mux_h I__4505 (
            .O(N__26372),
            .I(N__26363));
    LocalMux I__4504 (
            .O(N__26369),
            .I(r_Clock_Count_6_adj_2448));
    Odrv12 I__4503 (
            .O(N__26366),
            .I(r_Clock_Count_6_adj_2448));
    Odrv4 I__4502 (
            .O(N__26363),
            .I(r_Clock_Count_6_adj_2448));
    InMux I__4501 (
            .O(N__26356),
            .I(N__26353));
    LocalMux I__4500 (
            .O(N__26353),
            .I(\c0.n9585 ));
    InMux I__4499 (
            .O(N__26350),
            .I(N__26346));
    InMux I__4498 (
            .O(N__26349),
            .I(N__26343));
    LocalMux I__4497 (
            .O(N__26346),
            .I(N__26340));
    LocalMux I__4496 (
            .O(N__26343),
            .I(\c0.data_in_frame_2_2 ));
    Odrv4 I__4495 (
            .O(N__26340),
            .I(\c0.data_in_frame_2_2 ));
    InMux I__4494 (
            .O(N__26335),
            .I(N__26332));
    LocalMux I__4493 (
            .O(N__26332),
            .I(\c0.n22_adj_2301 ));
    CascadeMux I__4492 (
            .O(N__26329),
            .I(\c0.n9585_cascade_ ));
    InMux I__4491 (
            .O(N__26326),
            .I(N__26323));
    LocalMux I__4490 (
            .O(N__26323),
            .I(N__26319));
    InMux I__4489 (
            .O(N__26322),
            .I(N__26316));
    Sp12to4 I__4488 (
            .O(N__26319),
            .I(N__26313));
    LocalMux I__4487 (
            .O(N__26316),
            .I(data_in_frame_7_1));
    Odrv12 I__4486 (
            .O(N__26313),
            .I(data_in_frame_7_1));
    CascadeMux I__4485 (
            .O(N__26308),
            .I(N__26305));
    InMux I__4484 (
            .O(N__26305),
            .I(N__26301));
    InMux I__4483 (
            .O(N__26304),
            .I(N__26298));
    LocalMux I__4482 (
            .O(N__26301),
            .I(N__26295));
    LocalMux I__4481 (
            .O(N__26298),
            .I(N__26290));
    Span4Mux_v I__4480 (
            .O(N__26295),
            .I(N__26290));
    Odrv4 I__4479 (
            .O(N__26290),
            .I(data_in_frame_7_4));
    InMux I__4478 (
            .O(N__26287),
            .I(N__26283));
    InMux I__4477 (
            .O(N__26286),
            .I(N__26280));
    LocalMux I__4476 (
            .O(N__26283),
            .I(N__26277));
    LocalMux I__4475 (
            .O(N__26280),
            .I(\c0.data_in_frame_2_5 ));
    Odrv12 I__4474 (
            .O(N__26277),
            .I(\c0.data_in_frame_2_5 ));
    InMux I__4473 (
            .O(N__26272),
            .I(N__26268));
    InMux I__4472 (
            .O(N__26271),
            .I(N__26265));
    LocalMux I__4471 (
            .O(N__26268),
            .I(N__26262));
    LocalMux I__4470 (
            .O(N__26265),
            .I(\c0.data_in_frame_2_3 ));
    Odrv4 I__4469 (
            .O(N__26262),
            .I(\c0.data_in_frame_2_3 ));
    CascadeMux I__4468 (
            .O(N__26257),
            .I(\c0.n2336_cascade_ ));
    InMux I__4467 (
            .O(N__26254),
            .I(N__26250));
    InMux I__4466 (
            .O(N__26253),
            .I(N__26246));
    LocalMux I__4465 (
            .O(N__26250),
            .I(N__26243));
    InMux I__4464 (
            .O(N__26249),
            .I(N__26238));
    LocalMux I__4463 (
            .O(N__26246),
            .I(N__26235));
    Span4Mux_h I__4462 (
            .O(N__26243),
            .I(N__26232));
    InMux I__4461 (
            .O(N__26242),
            .I(N__26229));
    InMux I__4460 (
            .O(N__26241),
            .I(N__26226));
    LocalMux I__4459 (
            .O(N__26238),
            .I(\c0.data_in_frame_1_5 ));
    Odrv4 I__4458 (
            .O(N__26235),
            .I(\c0.data_in_frame_1_5 ));
    Odrv4 I__4457 (
            .O(N__26232),
            .I(\c0.data_in_frame_1_5 ));
    LocalMux I__4456 (
            .O(N__26229),
            .I(\c0.data_in_frame_1_5 ));
    LocalMux I__4455 (
            .O(N__26226),
            .I(\c0.data_in_frame_1_5 ));
    CascadeMux I__4454 (
            .O(N__26215),
            .I(\c0.n20_adj_2340_cascade_ ));
    InMux I__4453 (
            .O(N__26212),
            .I(N__26209));
    LocalMux I__4452 (
            .O(N__26209),
            .I(N__26204));
    InMux I__4451 (
            .O(N__26208),
            .I(N__26200));
    CascadeMux I__4450 (
            .O(N__26207),
            .I(N__26197));
    Span4Mux_h I__4449 (
            .O(N__26204),
            .I(N__26194));
    InMux I__4448 (
            .O(N__26203),
            .I(N__26191));
    LocalMux I__4447 (
            .O(N__26200),
            .I(N__26188));
    InMux I__4446 (
            .O(N__26197),
            .I(N__26185));
    Odrv4 I__4445 (
            .O(N__26194),
            .I(data_in_3_2));
    LocalMux I__4444 (
            .O(N__26191),
            .I(data_in_3_2));
    Odrv4 I__4443 (
            .O(N__26188),
            .I(data_in_3_2));
    LocalMux I__4442 (
            .O(N__26185),
            .I(data_in_3_2));
    InMux I__4441 (
            .O(N__26176),
            .I(N__26170));
    InMux I__4440 (
            .O(N__26175),
            .I(N__26165));
    InMux I__4439 (
            .O(N__26174),
            .I(N__26165));
    InMux I__4438 (
            .O(N__26173),
            .I(N__26162));
    LocalMux I__4437 (
            .O(N__26170),
            .I(N__26159));
    LocalMux I__4436 (
            .O(N__26165),
            .I(data_in_2_2));
    LocalMux I__4435 (
            .O(N__26162),
            .I(data_in_2_2));
    Odrv4 I__4434 (
            .O(N__26159),
            .I(data_in_2_2));
    InMux I__4433 (
            .O(N__26152),
            .I(N__26145));
    InMux I__4432 (
            .O(N__26151),
            .I(N__26145));
    InMux I__4431 (
            .O(N__26150),
            .I(N__26141));
    LocalMux I__4430 (
            .O(N__26145),
            .I(N__26138));
    InMux I__4429 (
            .O(N__26144),
            .I(N__26135));
    LocalMux I__4428 (
            .O(N__26141),
            .I(N__26132));
    Span4Mux_h I__4427 (
            .O(N__26138),
            .I(N__26126));
    LocalMux I__4426 (
            .O(N__26135),
            .I(N__26126));
    Span4Mux_h I__4425 (
            .O(N__26132),
            .I(N__26123));
    InMux I__4424 (
            .O(N__26131),
            .I(N__26120));
    Sp12to4 I__4423 (
            .O(N__26126),
            .I(N__26117));
    Odrv4 I__4422 (
            .O(N__26123),
            .I(data_in_1_2));
    LocalMux I__4421 (
            .O(N__26120),
            .I(data_in_1_2));
    Odrv12 I__4420 (
            .O(N__26117),
            .I(data_in_1_2));
    CascadeMux I__4419 (
            .O(N__26110),
            .I(N__26106));
    CascadeMux I__4418 (
            .O(N__26109),
            .I(N__26103));
    InMux I__4417 (
            .O(N__26106),
            .I(N__26100));
    InMux I__4416 (
            .O(N__26103),
            .I(N__26097));
    LocalMux I__4415 (
            .O(N__26100),
            .I(\c0.data_in_frame_10_3 ));
    LocalMux I__4414 (
            .O(N__26097),
            .I(\c0.data_in_frame_10_3 ));
    InMux I__4413 (
            .O(N__26092),
            .I(N__26088));
    InMux I__4412 (
            .O(N__26091),
            .I(N__26085));
    LocalMux I__4411 (
            .O(N__26088),
            .I(N__26082));
    LocalMux I__4410 (
            .O(N__26085),
            .I(data_in_frame_6_6));
    Odrv4 I__4409 (
            .O(N__26082),
            .I(data_in_frame_6_6));
    CascadeMux I__4408 (
            .O(N__26077),
            .I(N__26074));
    InMux I__4407 (
            .O(N__26074),
            .I(N__26071));
    LocalMux I__4406 (
            .O(N__26071),
            .I(N__26067));
    InMux I__4405 (
            .O(N__26070),
            .I(N__26064));
    Span4Mux_h I__4404 (
            .O(N__26067),
            .I(N__26061));
    LocalMux I__4403 (
            .O(N__26064),
            .I(data_in_frame_7_7));
    Odrv4 I__4402 (
            .O(N__26061),
            .I(data_in_frame_7_7));
    CascadeMux I__4401 (
            .O(N__26056),
            .I(\c0.n2351_cascade_ ));
    InMux I__4400 (
            .O(N__26053),
            .I(N__26050));
    LocalMux I__4399 (
            .O(N__26050),
            .I(N__26046));
    InMux I__4398 (
            .O(N__26049),
            .I(N__26043));
    Span4Mux_v I__4397 (
            .O(N__26046),
            .I(N__26040));
    LocalMux I__4396 (
            .O(N__26043),
            .I(data_in_frame_6_7));
    Odrv4 I__4395 (
            .O(N__26040),
            .I(data_in_frame_6_7));
    InMux I__4394 (
            .O(N__26035),
            .I(N__26031));
    InMux I__4393 (
            .O(N__26034),
            .I(N__26028));
    LocalMux I__4392 (
            .O(N__26031),
            .I(data_in_frame_6_1));
    LocalMux I__4391 (
            .O(N__26028),
            .I(data_in_frame_6_1));
    CascadeMux I__4390 (
            .O(N__26023),
            .I(\c0.n2352_cascade_ ));
    InMux I__4389 (
            .O(N__26020),
            .I(N__26017));
    LocalMux I__4388 (
            .O(N__26017),
            .I(N__26013));
    InMux I__4387 (
            .O(N__26016),
            .I(N__26010));
    Span4Mux_h I__4386 (
            .O(N__26013),
            .I(N__26007));
    LocalMux I__4385 (
            .O(N__26010),
            .I(data_in_frame_6_3));
    Odrv4 I__4384 (
            .O(N__26007),
            .I(data_in_frame_6_3));
    CascadeMux I__4383 (
            .O(N__26002),
            .I(N__25999));
    InMux I__4382 (
            .O(N__25999),
            .I(N__25996));
    LocalMux I__4381 (
            .O(N__25996),
            .I(N__25993));
    Span4Mux_v I__4380 (
            .O(N__25993),
            .I(N__25989));
    InMux I__4379 (
            .O(N__25992),
            .I(N__25986));
    Span4Mux_h I__4378 (
            .O(N__25989),
            .I(N__25983));
    LocalMux I__4377 (
            .O(N__25986),
            .I(data_in_frame_6_4));
    Odrv4 I__4376 (
            .O(N__25983),
            .I(data_in_frame_6_4));
    InMux I__4375 (
            .O(N__25978),
            .I(N__25975));
    LocalMux I__4374 (
            .O(N__25975),
            .I(\c0.n23_adj_2145 ));
    CascadeMux I__4373 (
            .O(N__25972),
            .I(\c0.n9541_cascade_ ));
    InMux I__4372 (
            .O(N__25969),
            .I(N__25966));
    LocalMux I__4371 (
            .O(N__25966),
            .I(N__25963));
    Span4Mux_h I__4370 (
            .O(N__25963),
            .I(N__25959));
    InMux I__4369 (
            .O(N__25962),
            .I(N__25956));
    Odrv4 I__4368 (
            .O(N__25959),
            .I(\c0.n16943 ));
    LocalMux I__4367 (
            .O(N__25956),
            .I(\c0.n16943 ));
    InMux I__4366 (
            .O(N__25951),
            .I(N__25945));
    InMux I__4365 (
            .O(N__25950),
            .I(N__25942));
    InMux I__4364 (
            .O(N__25949),
            .I(N__25937));
    InMux I__4363 (
            .O(N__25948),
            .I(N__25937));
    LocalMux I__4362 (
            .O(N__25945),
            .I(data_in_frame_0_2));
    LocalMux I__4361 (
            .O(N__25942),
            .I(data_in_frame_0_2));
    LocalMux I__4360 (
            .O(N__25937),
            .I(data_in_frame_0_2));
    InMux I__4359 (
            .O(N__25930),
            .I(N__25926));
    CascadeMux I__4358 (
            .O(N__25929),
            .I(N__25922));
    LocalMux I__4357 (
            .O(N__25926),
            .I(N__25919));
    InMux I__4356 (
            .O(N__25925),
            .I(N__25914));
    InMux I__4355 (
            .O(N__25922),
            .I(N__25914));
    Span4Mux_v I__4354 (
            .O(N__25919),
            .I(N__25909));
    LocalMux I__4353 (
            .O(N__25914),
            .I(N__25909));
    Span4Mux_h I__4352 (
            .O(N__25909),
            .I(N__25905));
    InMux I__4351 (
            .O(N__25908),
            .I(N__25902));
    Span4Mux_v I__4350 (
            .O(N__25905),
            .I(N__25899));
    LocalMux I__4349 (
            .O(N__25902),
            .I(data_in_3_5));
    Odrv4 I__4348 (
            .O(N__25899),
            .I(data_in_3_5));
    InMux I__4347 (
            .O(N__25894),
            .I(N__25891));
    LocalMux I__4346 (
            .O(N__25891),
            .I(N__25888));
    Span4Mux_v I__4345 (
            .O(N__25888),
            .I(N__25883));
    InMux I__4344 (
            .O(N__25887),
            .I(N__25880));
    CascadeMux I__4343 (
            .O(N__25886),
            .I(N__25876));
    Span4Mux_h I__4342 (
            .O(N__25883),
            .I(N__25871));
    LocalMux I__4341 (
            .O(N__25880),
            .I(N__25871));
    InMux I__4340 (
            .O(N__25879),
            .I(N__25866));
    InMux I__4339 (
            .O(N__25876),
            .I(N__25866));
    Odrv4 I__4338 (
            .O(N__25871),
            .I(data_in_2_5));
    LocalMux I__4337 (
            .O(N__25866),
            .I(data_in_2_5));
    InMux I__4336 (
            .O(N__25861),
            .I(N__25855));
    InMux I__4335 (
            .O(N__25860),
            .I(N__25855));
    LocalMux I__4334 (
            .O(N__25855),
            .I(N__25852));
    Span4Mux_v I__4333 (
            .O(N__25852),
            .I(N__25847));
    InMux I__4332 (
            .O(N__25851),
            .I(N__25842));
    InMux I__4331 (
            .O(N__25850),
            .I(N__25842));
    Odrv4 I__4330 (
            .O(N__25847),
            .I(data_in_2_7));
    LocalMux I__4329 (
            .O(N__25842),
            .I(data_in_2_7));
    InMux I__4328 (
            .O(N__25837),
            .I(N__25834));
    LocalMux I__4327 (
            .O(N__25834),
            .I(N__25831));
    Odrv4 I__4326 (
            .O(N__25831),
            .I(\c0.n8_adj_2157 ));
    CascadeMux I__4325 (
            .O(N__25828),
            .I(N__25825));
    InMux I__4324 (
            .O(N__25825),
            .I(N__25819));
    InMux I__4323 (
            .O(N__25824),
            .I(N__25819));
    LocalMux I__4322 (
            .O(N__25819),
            .I(N__25814));
    InMux I__4321 (
            .O(N__25818),
            .I(N__25809));
    InMux I__4320 (
            .O(N__25817),
            .I(N__25809));
    Span4Mux_h I__4319 (
            .O(N__25814),
            .I(N__25806));
    LocalMux I__4318 (
            .O(N__25809),
            .I(data_in_3_7));
    Odrv4 I__4317 (
            .O(N__25806),
            .I(data_in_3_7));
    InMux I__4316 (
            .O(N__25801),
            .I(N__25798));
    LocalMux I__4315 (
            .O(N__25798),
            .I(N__25795));
    Span4Mux_h I__4314 (
            .O(N__25795),
            .I(N__25791));
    InMux I__4313 (
            .O(N__25794),
            .I(N__25787));
    Span4Mux_h I__4312 (
            .O(N__25791),
            .I(N__25784));
    InMux I__4311 (
            .O(N__25790),
            .I(N__25781));
    LocalMux I__4310 (
            .O(N__25787),
            .I(data_in_3_3));
    Odrv4 I__4309 (
            .O(N__25784),
            .I(data_in_3_3));
    LocalMux I__4308 (
            .O(N__25781),
            .I(data_in_3_3));
    InMux I__4307 (
            .O(N__25774),
            .I(N__25771));
    LocalMux I__4306 (
            .O(N__25771),
            .I(N__25767));
    InMux I__4305 (
            .O(N__25770),
            .I(N__25764));
    Span4Mux_v I__4304 (
            .O(N__25767),
            .I(N__25761));
    LocalMux I__4303 (
            .O(N__25764),
            .I(data_in_frame_7_0));
    Odrv4 I__4302 (
            .O(N__25761),
            .I(data_in_frame_7_0));
    CascadeMux I__4301 (
            .O(N__25756),
            .I(N__25753));
    InMux I__4300 (
            .O(N__25753),
            .I(N__25750));
    LocalMux I__4299 (
            .O(N__25750),
            .I(N__25746));
    InMux I__4298 (
            .O(N__25749),
            .I(N__25743));
    Span4Mux_h I__4297 (
            .O(N__25746),
            .I(N__25740));
    LocalMux I__4296 (
            .O(N__25743),
            .I(data_in_frame_7_6));
    Odrv4 I__4295 (
            .O(N__25740),
            .I(data_in_frame_7_6));
    InMux I__4294 (
            .O(N__25735),
            .I(N__25732));
    LocalMux I__4293 (
            .O(N__25732),
            .I(N__25728));
    InMux I__4292 (
            .O(N__25731),
            .I(N__25725));
    Span4Mux_h I__4291 (
            .O(N__25728),
            .I(N__25719));
    LocalMux I__4290 (
            .O(N__25725),
            .I(N__25719));
    InMux I__4289 (
            .O(N__25724),
            .I(N__25716));
    Span4Mux_v I__4288 (
            .O(N__25719),
            .I(N__25706));
    LocalMux I__4287 (
            .O(N__25716),
            .I(N__25706));
    InMux I__4286 (
            .O(N__25715),
            .I(N__25703));
    InMux I__4285 (
            .O(N__25714),
            .I(N__25700));
    InMux I__4284 (
            .O(N__25713),
            .I(N__25695));
    InMux I__4283 (
            .O(N__25712),
            .I(N__25695));
    InMux I__4282 (
            .O(N__25711),
            .I(N__25692));
    Span4Mux_h I__4281 (
            .O(N__25706),
            .I(N__25689));
    LocalMux I__4280 (
            .O(N__25703),
            .I(N__25680));
    LocalMux I__4279 (
            .O(N__25700),
            .I(N__25680));
    LocalMux I__4278 (
            .O(N__25695),
            .I(N__25680));
    LocalMux I__4277 (
            .O(N__25692),
            .I(N__25680));
    Odrv4 I__4276 (
            .O(N__25689),
            .I(n16896));
    Odrv12 I__4275 (
            .O(N__25680),
            .I(n16896));
    CascadeMux I__4274 (
            .O(N__25675),
            .I(N__25669));
    CascadeMux I__4273 (
            .O(N__25674),
            .I(N__25666));
    InMux I__4272 (
            .O(N__25673),
            .I(N__25661));
    InMux I__4271 (
            .O(N__25672),
            .I(N__25658));
    InMux I__4270 (
            .O(N__25669),
            .I(N__25653));
    InMux I__4269 (
            .O(N__25666),
            .I(N__25653));
    CascadeMux I__4268 (
            .O(N__25665),
            .I(N__25650));
    InMux I__4267 (
            .O(N__25664),
            .I(N__25646));
    LocalMux I__4266 (
            .O(N__25661),
            .I(N__25643));
    LocalMux I__4265 (
            .O(N__25658),
            .I(N__25640));
    LocalMux I__4264 (
            .O(N__25653),
            .I(N__25635));
    InMux I__4263 (
            .O(N__25650),
            .I(N__25630));
    InMux I__4262 (
            .O(N__25649),
            .I(N__25630));
    LocalMux I__4261 (
            .O(N__25646),
            .I(N__25627));
    Span4Mux_h I__4260 (
            .O(N__25643),
            .I(N__25622));
    Span4Mux_h I__4259 (
            .O(N__25640),
            .I(N__25622));
    InMux I__4258 (
            .O(N__25639),
            .I(N__25619));
    InMux I__4257 (
            .O(N__25638),
            .I(N__25616));
    Odrv4 I__4256 (
            .O(N__25635),
            .I(rx_data_6));
    LocalMux I__4255 (
            .O(N__25630),
            .I(rx_data_6));
    Odrv4 I__4254 (
            .O(N__25627),
            .I(rx_data_6));
    Odrv4 I__4253 (
            .O(N__25622),
            .I(rx_data_6));
    LocalMux I__4252 (
            .O(N__25619),
            .I(rx_data_6));
    LocalMux I__4251 (
            .O(N__25616),
            .I(rx_data_6));
    InMux I__4250 (
            .O(N__25603),
            .I(N__25599));
    InMux I__4249 (
            .O(N__25602),
            .I(N__25596));
    LocalMux I__4248 (
            .O(N__25599),
            .I(N__25590));
    LocalMux I__4247 (
            .O(N__25596),
            .I(N__25586));
    CascadeMux I__4246 (
            .O(N__25595),
            .I(N__25582));
    InMux I__4245 (
            .O(N__25594),
            .I(N__25579));
    CascadeMux I__4244 (
            .O(N__25593),
            .I(N__25576));
    Sp12to4 I__4243 (
            .O(N__25590),
            .I(N__25573));
    CascadeMux I__4242 (
            .O(N__25589),
            .I(N__25570));
    Span4Mux_v I__4241 (
            .O(N__25586),
            .I(N__25567));
    InMux I__4240 (
            .O(N__25585),
            .I(N__25564));
    InMux I__4239 (
            .O(N__25582),
            .I(N__25559));
    LocalMux I__4238 (
            .O(N__25579),
            .I(N__25556));
    InMux I__4237 (
            .O(N__25576),
            .I(N__25553));
    Span12Mux_v I__4236 (
            .O(N__25573),
            .I(N__25550));
    InMux I__4235 (
            .O(N__25570),
            .I(N__25547));
    Span4Mux_s1_h I__4234 (
            .O(N__25567),
            .I(N__25542));
    LocalMux I__4233 (
            .O(N__25564),
            .I(N__25542));
    InMux I__4232 (
            .O(N__25563),
            .I(N__25539));
    InMux I__4231 (
            .O(N__25562),
            .I(N__25536));
    LocalMux I__4230 (
            .O(N__25559),
            .I(rx_data_0));
    Odrv4 I__4229 (
            .O(N__25556),
            .I(rx_data_0));
    LocalMux I__4228 (
            .O(N__25553),
            .I(rx_data_0));
    Odrv12 I__4227 (
            .O(N__25550),
            .I(rx_data_0));
    LocalMux I__4226 (
            .O(N__25547),
            .I(rx_data_0));
    Odrv4 I__4225 (
            .O(N__25542),
            .I(rx_data_0));
    LocalMux I__4224 (
            .O(N__25539),
            .I(rx_data_0));
    LocalMux I__4223 (
            .O(N__25536),
            .I(rx_data_0));
    InMux I__4222 (
            .O(N__25519),
            .I(N__25516));
    LocalMux I__4221 (
            .O(N__25516),
            .I(N__25510));
    InMux I__4220 (
            .O(N__25515),
            .I(N__25503));
    InMux I__4219 (
            .O(N__25514),
            .I(N__25503));
    InMux I__4218 (
            .O(N__25513),
            .I(N__25503));
    Odrv12 I__4217 (
            .O(N__25510),
            .I(\c0.FRAME_MATCHER_state_22 ));
    LocalMux I__4216 (
            .O(N__25503),
            .I(\c0.FRAME_MATCHER_state_22 ));
    SRMux I__4215 (
            .O(N__25498),
            .I(N__25495));
    LocalMux I__4214 (
            .O(N__25495),
            .I(N__25492));
    Span4Mux_v I__4213 (
            .O(N__25492),
            .I(N__25489));
    Odrv4 I__4212 (
            .O(N__25489),
            .I(\c0.n16365 ));
    InMux I__4211 (
            .O(N__25486),
            .I(N__25483));
    LocalMux I__4210 (
            .O(N__25483),
            .I(N__25480));
    Odrv4 I__4209 (
            .O(N__25480),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_12 ));
    CascadeMux I__4208 (
            .O(N__25477),
            .I(N__25474));
    InMux I__4207 (
            .O(N__25474),
            .I(N__25471));
    LocalMux I__4206 (
            .O(N__25471),
            .I(N__25466));
    InMux I__4205 (
            .O(N__25470),
            .I(N__25463));
    InMux I__4204 (
            .O(N__25469),
            .I(N__25460));
    Span4Mux_v I__4203 (
            .O(N__25466),
            .I(N__25455));
    LocalMux I__4202 (
            .O(N__25463),
            .I(N__25455));
    LocalMux I__4201 (
            .O(N__25460),
            .I(N__25452));
    Span4Mux_h I__4200 (
            .O(N__25455),
            .I(N__25446));
    Span4Mux_h I__4199 (
            .O(N__25452),
            .I(N__25446));
    InMux I__4198 (
            .O(N__25451),
            .I(N__25443));
    Odrv4 I__4197 (
            .O(N__25446),
            .I(\c0.FRAME_MATCHER_i_12 ));
    LocalMux I__4196 (
            .O(N__25443),
            .I(\c0.FRAME_MATCHER_i_12 ));
    SRMux I__4195 (
            .O(N__25438),
            .I(N__25435));
    LocalMux I__4194 (
            .O(N__25435),
            .I(N__25432));
    Span4Mux_h I__4193 (
            .O(N__25432),
            .I(N__25429));
    Odrv4 I__4192 (
            .O(N__25429),
            .I(\c0.n3_adj_2245 ));
    SRMux I__4191 (
            .O(N__25426),
            .I(N__25423));
    LocalMux I__4190 (
            .O(N__25423),
            .I(N__25420));
    Span4Mux_v I__4189 (
            .O(N__25420),
            .I(N__25417));
    Odrv4 I__4188 (
            .O(N__25417),
            .I(\c0.n16351 ));
    InMux I__4187 (
            .O(N__25414),
            .I(N__25409));
    CascadeMux I__4186 (
            .O(N__25413),
            .I(N__25405));
    InMux I__4185 (
            .O(N__25412),
            .I(N__25402));
    LocalMux I__4184 (
            .O(N__25409),
            .I(N__25399));
    InMux I__4183 (
            .O(N__25408),
            .I(N__25394));
    InMux I__4182 (
            .O(N__25405),
            .I(N__25394));
    LocalMux I__4181 (
            .O(N__25402),
            .I(\c0.FRAME_MATCHER_state_21 ));
    Odrv12 I__4180 (
            .O(N__25399),
            .I(\c0.FRAME_MATCHER_state_21 ));
    LocalMux I__4179 (
            .O(N__25394),
            .I(\c0.FRAME_MATCHER_state_21 ));
    SRMux I__4178 (
            .O(N__25387),
            .I(N__25384));
    LocalMux I__4177 (
            .O(N__25384),
            .I(N__25381));
    Span4Mux_v I__4176 (
            .O(N__25381),
            .I(N__25378));
    Odrv4 I__4175 (
            .O(N__25378),
            .I(\c0.n16367 ));
    InMux I__4174 (
            .O(N__25375),
            .I(N__25370));
    InMux I__4173 (
            .O(N__25374),
            .I(N__25367));
    InMux I__4172 (
            .O(N__25373),
            .I(N__25363));
    LocalMux I__4171 (
            .O(N__25370),
            .I(N__25360));
    LocalMux I__4170 (
            .O(N__25367),
            .I(N__25357));
    InMux I__4169 (
            .O(N__25366),
            .I(N__25354));
    LocalMux I__4168 (
            .O(N__25363),
            .I(\c0.FRAME_MATCHER_state_26 ));
    Odrv12 I__4167 (
            .O(N__25360),
            .I(\c0.FRAME_MATCHER_state_26 ));
    Odrv4 I__4166 (
            .O(N__25357),
            .I(\c0.FRAME_MATCHER_state_26 ));
    LocalMux I__4165 (
            .O(N__25354),
            .I(\c0.FRAME_MATCHER_state_26 ));
    SRMux I__4164 (
            .O(N__25345),
            .I(N__25342));
    LocalMux I__4163 (
            .O(N__25342),
            .I(N__25339));
    Span4Mux_v I__4162 (
            .O(N__25339),
            .I(N__25336));
    Odrv4 I__4161 (
            .O(N__25336),
            .I(\c0.n16357 ));
    InMux I__4160 (
            .O(N__25333),
            .I(N__25330));
    LocalMux I__4159 (
            .O(N__25330),
            .I(N__25325));
    InMux I__4158 (
            .O(N__25329),
            .I(N__25322));
    InMux I__4157 (
            .O(N__25328),
            .I(N__25319));
    Span4Mux_v I__4156 (
            .O(N__25325),
            .I(N__25314));
    LocalMux I__4155 (
            .O(N__25322),
            .I(N__25314));
    LocalMux I__4154 (
            .O(N__25319),
            .I(\c0.FRAME_MATCHER_state_27 ));
    Odrv4 I__4153 (
            .O(N__25314),
            .I(\c0.FRAME_MATCHER_state_27 ));
    SRMux I__4152 (
            .O(N__25309),
            .I(N__25306));
    LocalMux I__4151 (
            .O(N__25306),
            .I(N__25303));
    Span4Mux_s3_h I__4150 (
            .O(N__25303),
            .I(N__25300));
    Span4Mux_h I__4149 (
            .O(N__25300),
            .I(N__25297));
    Odrv4 I__4148 (
            .O(N__25297),
            .I(\c0.n16355 ));
    CascadeMux I__4147 (
            .O(N__25294),
            .I(N__25289));
    InMux I__4146 (
            .O(N__25293),
            .I(N__25286));
    InMux I__4145 (
            .O(N__25292),
            .I(N__25283));
    InMux I__4144 (
            .O(N__25289),
            .I(N__25280));
    LocalMux I__4143 (
            .O(N__25286),
            .I(N__25277));
    LocalMux I__4142 (
            .O(N__25283),
            .I(data_in_0_1));
    LocalMux I__4141 (
            .O(N__25280),
            .I(data_in_0_1));
    Odrv4 I__4140 (
            .O(N__25277),
            .I(data_in_0_1));
    InMux I__4139 (
            .O(N__25270),
            .I(N__25267));
    LocalMux I__4138 (
            .O(N__25267),
            .I(N__25264));
    Odrv4 I__4137 (
            .O(N__25264),
            .I(\c0.n17266 ));
    InMux I__4136 (
            .O(N__25261),
            .I(N__25256));
    InMux I__4135 (
            .O(N__25260),
            .I(N__25253));
    InMux I__4134 (
            .O(N__25259),
            .I(N__25250));
    LocalMux I__4133 (
            .O(N__25256),
            .I(N__25247));
    LocalMux I__4132 (
            .O(N__25253),
            .I(\c0.FRAME_MATCHER_state_10 ));
    LocalMux I__4131 (
            .O(N__25250),
            .I(\c0.FRAME_MATCHER_state_10 ));
    Odrv12 I__4130 (
            .O(N__25247),
            .I(\c0.FRAME_MATCHER_state_10 ));
    InMux I__4129 (
            .O(N__25240),
            .I(N__25237));
    LocalMux I__4128 (
            .O(N__25237),
            .I(N__25234));
    Odrv4 I__4127 (
            .O(N__25234),
            .I(\c0.n6_adj_2213 ));
    InMux I__4126 (
            .O(N__25231),
            .I(N__25228));
    LocalMux I__4125 (
            .O(N__25228),
            .I(\c0.n16869 ));
    CascadeMux I__4124 (
            .O(N__25225),
            .I(\c0.n16869_cascade_ ));
    CascadeMux I__4123 (
            .O(N__25222),
            .I(\c0.n16871_cascade_ ));
    InMux I__4122 (
            .O(N__25219),
            .I(N__25216));
    LocalMux I__4121 (
            .O(N__25216),
            .I(\c0.n16876 ));
    CascadeMux I__4120 (
            .O(N__25213),
            .I(N__25210));
    InMux I__4119 (
            .O(N__25210),
            .I(N__25207));
    LocalMux I__4118 (
            .O(N__25207),
            .I(\c0.n50 ));
    InMux I__4117 (
            .O(N__25204),
            .I(N__25201));
    LocalMux I__4116 (
            .O(N__25201),
            .I(N__25198));
    Span4Mux_h I__4115 (
            .O(N__25198),
            .I(N__25195));
    Span4Mux_v I__4114 (
            .O(N__25195),
            .I(N__25192));
    Odrv4 I__4113 (
            .O(N__25192),
            .I(\c0.n46 ));
    CascadeMux I__4112 (
            .O(N__25189),
            .I(\c0.n56_adj_2146_cascade_ ));
    InMux I__4111 (
            .O(N__25186),
            .I(N__25183));
    LocalMux I__4110 (
            .O(N__25183),
            .I(\c0.n51 ));
    InMux I__4109 (
            .O(N__25180),
            .I(N__25176));
    InMux I__4108 (
            .O(N__25179),
            .I(N__25172));
    LocalMux I__4107 (
            .O(N__25176),
            .I(N__25169));
    InMux I__4106 (
            .O(N__25175),
            .I(N__25165));
    LocalMux I__4105 (
            .O(N__25172),
            .I(N__25160));
    Span4Mux_v I__4104 (
            .O(N__25169),
            .I(N__25160));
    InMux I__4103 (
            .O(N__25168),
            .I(N__25157));
    LocalMux I__4102 (
            .O(N__25165),
            .I(N__25154));
    Span4Mux_v I__4101 (
            .O(N__25160),
            .I(N__25151));
    LocalMux I__4100 (
            .O(N__25157),
            .I(\c0.n9346 ));
    Odrv4 I__4099 (
            .O(N__25154),
            .I(\c0.n9346 ));
    Odrv4 I__4098 (
            .O(N__25151),
            .I(\c0.n9346 ));
    CascadeMux I__4097 (
            .O(N__25144),
            .I(N__25141));
    InMux I__4096 (
            .O(N__25141),
            .I(N__25137));
    CascadeMux I__4095 (
            .O(N__25140),
            .I(N__25134));
    LocalMux I__4094 (
            .O(N__25137),
            .I(N__25131));
    InMux I__4093 (
            .O(N__25134),
            .I(N__25128));
    Span4Mux_v I__4092 (
            .O(N__25131),
            .I(N__25123));
    LocalMux I__4091 (
            .O(N__25128),
            .I(N__25123));
    Span4Mux_h I__4090 (
            .O(N__25123),
            .I(N__25117));
    InMux I__4089 (
            .O(N__25122),
            .I(N__25113));
    InMux I__4088 (
            .O(N__25121),
            .I(N__25110));
    InMux I__4087 (
            .O(N__25120),
            .I(N__25107));
    Span4Mux_v I__4086 (
            .O(N__25117),
            .I(N__25104));
    InMux I__4085 (
            .O(N__25116),
            .I(N__25101));
    LocalMux I__4084 (
            .O(N__25113),
            .I(N__25096));
    LocalMux I__4083 (
            .O(N__25110),
            .I(N__25096));
    LocalMux I__4082 (
            .O(N__25107),
            .I(\c0.FRAME_MATCHER_i_3 ));
    Odrv4 I__4081 (
            .O(N__25104),
            .I(\c0.FRAME_MATCHER_i_3 ));
    LocalMux I__4080 (
            .O(N__25101),
            .I(\c0.FRAME_MATCHER_i_3 ));
    Odrv12 I__4079 (
            .O(N__25096),
            .I(\c0.FRAME_MATCHER_i_3 ));
    InMux I__4078 (
            .O(N__25087),
            .I(N__25081));
    InMux I__4077 (
            .O(N__25086),
            .I(N__25077));
    InMux I__4076 (
            .O(N__25085),
            .I(N__25074));
    InMux I__4075 (
            .O(N__25084),
            .I(N__25070));
    LocalMux I__4074 (
            .O(N__25081),
            .I(N__25067));
    CascadeMux I__4073 (
            .O(N__25080),
            .I(N__25063));
    LocalMux I__4072 (
            .O(N__25077),
            .I(N__25057));
    LocalMux I__4071 (
            .O(N__25074),
            .I(N__25057));
    CascadeMux I__4070 (
            .O(N__25073),
            .I(N__25054));
    LocalMux I__4069 (
            .O(N__25070),
            .I(N__25051));
    Span4Mux_v I__4068 (
            .O(N__25067),
            .I(N__25048));
    InMux I__4067 (
            .O(N__25066),
            .I(N__25045));
    InMux I__4066 (
            .O(N__25063),
            .I(N__25040));
    InMux I__4065 (
            .O(N__25062),
            .I(N__25040));
    Span4Mux_v I__4064 (
            .O(N__25057),
            .I(N__25037));
    InMux I__4063 (
            .O(N__25054),
            .I(N__25034));
    Span4Mux_v I__4062 (
            .O(N__25051),
            .I(N__25029));
    Span4Mux_h I__4061 (
            .O(N__25048),
            .I(N__25029));
    LocalMux I__4060 (
            .O(N__25045),
            .I(\c0.FRAME_MATCHER_i_2 ));
    LocalMux I__4059 (
            .O(N__25040),
            .I(\c0.FRAME_MATCHER_i_2 ));
    Odrv4 I__4058 (
            .O(N__25037),
            .I(\c0.FRAME_MATCHER_i_2 ));
    LocalMux I__4057 (
            .O(N__25034),
            .I(\c0.FRAME_MATCHER_i_2 ));
    Odrv4 I__4056 (
            .O(N__25029),
            .I(\c0.FRAME_MATCHER_i_2 ));
    CascadeMux I__4055 (
            .O(N__25018),
            .I(N__25013));
    InMux I__4054 (
            .O(N__25017),
            .I(N__25010));
    CascadeMux I__4053 (
            .O(N__25016),
            .I(N__25007));
    InMux I__4052 (
            .O(N__25013),
            .I(N__25004));
    LocalMux I__4051 (
            .O(N__25010),
            .I(N__25001));
    InMux I__4050 (
            .O(N__25007),
            .I(N__24998));
    LocalMux I__4049 (
            .O(N__25004),
            .I(N__24994));
    Span4Mux_v I__4048 (
            .O(N__25001),
            .I(N__24989));
    LocalMux I__4047 (
            .O(N__24998),
            .I(N__24989));
    InMux I__4046 (
            .O(N__24997),
            .I(N__24986));
    Span4Mux_v I__4045 (
            .O(N__24994),
            .I(N__24983));
    Span4Mux_h I__4044 (
            .O(N__24989),
            .I(N__24980));
    LocalMux I__4043 (
            .O(N__24986),
            .I(N__24975));
    Span4Mux_v I__4042 (
            .O(N__24983),
            .I(N__24975));
    Span4Mux_v I__4041 (
            .O(N__24980),
            .I(N__24972));
    Odrv4 I__4040 (
            .O(N__24975),
            .I(\c0.FRAME_MATCHER_i_28 ));
    Odrv4 I__4039 (
            .O(N__24972),
            .I(\c0.FRAME_MATCHER_i_28 ));
    InMux I__4038 (
            .O(N__24967),
            .I(N__24964));
    LocalMux I__4037 (
            .O(N__24964),
            .I(\c0.n45 ));
    CascadeMux I__4036 (
            .O(N__24961),
            .I(N__24957));
    InMux I__4035 (
            .O(N__24960),
            .I(N__24952));
    InMux I__4034 (
            .O(N__24957),
            .I(N__24949));
    InMux I__4033 (
            .O(N__24956),
            .I(N__24946));
    InMux I__4032 (
            .O(N__24955),
            .I(N__24943));
    LocalMux I__4031 (
            .O(N__24952),
            .I(N__24940));
    LocalMux I__4030 (
            .O(N__24949),
            .I(N__24937));
    LocalMux I__4029 (
            .O(N__24946),
            .I(N__24934));
    LocalMux I__4028 (
            .O(N__24943),
            .I(N__24931));
    Span4Mux_v I__4027 (
            .O(N__24940),
            .I(N__24924));
    Span4Mux_v I__4026 (
            .O(N__24937),
            .I(N__24924));
    Span4Mux_h I__4025 (
            .O(N__24934),
            .I(N__24924));
    Span4Mux_v I__4024 (
            .O(N__24931),
            .I(N__24921));
    Span4Mux_h I__4023 (
            .O(N__24924),
            .I(N__24918));
    Odrv4 I__4022 (
            .O(N__24921),
            .I(\c0.FRAME_MATCHER_i_27 ));
    Odrv4 I__4021 (
            .O(N__24918),
            .I(\c0.FRAME_MATCHER_i_27 ));
    CascadeMux I__4020 (
            .O(N__24913),
            .I(N__24910));
    InMux I__4019 (
            .O(N__24910),
            .I(N__24904));
    InMux I__4018 (
            .O(N__24909),
            .I(N__24901));
    CascadeMux I__4017 (
            .O(N__24908),
            .I(N__24898));
    InMux I__4016 (
            .O(N__24907),
            .I(N__24895));
    LocalMux I__4015 (
            .O(N__24904),
            .I(N__24892));
    LocalMux I__4014 (
            .O(N__24901),
            .I(N__24889));
    InMux I__4013 (
            .O(N__24898),
            .I(N__24886));
    LocalMux I__4012 (
            .O(N__24895),
            .I(N__24883));
    Span4Mux_v I__4011 (
            .O(N__24892),
            .I(N__24880));
    Span4Mux_v I__4010 (
            .O(N__24889),
            .I(N__24877));
    LocalMux I__4009 (
            .O(N__24886),
            .I(\c0.FRAME_MATCHER_i_30 ));
    Odrv12 I__4008 (
            .O(N__24883),
            .I(\c0.FRAME_MATCHER_i_30 ));
    Odrv4 I__4007 (
            .O(N__24880),
            .I(\c0.FRAME_MATCHER_i_30 ));
    Odrv4 I__4006 (
            .O(N__24877),
            .I(\c0.FRAME_MATCHER_i_30 ));
    CascadeMux I__4005 (
            .O(N__24868),
            .I(N__24865));
    InMux I__4004 (
            .O(N__24865),
            .I(N__24861));
    CascadeMux I__4003 (
            .O(N__24864),
            .I(N__24857));
    LocalMux I__4002 (
            .O(N__24861),
            .I(N__24854));
    InMux I__4001 (
            .O(N__24860),
            .I(N__24851));
    InMux I__4000 (
            .O(N__24857),
            .I(N__24848));
    Span4Mux_v I__3999 (
            .O(N__24854),
            .I(N__24840));
    LocalMux I__3998 (
            .O(N__24851),
            .I(N__24840));
    LocalMux I__3997 (
            .O(N__24848),
            .I(N__24840));
    InMux I__3996 (
            .O(N__24847),
            .I(N__24837));
    Span4Mux_h I__3995 (
            .O(N__24840),
            .I(N__24834));
    LocalMux I__3994 (
            .O(N__24837),
            .I(N__24831));
    Span4Mux_h I__3993 (
            .O(N__24834),
            .I(N__24828));
    Odrv4 I__3992 (
            .O(N__24831),
            .I(\c0.FRAME_MATCHER_i_8 ));
    Odrv4 I__3991 (
            .O(N__24828),
            .I(\c0.FRAME_MATCHER_i_8 ));
    CascadeMux I__3990 (
            .O(N__24823),
            .I(N__24819));
    CascadeMux I__3989 (
            .O(N__24822),
            .I(N__24815));
    InMux I__3988 (
            .O(N__24819),
            .I(N__24812));
    InMux I__3987 (
            .O(N__24818),
            .I(N__24809));
    InMux I__3986 (
            .O(N__24815),
            .I(N__24805));
    LocalMux I__3985 (
            .O(N__24812),
            .I(N__24800));
    LocalMux I__3984 (
            .O(N__24809),
            .I(N__24800));
    InMux I__3983 (
            .O(N__24808),
            .I(N__24797));
    LocalMux I__3982 (
            .O(N__24805),
            .I(N__24794));
    Span4Mux_v I__3981 (
            .O(N__24800),
            .I(N__24789));
    LocalMux I__3980 (
            .O(N__24797),
            .I(N__24789));
    Span4Mux_v I__3979 (
            .O(N__24794),
            .I(N__24784));
    Span4Mux_h I__3978 (
            .O(N__24789),
            .I(N__24784));
    Span4Mux_h I__3977 (
            .O(N__24784),
            .I(N__24781));
    Odrv4 I__3976 (
            .O(N__24781),
            .I(\c0.FRAME_MATCHER_i_26 ));
    InMux I__3975 (
            .O(N__24778),
            .I(N__24775));
    LocalMux I__3974 (
            .O(N__24775),
            .I(\c0.n47_adj_2144 ));
    CascadeMux I__3973 (
            .O(N__24772),
            .I(N__24769));
    InMux I__3972 (
            .O(N__24769),
            .I(N__24765));
    InMux I__3971 (
            .O(N__24768),
            .I(N__24762));
    LocalMux I__3970 (
            .O(N__24765),
            .I(N__24758));
    LocalMux I__3969 (
            .O(N__24762),
            .I(N__24755));
    InMux I__3968 (
            .O(N__24761),
            .I(N__24752));
    Span4Mux_h I__3967 (
            .O(N__24758),
            .I(N__24748));
    Span4Mux_h I__3966 (
            .O(N__24755),
            .I(N__24743));
    LocalMux I__3965 (
            .O(N__24752),
            .I(N__24743));
    InMux I__3964 (
            .O(N__24751),
            .I(N__24740));
    Span4Mux_h I__3963 (
            .O(N__24748),
            .I(N__24735));
    Span4Mux_h I__3962 (
            .O(N__24743),
            .I(N__24735));
    LocalMux I__3961 (
            .O(N__24740),
            .I(N__24732));
    Odrv4 I__3960 (
            .O(N__24735),
            .I(\c0.FRAME_MATCHER_i_22 ));
    Odrv12 I__3959 (
            .O(N__24732),
            .I(\c0.FRAME_MATCHER_i_22 ));
    CascadeMux I__3958 (
            .O(N__24727),
            .I(N__24723));
    CascadeMux I__3957 (
            .O(N__24726),
            .I(N__24719));
    InMux I__3956 (
            .O(N__24723),
            .I(N__24716));
    InMux I__3955 (
            .O(N__24722),
            .I(N__24713));
    InMux I__3954 (
            .O(N__24719),
            .I(N__24709));
    LocalMux I__3953 (
            .O(N__24716),
            .I(N__24704));
    LocalMux I__3952 (
            .O(N__24713),
            .I(N__24704));
    InMux I__3951 (
            .O(N__24712),
            .I(N__24701));
    LocalMux I__3950 (
            .O(N__24709),
            .I(N__24698));
    Span4Mux_v I__3949 (
            .O(N__24704),
            .I(N__24693));
    LocalMux I__3948 (
            .O(N__24701),
            .I(N__24693));
    Span4Mux_v I__3947 (
            .O(N__24698),
            .I(N__24688));
    Span4Mux_h I__3946 (
            .O(N__24693),
            .I(N__24688));
    Span4Mux_h I__3945 (
            .O(N__24688),
            .I(N__24685));
    Odrv4 I__3944 (
            .O(N__24685),
            .I(\c0.FRAME_MATCHER_i_23 ));
    InMux I__3943 (
            .O(N__24682),
            .I(N__24677));
    InMux I__3942 (
            .O(N__24681),
            .I(N__24674));
    InMux I__3941 (
            .O(N__24680),
            .I(N__24671));
    LocalMux I__3940 (
            .O(N__24677),
            .I(N__24668));
    LocalMux I__3939 (
            .O(N__24674),
            .I(N__24664));
    LocalMux I__3938 (
            .O(N__24671),
            .I(N__24661));
    Span4Mux_h I__3937 (
            .O(N__24668),
            .I(N__24658));
    InMux I__3936 (
            .O(N__24667),
            .I(N__24655));
    Span4Mux_h I__3935 (
            .O(N__24664),
            .I(N__24652));
    Odrv4 I__3934 (
            .O(N__24661),
            .I(\c0.FRAME_MATCHER_i_25 ));
    Odrv4 I__3933 (
            .O(N__24658),
            .I(\c0.FRAME_MATCHER_i_25 ));
    LocalMux I__3932 (
            .O(N__24655),
            .I(\c0.FRAME_MATCHER_i_25 ));
    Odrv4 I__3931 (
            .O(N__24652),
            .I(\c0.FRAME_MATCHER_i_25 ));
    InMux I__3930 (
            .O(N__24643),
            .I(N__24640));
    LocalMux I__3929 (
            .O(N__24640),
            .I(\c0.n49 ));
    InMux I__3928 (
            .O(N__24637),
            .I(N__24634));
    LocalMux I__3927 (
            .O(N__24634),
            .I(N__24631));
    Odrv4 I__3926 (
            .O(N__24631),
            .I(\c0.n59 ));
    CascadeMux I__3925 (
            .O(N__24628),
            .I(\c0.n61_cascade_ ));
    InMux I__3924 (
            .O(N__24625),
            .I(N__24622));
    LocalMux I__3923 (
            .O(N__24622),
            .I(\c0.n10_adj_2336 ));
    CascadeMux I__3922 (
            .O(N__24619),
            .I(\c0.n16133_cascade_ ));
    InMux I__3921 (
            .O(N__24616),
            .I(N__24612));
    InMux I__3920 (
            .O(N__24615),
            .I(N__24609));
    LocalMux I__3919 (
            .O(N__24612),
            .I(\c0.n16898 ));
    LocalMux I__3918 (
            .O(N__24609),
            .I(\c0.n16898 ));
    InMux I__3917 (
            .O(N__24604),
            .I(N__24596));
    InMux I__3916 (
            .O(N__24603),
            .I(N__24596));
    InMux I__3915 (
            .O(N__24602),
            .I(N__24593));
    InMux I__3914 (
            .O(N__24601),
            .I(N__24590));
    LocalMux I__3913 (
            .O(N__24596),
            .I(N__24587));
    LocalMux I__3912 (
            .O(N__24593),
            .I(\c0.FRAME_MATCHER_state_19 ));
    LocalMux I__3911 (
            .O(N__24590),
            .I(\c0.FRAME_MATCHER_state_19 ));
    Odrv12 I__3910 (
            .O(N__24587),
            .I(\c0.FRAME_MATCHER_state_19 ));
    InMux I__3909 (
            .O(N__24580),
            .I(N__24577));
    LocalMux I__3908 (
            .O(N__24577),
            .I(\c0.n52 ));
    InMux I__3907 (
            .O(N__24574),
            .I(N__24571));
    LocalMux I__3906 (
            .O(N__24571),
            .I(N__24568));
    Span4Mux_h I__3905 (
            .O(N__24568),
            .I(N__24565));
    Odrv4 I__3904 (
            .O(N__24565),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_4 ));
    SRMux I__3903 (
            .O(N__24562),
            .I(N__24559));
    LocalMux I__3902 (
            .O(N__24559),
            .I(N__24556));
    Span4Mux_h I__3901 (
            .O(N__24556),
            .I(N__24553));
    Odrv4 I__3900 (
            .O(N__24553),
            .I(\c0.n3_adj_2257 ));
    CascadeMux I__3899 (
            .O(N__24550),
            .I(N__24547));
    InMux I__3898 (
            .O(N__24547),
            .I(N__24542));
    InMux I__3897 (
            .O(N__24546),
            .I(N__24539));
    CascadeMux I__3896 (
            .O(N__24545),
            .I(N__24536));
    LocalMux I__3895 (
            .O(N__24542),
            .I(N__24530));
    LocalMux I__3894 (
            .O(N__24539),
            .I(N__24530));
    InMux I__3893 (
            .O(N__24536),
            .I(N__24527));
    InMux I__3892 (
            .O(N__24535),
            .I(N__24524));
    Span4Mux_v I__3891 (
            .O(N__24530),
            .I(N__24521));
    LocalMux I__3890 (
            .O(N__24527),
            .I(N__24516));
    LocalMux I__3889 (
            .O(N__24524),
            .I(N__24516));
    Odrv4 I__3888 (
            .O(N__24521),
            .I(\c0.FRAME_MATCHER_i_20 ));
    Odrv12 I__3887 (
            .O(N__24516),
            .I(\c0.FRAME_MATCHER_i_20 ));
    CascadeMux I__3886 (
            .O(N__24511),
            .I(N__24506));
    InMux I__3885 (
            .O(N__24510),
            .I(N__24503));
    InMux I__3884 (
            .O(N__24509),
            .I(N__24500));
    InMux I__3883 (
            .O(N__24506),
            .I(N__24497));
    LocalMux I__3882 (
            .O(N__24503),
            .I(N__24492));
    LocalMux I__3881 (
            .O(N__24500),
            .I(N__24492));
    LocalMux I__3880 (
            .O(N__24497),
            .I(N__24487));
    Span4Mux_h I__3879 (
            .O(N__24492),
            .I(N__24484));
    InMux I__3878 (
            .O(N__24491),
            .I(N__24479));
    InMux I__3877 (
            .O(N__24490),
            .I(N__24479));
    Span4Mux_h I__3876 (
            .O(N__24487),
            .I(N__24476));
    Span4Mux_v I__3875 (
            .O(N__24484),
            .I(N__24472));
    LocalMux I__3874 (
            .O(N__24479),
            .I(N__24469));
    Span4Mux_h I__3873 (
            .O(N__24476),
            .I(N__24466));
    InMux I__3872 (
            .O(N__24475),
            .I(N__24463));
    Odrv4 I__3871 (
            .O(N__24472),
            .I(\c0.FRAME_MATCHER_i_4 ));
    Odrv12 I__3870 (
            .O(N__24469),
            .I(\c0.FRAME_MATCHER_i_4 ));
    Odrv4 I__3869 (
            .O(N__24466),
            .I(\c0.FRAME_MATCHER_i_4 ));
    LocalMux I__3868 (
            .O(N__24463),
            .I(\c0.FRAME_MATCHER_i_4 ));
    InMux I__3867 (
            .O(N__24454),
            .I(N__24450));
    InMux I__3866 (
            .O(N__24453),
            .I(N__24447));
    LocalMux I__3865 (
            .O(N__24450),
            .I(N__24441));
    LocalMux I__3864 (
            .O(N__24447),
            .I(N__24441));
    InMux I__3863 (
            .O(N__24446),
            .I(N__24437));
    Span4Mux_h I__3862 (
            .O(N__24441),
            .I(N__24434));
    CascadeMux I__3861 (
            .O(N__24440),
            .I(N__24430));
    LocalMux I__3860 (
            .O(N__24437),
            .I(N__24426));
    Sp12to4 I__3859 (
            .O(N__24434),
            .I(N__24423));
    InMux I__3858 (
            .O(N__24433),
            .I(N__24420));
    InMux I__3857 (
            .O(N__24430),
            .I(N__24415));
    InMux I__3856 (
            .O(N__24429),
            .I(N__24415));
    Span4Mux_h I__3855 (
            .O(N__24426),
            .I(N__24412));
    Odrv12 I__3854 (
            .O(N__24423),
            .I(\c0.FRAME_MATCHER_i_5 ));
    LocalMux I__3853 (
            .O(N__24420),
            .I(\c0.FRAME_MATCHER_i_5 ));
    LocalMux I__3852 (
            .O(N__24415),
            .I(\c0.FRAME_MATCHER_i_5 ));
    Odrv4 I__3851 (
            .O(N__24412),
            .I(\c0.FRAME_MATCHER_i_5 ));
    InMux I__3850 (
            .O(N__24403),
            .I(N__24399));
    InMux I__3849 (
            .O(N__24402),
            .I(N__24395));
    LocalMux I__3848 (
            .O(N__24399),
            .I(N__24392));
    InMux I__3847 (
            .O(N__24398),
            .I(N__24389));
    LocalMux I__3846 (
            .O(N__24395),
            .I(N__24385));
    Span4Mux_v I__3845 (
            .O(N__24392),
            .I(N__24382));
    LocalMux I__3844 (
            .O(N__24389),
            .I(N__24379));
    CascadeMux I__3843 (
            .O(N__24388),
            .I(N__24376));
    Span4Mux_v I__3842 (
            .O(N__24385),
            .I(N__24373));
    Span4Mux_s3_h I__3841 (
            .O(N__24382),
            .I(N__24368));
    Span4Mux_h I__3840 (
            .O(N__24379),
            .I(N__24368));
    InMux I__3839 (
            .O(N__24376),
            .I(N__24365));
    Span4Mux_v I__3838 (
            .O(N__24373),
            .I(N__24362));
    Span4Mux_v I__3837 (
            .O(N__24368),
            .I(N__24359));
    LocalMux I__3836 (
            .O(N__24365),
            .I(\c0.FRAME_MATCHER_i_21 ));
    Odrv4 I__3835 (
            .O(N__24362),
            .I(\c0.FRAME_MATCHER_i_21 ));
    Odrv4 I__3834 (
            .O(N__24359),
            .I(\c0.FRAME_MATCHER_i_21 ));
    CascadeMux I__3833 (
            .O(N__24352),
            .I(\c0.n30_cascade_ ));
    CascadeMux I__3832 (
            .O(N__24349),
            .I(N__24344));
    InMux I__3831 (
            .O(N__24348),
            .I(N__24341));
    CascadeMux I__3830 (
            .O(N__24347),
            .I(N__24338));
    InMux I__3829 (
            .O(N__24344),
            .I(N__24334));
    LocalMux I__3828 (
            .O(N__24341),
            .I(N__24331));
    InMux I__3827 (
            .O(N__24338),
            .I(N__24326));
    InMux I__3826 (
            .O(N__24337),
            .I(N__24326));
    LocalMux I__3825 (
            .O(N__24334),
            .I(N__24323));
    Span4Mux_v I__3824 (
            .O(N__24331),
            .I(N__24320));
    LocalMux I__3823 (
            .O(N__24326),
            .I(\c0.FRAME_MATCHER_i_13 ));
    Odrv4 I__3822 (
            .O(N__24323),
            .I(\c0.FRAME_MATCHER_i_13 ));
    Odrv4 I__3821 (
            .O(N__24320),
            .I(\c0.FRAME_MATCHER_i_13 ));
    InMux I__3820 (
            .O(N__24313),
            .I(N__24309));
    InMux I__3819 (
            .O(N__24312),
            .I(N__24306));
    LocalMux I__3818 (
            .O(N__24309),
            .I(\c0.n56 ));
    LocalMux I__3817 (
            .O(N__24306),
            .I(\c0.n56 ));
    InMux I__3816 (
            .O(N__24301),
            .I(N__24297));
    InMux I__3815 (
            .O(N__24300),
            .I(N__24294));
    LocalMux I__3814 (
            .O(N__24297),
            .I(N__24291));
    LocalMux I__3813 (
            .O(N__24294),
            .I(\c0.n446 ));
    Odrv12 I__3812 (
            .O(N__24291),
            .I(\c0.n446 ));
    CascadeMux I__3811 (
            .O(N__24286),
            .I(\c0.n446_cascade_ ));
    InMux I__3810 (
            .O(N__24283),
            .I(N__24277));
    InMux I__3809 (
            .O(N__24282),
            .I(N__24277));
    LocalMux I__3808 (
            .O(N__24277),
            .I(\c0.n456 ));
    SRMux I__3807 (
            .O(N__24274),
            .I(N__24271));
    LocalMux I__3806 (
            .O(N__24271),
            .I(N__24268));
    Span4Mux_h I__3805 (
            .O(N__24268),
            .I(N__24265));
    Odrv4 I__3804 (
            .O(N__24265),
            .I(\c0.n16371 ));
    SRMux I__3803 (
            .O(N__24262),
            .I(N__24259));
    LocalMux I__3802 (
            .O(N__24259),
            .I(N__24256));
    Odrv4 I__3801 (
            .O(N__24256),
            .I(\c0.n16453 ));
    CascadeMux I__3800 (
            .O(N__24253),
            .I(\c0.n8938_cascade_ ));
    InMux I__3799 (
            .O(N__24250),
            .I(N__24247));
    LocalMux I__3798 (
            .O(N__24247),
            .I(N__24244));
    Odrv4 I__3797 (
            .O(N__24244),
            .I(\c0.n22_adj_2164 ));
    CascadeMux I__3796 (
            .O(N__24241),
            .I(\c0.n22_adj_2164_cascade_ ));
    InMux I__3795 (
            .O(N__24238),
            .I(N__24232));
    InMux I__3794 (
            .O(N__24237),
            .I(N__24232));
    LocalMux I__3793 (
            .O(N__24232),
            .I(\c0.tx_transmit_N_1949_1 ));
    CascadeMux I__3792 (
            .O(N__24229),
            .I(\c0.n15868_cascade_ ));
    InMux I__3791 (
            .O(N__24226),
            .I(N__24223));
    LocalMux I__3790 (
            .O(N__24223),
            .I(\c0.n8631 ));
    CascadeMux I__3789 (
            .O(N__24220),
            .I(n10141_cascade_));
    InMux I__3788 (
            .O(N__24217),
            .I(\c0.n15653 ));
    InMux I__3787 (
            .O(N__24214),
            .I(\c0.n15654 ));
    InMux I__3786 (
            .O(N__24211),
            .I(\c0.n15655 ));
    InMux I__3785 (
            .O(N__24208),
            .I(\c0.n15656 ));
    InMux I__3784 (
            .O(N__24205),
            .I(\c0.n15657 ));
    InMux I__3783 (
            .O(N__24202),
            .I(\c0.n15658 ));
    InMux I__3782 (
            .O(N__24199),
            .I(\c0.n15659 ));
    InMux I__3781 (
            .O(N__24196),
            .I(N__24193));
    LocalMux I__3780 (
            .O(N__24193),
            .I(\c0.n25_adj_2324 ));
    CascadeMux I__3779 (
            .O(N__24190),
            .I(n4_adj_2458_cascade_));
    CascadeMux I__3778 (
            .O(N__24187),
            .I(N__24184));
    InMux I__3777 (
            .O(N__24184),
            .I(N__24179));
    InMux I__3776 (
            .O(N__24183),
            .I(N__24174));
    InMux I__3775 (
            .O(N__24182),
            .I(N__24174));
    LocalMux I__3774 (
            .O(N__24179),
            .I(N__24166));
    LocalMux I__3773 (
            .O(N__24174),
            .I(N__24163));
    InMux I__3772 (
            .O(N__24173),
            .I(N__24160));
    InMux I__3771 (
            .O(N__24172),
            .I(N__24157));
    CascadeMux I__3770 (
            .O(N__24171),
            .I(N__24153));
    CascadeMux I__3769 (
            .O(N__24170),
            .I(N__24150));
    InMux I__3768 (
            .O(N__24169),
            .I(N__24147));
    Span4Mux_h I__3767 (
            .O(N__24166),
            .I(N__24144));
    Span4Mux_h I__3766 (
            .O(N__24163),
            .I(N__24139));
    LocalMux I__3765 (
            .O(N__24160),
            .I(N__24139));
    LocalMux I__3764 (
            .O(N__24157),
            .I(N__24136));
    InMux I__3763 (
            .O(N__24156),
            .I(N__24131));
    InMux I__3762 (
            .O(N__24153),
            .I(N__24131));
    InMux I__3761 (
            .O(N__24150),
            .I(N__24128));
    LocalMux I__3760 (
            .O(N__24147),
            .I(r_SM_Main_0));
    Odrv4 I__3759 (
            .O(N__24144),
            .I(r_SM_Main_0));
    Odrv4 I__3758 (
            .O(N__24139),
            .I(r_SM_Main_0));
    Odrv12 I__3757 (
            .O(N__24136),
            .I(r_SM_Main_0));
    LocalMux I__3756 (
            .O(N__24131),
            .I(r_SM_Main_0));
    LocalMux I__3755 (
            .O(N__24128),
            .I(r_SM_Main_0));
    InMux I__3754 (
            .O(N__24115),
            .I(N__24110));
    InMux I__3753 (
            .O(N__24114),
            .I(N__24105));
    InMux I__3752 (
            .O(N__24113),
            .I(N__24105));
    LocalMux I__3751 (
            .O(N__24110),
            .I(N__24100));
    LocalMux I__3750 (
            .O(N__24105),
            .I(N__24097));
    InMux I__3749 (
            .O(N__24104),
            .I(N__24094));
    InMux I__3748 (
            .O(N__24103),
            .I(N__24091));
    Span4Mux_s1_v I__3747 (
            .O(N__24100),
            .I(N__24088));
    Span4Mux_h I__3746 (
            .O(N__24097),
            .I(N__24083));
    LocalMux I__3745 (
            .O(N__24094),
            .I(N__24083));
    LocalMux I__3744 (
            .O(N__24091),
            .I(n14060));
    Odrv4 I__3743 (
            .O(N__24088),
            .I(n14060));
    Odrv4 I__3742 (
            .O(N__24083),
            .I(n14060));
    CascadeMux I__3741 (
            .O(N__24076),
            .I(N__24071));
    CascadeMux I__3740 (
            .O(N__24075),
            .I(N__24068));
    InMux I__3739 (
            .O(N__24074),
            .I(N__24056));
    InMux I__3738 (
            .O(N__24071),
            .I(N__24056));
    InMux I__3737 (
            .O(N__24068),
            .I(N__24056));
    InMux I__3736 (
            .O(N__24067),
            .I(N__24053));
    InMux I__3735 (
            .O(N__24066),
            .I(N__24050));
    InMux I__3734 (
            .O(N__24065),
            .I(N__24046));
    CascadeMux I__3733 (
            .O(N__24064),
            .I(N__24040));
    InMux I__3732 (
            .O(N__24063),
            .I(N__24035));
    LocalMux I__3731 (
            .O(N__24056),
            .I(N__24030));
    LocalMux I__3730 (
            .O(N__24053),
            .I(N__24030));
    LocalMux I__3729 (
            .O(N__24050),
            .I(N__24027));
    CascadeMux I__3728 (
            .O(N__24049),
            .I(N__24024));
    LocalMux I__3727 (
            .O(N__24046),
            .I(N__24020));
    InMux I__3726 (
            .O(N__24045),
            .I(N__24015));
    InMux I__3725 (
            .O(N__24044),
            .I(N__24015));
    InMux I__3724 (
            .O(N__24043),
            .I(N__24012));
    InMux I__3723 (
            .O(N__24040),
            .I(N__24007));
    InMux I__3722 (
            .O(N__24039),
            .I(N__24007));
    InMux I__3721 (
            .O(N__24038),
            .I(N__24004));
    LocalMux I__3720 (
            .O(N__24035),
            .I(N__24001));
    Span4Mux_v I__3719 (
            .O(N__24030),
            .I(N__23996));
    Span4Mux_v I__3718 (
            .O(N__24027),
            .I(N__23996));
    InMux I__3717 (
            .O(N__24024),
            .I(N__23991));
    InMux I__3716 (
            .O(N__24023),
            .I(N__23991));
    Span4Mux_s3_h I__3715 (
            .O(N__24020),
            .I(N__23982));
    LocalMux I__3714 (
            .O(N__24015),
            .I(N__23982));
    LocalMux I__3713 (
            .O(N__24012),
            .I(N__23982));
    LocalMux I__3712 (
            .O(N__24007),
            .I(N__23982));
    LocalMux I__3711 (
            .O(N__24004),
            .I(r_SM_Main_1));
    Odrv12 I__3710 (
            .O(N__24001),
            .I(r_SM_Main_1));
    Odrv4 I__3709 (
            .O(N__23996),
            .I(r_SM_Main_1));
    LocalMux I__3708 (
            .O(N__23991),
            .I(r_SM_Main_1));
    Odrv4 I__3707 (
            .O(N__23982),
            .I(r_SM_Main_1));
    InMux I__3706 (
            .O(N__23971),
            .I(N__23965));
    InMux I__3705 (
            .O(N__23970),
            .I(N__23950));
    InMux I__3704 (
            .O(N__23969),
            .I(N__23945));
    InMux I__3703 (
            .O(N__23968),
            .I(N__23945));
    LocalMux I__3702 (
            .O(N__23965),
            .I(N__23942));
    InMux I__3701 (
            .O(N__23964),
            .I(N__23937));
    InMux I__3700 (
            .O(N__23963),
            .I(N__23937));
    InMux I__3699 (
            .O(N__23962),
            .I(N__23934));
    InMux I__3698 (
            .O(N__23961),
            .I(N__23930));
    InMux I__3697 (
            .O(N__23960),
            .I(N__23925));
    InMux I__3696 (
            .O(N__23959),
            .I(N__23925));
    InMux I__3695 (
            .O(N__23958),
            .I(N__23922));
    InMux I__3694 (
            .O(N__23957),
            .I(N__23919));
    InMux I__3693 (
            .O(N__23956),
            .I(N__23914));
    InMux I__3692 (
            .O(N__23955),
            .I(N__23914));
    InMux I__3691 (
            .O(N__23954),
            .I(N__23909));
    InMux I__3690 (
            .O(N__23953),
            .I(N__23909));
    LocalMux I__3689 (
            .O(N__23950),
            .I(N__23906));
    LocalMux I__3688 (
            .O(N__23945),
            .I(N__23903));
    Span4Mux_v I__3687 (
            .O(N__23942),
            .I(N__23896));
    LocalMux I__3686 (
            .O(N__23937),
            .I(N__23896));
    LocalMux I__3685 (
            .O(N__23934),
            .I(N__23896));
    CascadeMux I__3684 (
            .O(N__23933),
            .I(N__23893));
    LocalMux I__3683 (
            .O(N__23930),
            .I(N__23879));
    LocalMux I__3682 (
            .O(N__23925),
            .I(N__23879));
    LocalMux I__3681 (
            .O(N__23922),
            .I(N__23879));
    LocalMux I__3680 (
            .O(N__23919),
            .I(N__23879));
    LocalMux I__3679 (
            .O(N__23914),
            .I(N__23879));
    LocalMux I__3678 (
            .O(N__23909),
            .I(N__23879));
    Span4Mux_v I__3677 (
            .O(N__23906),
            .I(N__23872));
    Span4Mux_s1_h I__3676 (
            .O(N__23903),
            .I(N__23872));
    Span4Mux_s3_v I__3675 (
            .O(N__23896),
            .I(N__23869));
    InMux I__3674 (
            .O(N__23893),
            .I(N__23864));
    InMux I__3673 (
            .O(N__23892),
            .I(N__23864));
    Span4Mux_s3_v I__3672 (
            .O(N__23879),
            .I(N__23861));
    InMux I__3671 (
            .O(N__23878),
            .I(N__23858));
    InMux I__3670 (
            .O(N__23877),
            .I(N__23855));
    Span4Mux_h I__3669 (
            .O(N__23872),
            .I(N__23852));
    Span4Mux_s3_h I__3668 (
            .O(N__23869),
            .I(N__23849));
    LocalMux I__3667 (
            .O(N__23864),
            .I(N__23844));
    Span4Mux_s2_h I__3666 (
            .O(N__23861),
            .I(N__23844));
    LocalMux I__3665 (
            .O(N__23858),
            .I(r_SM_Main_2));
    LocalMux I__3664 (
            .O(N__23855),
            .I(r_SM_Main_2));
    Odrv4 I__3663 (
            .O(N__23852),
            .I(r_SM_Main_2));
    Odrv4 I__3662 (
            .O(N__23849),
            .I(r_SM_Main_2));
    Odrv4 I__3661 (
            .O(N__23844),
            .I(r_SM_Main_2));
    InMux I__3660 (
            .O(N__23833),
            .I(N__23830));
    LocalMux I__3659 (
            .O(N__23830),
            .I(N__23827));
    Odrv4 I__3658 (
            .O(N__23827),
            .I(n17395));
    InMux I__3657 (
            .O(N__23824),
            .I(N__23821));
    LocalMux I__3656 (
            .O(N__23821),
            .I(\c0.tx_active_prev ));
    InMux I__3655 (
            .O(N__23818),
            .I(N__23815));
    LocalMux I__3654 (
            .O(N__23815),
            .I(\c0.n65 ));
    CascadeMux I__3653 (
            .O(N__23812),
            .I(N__23808));
    InMux I__3652 (
            .O(N__23811),
            .I(N__23805));
    InMux I__3651 (
            .O(N__23808),
            .I(N__23802));
    LocalMux I__3650 (
            .O(N__23805),
            .I(\c0.data_in_frame_2_7 ));
    LocalMux I__3649 (
            .O(N__23802),
            .I(\c0.data_in_frame_2_7 ));
    CascadeMux I__3648 (
            .O(N__23797),
            .I(N__23793));
    CascadeMux I__3647 (
            .O(N__23796),
            .I(N__23790));
    InMux I__3646 (
            .O(N__23793),
            .I(N__23785));
    InMux I__3645 (
            .O(N__23790),
            .I(N__23785));
    LocalMux I__3644 (
            .O(N__23785),
            .I(\c0.data_in_frame_10_1 ));
    InMux I__3643 (
            .O(N__23782),
            .I(N__23775));
    InMux I__3642 (
            .O(N__23781),
            .I(N__23775));
    InMux I__3641 (
            .O(N__23780),
            .I(N__23772));
    LocalMux I__3640 (
            .O(N__23775),
            .I(\c0.n9743 ));
    LocalMux I__3639 (
            .O(N__23772),
            .I(\c0.n9743 ));
    CascadeMux I__3638 (
            .O(N__23767),
            .I(\c0.n16954_cascade_ ));
    InMux I__3637 (
            .O(N__23764),
            .I(N__23758));
    InMux I__3636 (
            .O(N__23763),
            .I(N__23758));
    LocalMux I__3635 (
            .O(N__23758),
            .I(\c0.data_in_frame_10_6 ));
    CascadeMux I__3634 (
            .O(N__23755),
            .I(\c0.n18_adj_2174_cascade_ ));
    InMux I__3633 (
            .O(N__23752),
            .I(N__23749));
    LocalMux I__3632 (
            .O(N__23749),
            .I(\c0.n17015 ));
    InMux I__3631 (
            .O(N__23746),
            .I(N__23742));
    InMux I__3630 (
            .O(N__23745),
            .I(N__23739));
    LocalMux I__3629 (
            .O(N__23742),
            .I(\c0.data_in_frame_9_4 ));
    LocalMux I__3628 (
            .O(N__23739),
            .I(\c0.data_in_frame_9_4 ));
    CascadeMux I__3627 (
            .O(N__23734),
            .I(N__23731));
    InMux I__3626 (
            .O(N__23731),
            .I(N__23728));
    LocalMux I__3625 (
            .O(N__23728),
            .I(N__23725));
    Odrv4 I__3624 (
            .O(N__23725),
            .I(\c0.n6_adj_2152 ));
    InMux I__3623 (
            .O(N__23722),
            .I(N__23718));
    InMux I__3622 (
            .O(N__23721),
            .I(N__23715));
    LocalMux I__3621 (
            .O(N__23718),
            .I(N__23709));
    LocalMux I__3620 (
            .O(N__23715),
            .I(N__23709));
    InMux I__3619 (
            .O(N__23714),
            .I(N__23706));
    Span4Mux_v I__3618 (
            .O(N__23709),
            .I(N__23703));
    LocalMux I__3617 (
            .O(N__23706),
            .I(N__23700));
    Odrv4 I__3616 (
            .O(N__23703),
            .I(\c0.n13272 ));
    Odrv12 I__3615 (
            .O(N__23700),
            .I(\c0.n13272 ));
    CascadeMux I__3614 (
            .O(N__23695),
            .I(\c0.n16882_cascade_ ));
    InMux I__3613 (
            .O(N__23692),
            .I(N__23688));
    InMux I__3612 (
            .O(N__23691),
            .I(N__23685));
    LocalMux I__3611 (
            .O(N__23688),
            .I(\c0.data_in_frame_10_4 ));
    LocalMux I__3610 (
            .O(N__23685),
            .I(\c0.data_in_frame_10_4 ));
    InMux I__3609 (
            .O(N__23680),
            .I(N__23676));
    InMux I__3608 (
            .O(N__23679),
            .I(N__23673));
    LocalMux I__3607 (
            .O(N__23676),
            .I(\c0.data_in_frame_9_6 ));
    LocalMux I__3606 (
            .O(N__23673),
            .I(\c0.data_in_frame_9_6 ));
    InMux I__3605 (
            .O(N__23668),
            .I(N__23665));
    LocalMux I__3604 (
            .O(N__23665),
            .I(N__23661));
    CascadeMux I__3603 (
            .O(N__23664),
            .I(N__23658));
    Span4Mux_h I__3602 (
            .O(N__23661),
            .I(N__23655));
    InMux I__3601 (
            .O(N__23658),
            .I(N__23652));
    Span4Mux_h I__3600 (
            .O(N__23655),
            .I(N__23649));
    LocalMux I__3599 (
            .O(N__23652),
            .I(\c0.data_in_frame_10_0 ));
    Odrv4 I__3598 (
            .O(N__23649),
            .I(\c0.data_in_frame_10_0 ));
    CascadeMux I__3597 (
            .O(N__23644),
            .I(\c0.n17013_cascade_ ));
    InMux I__3596 (
            .O(N__23641),
            .I(N__23638));
    LocalMux I__3595 (
            .O(N__23638),
            .I(N__23635));
    Odrv4 I__3594 (
            .O(N__23635),
            .I(\c0.n17013 ));
    CascadeMux I__3593 (
            .O(N__23632),
            .I(N__23629));
    InMux I__3592 (
            .O(N__23629),
            .I(N__23626));
    LocalMux I__3591 (
            .O(N__23626),
            .I(N__23622));
    InMux I__3590 (
            .O(N__23625),
            .I(N__23619));
    Span4Mux_h I__3589 (
            .O(N__23622),
            .I(N__23616));
    LocalMux I__3588 (
            .O(N__23619),
            .I(\c0.data_in_frame_9_7 ));
    Odrv4 I__3587 (
            .O(N__23616),
            .I(\c0.data_in_frame_9_7 ));
    InMux I__3586 (
            .O(N__23611),
            .I(N__23608));
    LocalMux I__3585 (
            .O(N__23608),
            .I(N__23601));
    InMux I__3584 (
            .O(N__23607),
            .I(N__23596));
    InMux I__3583 (
            .O(N__23606),
            .I(N__23596));
    InMux I__3582 (
            .O(N__23605),
            .I(N__23591));
    InMux I__3581 (
            .O(N__23604),
            .I(N__23591));
    Span4Mux_h I__3580 (
            .O(N__23601),
            .I(N__23588));
    LocalMux I__3579 (
            .O(N__23596),
            .I(data_in_3_6));
    LocalMux I__3578 (
            .O(N__23591),
            .I(data_in_3_6));
    Odrv4 I__3577 (
            .O(N__23588),
            .I(data_in_3_6));
    InMux I__3576 (
            .O(N__23581),
            .I(N__23577));
    InMux I__3575 (
            .O(N__23580),
            .I(N__23574));
    LocalMux I__3574 (
            .O(N__23577),
            .I(N__23569));
    LocalMux I__3573 (
            .O(N__23574),
            .I(N__23566));
    InMux I__3572 (
            .O(N__23573),
            .I(N__23561));
    InMux I__3571 (
            .O(N__23572),
            .I(N__23561));
    Span4Mux_h I__3570 (
            .O(N__23569),
            .I(N__23558));
    Span4Mux_v I__3569 (
            .O(N__23566),
            .I(N__23555));
    LocalMux I__3568 (
            .O(N__23561),
            .I(data_in_2_0));
    Odrv4 I__3567 (
            .O(N__23558),
            .I(data_in_2_0));
    Odrv4 I__3566 (
            .O(N__23555),
            .I(data_in_2_0));
    InMux I__3565 (
            .O(N__23548),
            .I(N__23545));
    LocalMux I__3564 (
            .O(N__23545),
            .I(N__23542));
    Odrv12 I__3563 (
            .O(N__23542),
            .I(\c0.n17268 ));
    InMux I__3562 (
            .O(N__23539),
            .I(N__23536));
    LocalMux I__3561 (
            .O(N__23536),
            .I(N__23532));
    InMux I__3560 (
            .O(N__23535),
            .I(N__23527));
    Span4Mux_h I__3559 (
            .O(N__23532),
            .I(N__23524));
    InMux I__3558 (
            .O(N__23531),
            .I(N__23519));
    InMux I__3557 (
            .O(N__23530),
            .I(N__23519));
    LocalMux I__3556 (
            .O(N__23527),
            .I(data_in_1_7));
    Odrv4 I__3555 (
            .O(N__23524),
            .I(data_in_1_7));
    LocalMux I__3554 (
            .O(N__23519),
            .I(data_in_1_7));
    CascadeMux I__3553 (
            .O(N__23512),
            .I(N__23508));
    InMux I__3552 (
            .O(N__23511),
            .I(N__23504));
    InMux I__3551 (
            .O(N__23508),
            .I(N__23499));
    InMux I__3550 (
            .O(N__23507),
            .I(N__23499));
    LocalMux I__3549 (
            .O(N__23504),
            .I(data_in_0_3));
    LocalMux I__3548 (
            .O(N__23499),
            .I(data_in_0_3));
    InMux I__3547 (
            .O(N__23494),
            .I(N__23491));
    LocalMux I__3546 (
            .O(N__23491),
            .I(N__23488));
    Odrv4 I__3545 (
            .O(N__23488),
            .I(\c0.n19_adj_2199 ));
    InMux I__3544 (
            .O(N__23485),
            .I(N__23480));
    CascadeMux I__3543 (
            .O(N__23484),
            .I(N__23476));
    InMux I__3542 (
            .O(N__23483),
            .I(N__23473));
    LocalMux I__3541 (
            .O(N__23480),
            .I(N__23470));
    InMux I__3540 (
            .O(N__23479),
            .I(N__23467));
    InMux I__3539 (
            .O(N__23476),
            .I(N__23464));
    LocalMux I__3538 (
            .O(N__23473),
            .I(N__23461));
    Span4Mux_v I__3537 (
            .O(N__23470),
            .I(N__23458));
    LocalMux I__3536 (
            .O(N__23467),
            .I(\c0.FRAME_MATCHER_i_18 ));
    LocalMux I__3535 (
            .O(N__23464),
            .I(\c0.FRAME_MATCHER_i_18 ));
    Odrv4 I__3534 (
            .O(N__23461),
            .I(\c0.FRAME_MATCHER_i_18 ));
    Odrv4 I__3533 (
            .O(N__23458),
            .I(\c0.FRAME_MATCHER_i_18 ));
    SRMux I__3532 (
            .O(N__23449),
            .I(N__23446));
    LocalMux I__3531 (
            .O(N__23446),
            .I(N__23443));
    Odrv4 I__3530 (
            .O(N__23443),
            .I(\c0.n3_adj_2239 ));
    InMux I__3529 (
            .O(N__23440),
            .I(N__23437));
    LocalMux I__3528 (
            .O(N__23437),
            .I(N__23434));
    Odrv12 I__3527 (
            .O(N__23434),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_17 ));
    InMux I__3526 (
            .O(N__23431),
            .I(N__23423));
    InMux I__3525 (
            .O(N__23430),
            .I(N__23410));
    InMux I__3524 (
            .O(N__23429),
            .I(N__23410));
    InMux I__3523 (
            .O(N__23428),
            .I(N__23403));
    InMux I__3522 (
            .O(N__23427),
            .I(N__23403));
    InMux I__3521 (
            .O(N__23426),
            .I(N__23403));
    LocalMux I__3520 (
            .O(N__23423),
            .I(N__23399));
    InMux I__3519 (
            .O(N__23422),
            .I(N__23394));
    InMux I__3518 (
            .O(N__23421),
            .I(N__23394));
    InMux I__3517 (
            .O(N__23420),
            .I(N__23391));
    InMux I__3516 (
            .O(N__23419),
            .I(N__23388));
    InMux I__3515 (
            .O(N__23418),
            .I(N__23379));
    InMux I__3514 (
            .O(N__23417),
            .I(N__23379));
    InMux I__3513 (
            .O(N__23416),
            .I(N__23379));
    InMux I__3512 (
            .O(N__23415),
            .I(N__23379));
    LocalMux I__3511 (
            .O(N__23410),
            .I(N__23359));
    LocalMux I__3510 (
            .O(N__23403),
            .I(N__23359));
    InMux I__3509 (
            .O(N__23402),
            .I(N__23348));
    Span4Mux_v I__3508 (
            .O(N__23399),
            .I(N__23339));
    LocalMux I__3507 (
            .O(N__23394),
            .I(N__23339));
    LocalMux I__3506 (
            .O(N__23391),
            .I(N__23339));
    LocalMux I__3505 (
            .O(N__23388),
            .I(N__23339));
    LocalMux I__3504 (
            .O(N__23379),
            .I(N__23336));
    InMux I__3503 (
            .O(N__23378),
            .I(N__23327));
    InMux I__3502 (
            .O(N__23377),
            .I(N__23327));
    InMux I__3501 (
            .O(N__23376),
            .I(N__23327));
    InMux I__3500 (
            .O(N__23375),
            .I(N__23327));
    InMux I__3499 (
            .O(N__23374),
            .I(N__23312));
    InMux I__3498 (
            .O(N__23373),
            .I(N__23312));
    InMux I__3497 (
            .O(N__23372),
            .I(N__23312));
    InMux I__3496 (
            .O(N__23371),
            .I(N__23312));
    InMux I__3495 (
            .O(N__23370),
            .I(N__23312));
    InMux I__3494 (
            .O(N__23369),
            .I(N__23312));
    InMux I__3493 (
            .O(N__23368),
            .I(N__23312));
    InMux I__3492 (
            .O(N__23367),
            .I(N__23303));
    InMux I__3491 (
            .O(N__23366),
            .I(N__23303));
    InMux I__3490 (
            .O(N__23365),
            .I(N__23303));
    InMux I__3489 (
            .O(N__23364),
            .I(N__23303));
    Span4Mux_v I__3488 (
            .O(N__23359),
            .I(N__23300));
    InMux I__3487 (
            .O(N__23358),
            .I(N__23291));
    InMux I__3486 (
            .O(N__23357),
            .I(N__23291));
    InMux I__3485 (
            .O(N__23356),
            .I(N__23291));
    InMux I__3484 (
            .O(N__23355),
            .I(N__23291));
    InMux I__3483 (
            .O(N__23354),
            .I(N__23282));
    InMux I__3482 (
            .O(N__23353),
            .I(N__23282));
    InMux I__3481 (
            .O(N__23352),
            .I(N__23282));
    InMux I__3480 (
            .O(N__23351),
            .I(N__23282));
    LocalMux I__3479 (
            .O(N__23348),
            .I(N__23277));
    Span4Mux_v I__3478 (
            .O(N__23339),
            .I(N__23277));
    Odrv4 I__3477 (
            .O(N__23336),
            .I(\c0.n127_adj_2136 ));
    LocalMux I__3476 (
            .O(N__23327),
            .I(\c0.n127_adj_2136 ));
    LocalMux I__3475 (
            .O(N__23312),
            .I(\c0.n127_adj_2136 ));
    LocalMux I__3474 (
            .O(N__23303),
            .I(\c0.n127_adj_2136 ));
    Odrv4 I__3473 (
            .O(N__23300),
            .I(\c0.n127_adj_2136 ));
    LocalMux I__3472 (
            .O(N__23291),
            .I(\c0.n127_adj_2136 ));
    LocalMux I__3471 (
            .O(N__23282),
            .I(\c0.n127_adj_2136 ));
    Odrv4 I__3470 (
            .O(N__23277),
            .I(\c0.n127_adj_2136 ));
    InMux I__3469 (
            .O(N__23260),
            .I(N__23246));
    InMux I__3468 (
            .O(N__23259),
            .I(N__23246));
    InMux I__3467 (
            .O(N__23258),
            .I(N__23246));
    InMux I__3466 (
            .O(N__23257),
            .I(N__23241));
    InMux I__3465 (
            .O(N__23256),
            .I(N__23241));
    InMux I__3464 (
            .O(N__23255),
            .I(N__23226));
    InMux I__3463 (
            .O(N__23254),
            .I(N__23226));
    InMux I__3462 (
            .O(N__23253),
            .I(N__23226));
    LocalMux I__3461 (
            .O(N__23246),
            .I(N__23218));
    LocalMux I__3460 (
            .O(N__23241),
            .I(N__23218));
    InMux I__3459 (
            .O(N__23240),
            .I(N__23215));
    InMux I__3458 (
            .O(N__23239),
            .I(N__23206));
    InMux I__3457 (
            .O(N__23238),
            .I(N__23206));
    InMux I__3456 (
            .O(N__23237),
            .I(N__23206));
    InMux I__3455 (
            .O(N__23236),
            .I(N__23206));
    CascadeMux I__3454 (
            .O(N__23235),
            .I(N__23192));
    InMux I__3453 (
            .O(N__23234),
            .I(N__23177));
    InMux I__3452 (
            .O(N__23233),
            .I(N__23177));
    LocalMux I__3451 (
            .O(N__23226),
            .I(N__23174));
    InMux I__3450 (
            .O(N__23225),
            .I(N__23171));
    InMux I__3449 (
            .O(N__23224),
            .I(N__23166));
    InMux I__3448 (
            .O(N__23223),
            .I(N__23166));
    Span4Mux_h I__3447 (
            .O(N__23218),
            .I(N__23163));
    LocalMux I__3446 (
            .O(N__23215),
            .I(N__23160));
    LocalMux I__3445 (
            .O(N__23206),
            .I(N__23157));
    InMux I__3444 (
            .O(N__23205),
            .I(N__23148));
    InMux I__3443 (
            .O(N__23204),
            .I(N__23148));
    InMux I__3442 (
            .O(N__23203),
            .I(N__23148));
    InMux I__3441 (
            .O(N__23202),
            .I(N__23148));
    InMux I__3440 (
            .O(N__23201),
            .I(N__23133));
    InMux I__3439 (
            .O(N__23200),
            .I(N__23133));
    InMux I__3438 (
            .O(N__23199),
            .I(N__23133));
    InMux I__3437 (
            .O(N__23198),
            .I(N__23133));
    InMux I__3436 (
            .O(N__23197),
            .I(N__23133));
    InMux I__3435 (
            .O(N__23196),
            .I(N__23133));
    InMux I__3434 (
            .O(N__23195),
            .I(N__23133));
    InMux I__3433 (
            .O(N__23192),
            .I(N__23124));
    InMux I__3432 (
            .O(N__23191),
            .I(N__23124));
    InMux I__3431 (
            .O(N__23190),
            .I(N__23124));
    InMux I__3430 (
            .O(N__23189),
            .I(N__23124));
    InMux I__3429 (
            .O(N__23188),
            .I(N__23113));
    InMux I__3428 (
            .O(N__23187),
            .I(N__23113));
    InMux I__3427 (
            .O(N__23186),
            .I(N__23113));
    InMux I__3426 (
            .O(N__23185),
            .I(N__23113));
    InMux I__3425 (
            .O(N__23184),
            .I(N__23113));
    InMux I__3424 (
            .O(N__23183),
            .I(N__23108));
    InMux I__3423 (
            .O(N__23182),
            .I(N__23108));
    LocalMux I__3422 (
            .O(N__23177),
            .I(N__23103));
    Span4Mux_h I__3421 (
            .O(N__23174),
            .I(N__23103));
    LocalMux I__3420 (
            .O(N__23171),
            .I(N__23098));
    LocalMux I__3419 (
            .O(N__23166),
            .I(N__23098));
    Odrv4 I__3418 (
            .O(N__23163),
            .I(n127));
    Odrv4 I__3417 (
            .O(N__23160),
            .I(n127));
    Odrv4 I__3416 (
            .O(N__23157),
            .I(n127));
    LocalMux I__3415 (
            .O(N__23148),
            .I(n127));
    LocalMux I__3414 (
            .O(N__23133),
            .I(n127));
    LocalMux I__3413 (
            .O(N__23124),
            .I(n127));
    LocalMux I__3412 (
            .O(N__23113),
            .I(n127));
    LocalMux I__3411 (
            .O(N__23108),
            .I(n127));
    Odrv4 I__3410 (
            .O(N__23103),
            .I(n127));
    Odrv12 I__3409 (
            .O(N__23098),
            .I(n127));
    InMux I__3408 (
            .O(N__23077),
            .I(N__23074));
    LocalMux I__3407 (
            .O(N__23074),
            .I(N__23071));
    Span4Mux_h I__3406 (
            .O(N__23071),
            .I(N__23068));
    Odrv4 I__3405 (
            .O(N__23068),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_16 ));
    CascadeMux I__3404 (
            .O(N__23065),
            .I(N__23053));
    CascadeMux I__3403 (
            .O(N__23064),
            .I(N__23050));
    InMux I__3402 (
            .O(N__23063),
            .I(N__23022));
    InMux I__3401 (
            .O(N__23062),
            .I(N__23022));
    InMux I__3400 (
            .O(N__23061),
            .I(N__23022));
    InMux I__3399 (
            .O(N__23060),
            .I(N__23022));
    InMux I__3398 (
            .O(N__23059),
            .I(N__23022));
    InMux I__3397 (
            .O(N__23058),
            .I(N__23022));
    InMux I__3396 (
            .O(N__23057),
            .I(N__23017));
    InMux I__3395 (
            .O(N__23056),
            .I(N__23017));
    InMux I__3394 (
            .O(N__23053),
            .I(N__23009));
    InMux I__3393 (
            .O(N__23050),
            .I(N__23009));
    InMux I__3392 (
            .O(N__23049),
            .I(N__23009));
    CascadeMux I__3391 (
            .O(N__23048),
            .I(N__23003));
    CascadeMux I__3390 (
            .O(N__23047),
            .I(N__23000));
    CascadeMux I__3389 (
            .O(N__23046),
            .I(N__22997));
    InMux I__3388 (
            .O(N__23045),
            .I(N__22983));
    InMux I__3387 (
            .O(N__23044),
            .I(N__22983));
    InMux I__3386 (
            .O(N__23043),
            .I(N__22980));
    CascadeMux I__3385 (
            .O(N__23042),
            .I(N__22972));
    InMux I__3384 (
            .O(N__23041),
            .I(N__22966));
    InMux I__3383 (
            .O(N__23040),
            .I(N__22966));
    InMux I__3382 (
            .O(N__23039),
            .I(N__22955));
    InMux I__3381 (
            .O(N__23038),
            .I(N__22955));
    InMux I__3380 (
            .O(N__23037),
            .I(N__22955));
    InMux I__3379 (
            .O(N__23036),
            .I(N__22955));
    InMux I__3378 (
            .O(N__23035),
            .I(N__22955));
    LocalMux I__3377 (
            .O(N__23022),
            .I(N__22949));
    LocalMux I__3376 (
            .O(N__23017),
            .I(N__22949));
    InMux I__3375 (
            .O(N__23016),
            .I(N__22946));
    LocalMux I__3374 (
            .O(N__23009),
            .I(N__22943));
    InMux I__3373 (
            .O(N__23008),
            .I(N__22928));
    InMux I__3372 (
            .O(N__23007),
            .I(N__22928));
    InMux I__3371 (
            .O(N__23006),
            .I(N__22928));
    InMux I__3370 (
            .O(N__23003),
            .I(N__22928));
    InMux I__3369 (
            .O(N__23000),
            .I(N__22928));
    InMux I__3368 (
            .O(N__22997),
            .I(N__22928));
    InMux I__3367 (
            .O(N__22996),
            .I(N__22928));
    CascadeMux I__3366 (
            .O(N__22995),
            .I(N__22922));
    CascadeMux I__3365 (
            .O(N__22994),
            .I(N__22919));
    CascadeMux I__3364 (
            .O(N__22993),
            .I(N__22916));
    CascadeMux I__3363 (
            .O(N__22992),
            .I(N__22912));
    CascadeMux I__3362 (
            .O(N__22991),
            .I(N__22909));
    CascadeMux I__3361 (
            .O(N__22990),
            .I(N__22906));
    CascadeMux I__3360 (
            .O(N__22989),
            .I(N__22892));
    CascadeMux I__3359 (
            .O(N__22988),
            .I(N__22888));
    LocalMux I__3358 (
            .O(N__22983),
            .I(N__22881));
    LocalMux I__3357 (
            .O(N__22980),
            .I(N__22881));
    InMux I__3356 (
            .O(N__22979),
            .I(N__22866));
    InMux I__3355 (
            .O(N__22978),
            .I(N__22866));
    InMux I__3354 (
            .O(N__22977),
            .I(N__22866));
    InMux I__3353 (
            .O(N__22976),
            .I(N__22866));
    InMux I__3352 (
            .O(N__22975),
            .I(N__22866));
    InMux I__3351 (
            .O(N__22972),
            .I(N__22866));
    InMux I__3350 (
            .O(N__22971),
            .I(N__22866));
    LocalMux I__3349 (
            .O(N__22966),
            .I(N__22863));
    LocalMux I__3348 (
            .O(N__22955),
            .I(N__22860));
    CascadeMux I__3347 (
            .O(N__22954),
            .I(N__22857));
    Span4Mux_v I__3346 (
            .O(N__22949),
            .I(N__22852));
    LocalMux I__3345 (
            .O(N__22946),
            .I(N__22849));
    Span4Mux_v I__3344 (
            .O(N__22943),
            .I(N__22844));
    LocalMux I__3343 (
            .O(N__22928),
            .I(N__22844));
    InMux I__3342 (
            .O(N__22927),
            .I(N__22829));
    InMux I__3341 (
            .O(N__22926),
            .I(N__22829));
    InMux I__3340 (
            .O(N__22925),
            .I(N__22829));
    InMux I__3339 (
            .O(N__22922),
            .I(N__22829));
    InMux I__3338 (
            .O(N__22919),
            .I(N__22829));
    InMux I__3337 (
            .O(N__22916),
            .I(N__22829));
    InMux I__3336 (
            .O(N__22915),
            .I(N__22829));
    InMux I__3335 (
            .O(N__22912),
            .I(N__22814));
    InMux I__3334 (
            .O(N__22909),
            .I(N__22814));
    InMux I__3333 (
            .O(N__22906),
            .I(N__22814));
    InMux I__3332 (
            .O(N__22905),
            .I(N__22814));
    InMux I__3331 (
            .O(N__22904),
            .I(N__22814));
    InMux I__3330 (
            .O(N__22903),
            .I(N__22814));
    InMux I__3329 (
            .O(N__22902),
            .I(N__22814));
    InMux I__3328 (
            .O(N__22901),
            .I(N__22799));
    InMux I__3327 (
            .O(N__22900),
            .I(N__22799));
    InMux I__3326 (
            .O(N__22899),
            .I(N__22799));
    InMux I__3325 (
            .O(N__22898),
            .I(N__22799));
    InMux I__3324 (
            .O(N__22897),
            .I(N__22799));
    InMux I__3323 (
            .O(N__22896),
            .I(N__22799));
    InMux I__3322 (
            .O(N__22895),
            .I(N__22799));
    InMux I__3321 (
            .O(N__22892),
            .I(N__22788));
    InMux I__3320 (
            .O(N__22891),
            .I(N__22788));
    InMux I__3319 (
            .O(N__22888),
            .I(N__22788));
    InMux I__3318 (
            .O(N__22887),
            .I(N__22788));
    InMux I__3317 (
            .O(N__22886),
            .I(N__22788));
    Span4Mux_v I__3316 (
            .O(N__22881),
            .I(N__22779));
    LocalMux I__3315 (
            .O(N__22866),
            .I(N__22779));
    Span4Mux_h I__3314 (
            .O(N__22863),
            .I(N__22779));
    Span4Mux_h I__3313 (
            .O(N__22860),
            .I(N__22779));
    InMux I__3312 (
            .O(N__22857),
            .I(N__22772));
    InMux I__3311 (
            .O(N__22856),
            .I(N__22772));
    InMux I__3310 (
            .O(N__22855),
            .I(N__22772));
    Odrv4 I__3309 (
            .O(N__22852),
            .I(n127_adj_2418));
    Odrv4 I__3308 (
            .O(N__22849),
            .I(n127_adj_2418));
    Odrv4 I__3307 (
            .O(N__22844),
            .I(n127_adj_2418));
    LocalMux I__3306 (
            .O(N__22829),
            .I(n127_adj_2418));
    LocalMux I__3305 (
            .O(N__22814),
            .I(n127_adj_2418));
    LocalMux I__3304 (
            .O(N__22799),
            .I(n127_adj_2418));
    LocalMux I__3303 (
            .O(N__22788),
            .I(n127_adj_2418));
    Odrv4 I__3302 (
            .O(N__22779),
            .I(n127_adj_2418));
    LocalMux I__3301 (
            .O(N__22772),
            .I(n127_adj_2418));
    CascadeMux I__3300 (
            .O(N__22753),
            .I(N__22748));
    InMux I__3299 (
            .O(N__22752),
            .I(N__22745));
    CascadeMux I__3298 (
            .O(N__22751),
            .I(N__22742));
    InMux I__3297 (
            .O(N__22748),
            .I(N__22739));
    LocalMux I__3296 (
            .O(N__22745),
            .I(N__22736));
    InMux I__3295 (
            .O(N__22742),
            .I(N__22733));
    LocalMux I__3294 (
            .O(N__22739),
            .I(N__22730));
    Span4Mux_v I__3293 (
            .O(N__22736),
            .I(N__22727));
    LocalMux I__3292 (
            .O(N__22733),
            .I(N__22721));
    Sp12to4 I__3291 (
            .O(N__22730),
            .I(N__22721));
    Span4Mux_v I__3290 (
            .O(N__22727),
            .I(N__22718));
    InMux I__3289 (
            .O(N__22726),
            .I(N__22715));
    Odrv12 I__3288 (
            .O(N__22721),
            .I(\c0.FRAME_MATCHER_i_16 ));
    Odrv4 I__3287 (
            .O(N__22718),
            .I(\c0.FRAME_MATCHER_i_16 ));
    LocalMux I__3286 (
            .O(N__22715),
            .I(\c0.FRAME_MATCHER_i_16 ));
    InMux I__3285 (
            .O(N__22708),
            .I(N__22683));
    InMux I__3284 (
            .O(N__22707),
            .I(N__22683));
    InMux I__3283 (
            .O(N__22706),
            .I(N__22683));
    InMux I__3282 (
            .O(N__22705),
            .I(N__22676));
    InMux I__3281 (
            .O(N__22704),
            .I(N__22676));
    InMux I__3280 (
            .O(N__22703),
            .I(N__22676));
    CascadeMux I__3279 (
            .O(N__22702),
            .I(N__22669));
    CascadeMux I__3278 (
            .O(N__22701),
            .I(N__22662));
    CascadeMux I__3277 (
            .O(N__22700),
            .I(N__22659));
    InMux I__3276 (
            .O(N__22699),
            .I(N__22652));
    InMux I__3275 (
            .O(N__22698),
            .I(N__22652));
    InMux I__3274 (
            .O(N__22697),
            .I(N__22652));
    InMux I__3273 (
            .O(N__22696),
            .I(N__22641));
    InMux I__3272 (
            .O(N__22695),
            .I(N__22641));
    InMux I__3271 (
            .O(N__22694),
            .I(N__22641));
    InMux I__3270 (
            .O(N__22693),
            .I(N__22641));
    InMux I__3269 (
            .O(N__22692),
            .I(N__22641));
    InMux I__3268 (
            .O(N__22691),
            .I(N__22636));
    InMux I__3267 (
            .O(N__22690),
            .I(N__22636));
    LocalMux I__3266 (
            .O(N__22683),
            .I(N__22633));
    LocalMux I__3265 (
            .O(N__22676),
            .I(N__22630));
    InMux I__3264 (
            .O(N__22675),
            .I(N__22621));
    InMux I__3263 (
            .O(N__22674),
            .I(N__22621));
    InMux I__3262 (
            .O(N__22673),
            .I(N__22621));
    InMux I__3261 (
            .O(N__22672),
            .I(N__22621));
    InMux I__3260 (
            .O(N__22669),
            .I(N__22618));
    InMux I__3259 (
            .O(N__22668),
            .I(N__22615));
    InMux I__3258 (
            .O(N__22667),
            .I(N__22604));
    InMux I__3257 (
            .O(N__22666),
            .I(N__22604));
    InMux I__3256 (
            .O(N__22665),
            .I(N__22604));
    InMux I__3255 (
            .O(N__22662),
            .I(N__22604));
    InMux I__3254 (
            .O(N__22659),
            .I(N__22604));
    LocalMux I__3253 (
            .O(N__22652),
            .I(N__22599));
    LocalMux I__3252 (
            .O(N__22641),
            .I(N__22599));
    LocalMux I__3251 (
            .O(N__22636),
            .I(N__22594));
    Span4Mux_v I__3250 (
            .O(N__22633),
            .I(N__22594));
    Span4Mux_v I__3249 (
            .O(N__22630),
            .I(N__22587));
    LocalMux I__3248 (
            .O(N__22621),
            .I(N__22587));
    LocalMux I__3247 (
            .O(N__22618),
            .I(N__22587));
    LocalMux I__3246 (
            .O(N__22615),
            .I(\c0.n7212 ));
    LocalMux I__3245 (
            .O(N__22604),
            .I(\c0.n7212 ));
    Odrv4 I__3244 (
            .O(N__22599),
            .I(\c0.n7212 ));
    Odrv4 I__3243 (
            .O(N__22594),
            .I(\c0.n7212 ));
    Odrv4 I__3242 (
            .O(N__22587),
            .I(\c0.n7212 ));
    SRMux I__3241 (
            .O(N__22576),
            .I(N__22573));
    LocalMux I__3240 (
            .O(N__22573),
            .I(N__22570));
    Span12Mux_v I__3239 (
            .O(N__22570),
            .I(N__22567));
    Odrv12 I__3238 (
            .O(N__22567),
            .I(\c0.n3_adj_2241 ));
    InMux I__3237 (
            .O(N__22564),
            .I(N__22560));
    CascadeMux I__3236 (
            .O(N__22563),
            .I(N__22557));
    LocalMux I__3235 (
            .O(N__22560),
            .I(N__22554));
    InMux I__3234 (
            .O(N__22557),
            .I(N__22551));
    Span4Mux_h I__3233 (
            .O(N__22554),
            .I(N__22548));
    LocalMux I__3232 (
            .O(N__22551),
            .I(\c0.data_in_frame_9_2 ));
    Odrv4 I__3231 (
            .O(N__22548),
            .I(\c0.data_in_frame_9_2 ));
    CascadeMux I__3230 (
            .O(N__22543),
            .I(N__22540));
    InMux I__3229 (
            .O(N__22540),
            .I(N__22537));
    LocalMux I__3228 (
            .O(N__22537),
            .I(N__22534));
    Odrv4 I__3227 (
            .O(N__22534),
            .I(\c0.n15939 ));
    InMux I__3226 (
            .O(N__22531),
            .I(N__22528));
    LocalMux I__3225 (
            .O(N__22528),
            .I(N__22525));
    Span4Mux_v I__3224 (
            .O(N__22525),
            .I(N__22522));
    Odrv4 I__3223 (
            .O(N__22522),
            .I(\c0.n17264 ));
    InMux I__3222 (
            .O(N__22519),
            .I(N__22516));
    LocalMux I__3221 (
            .O(N__22516),
            .I(N__22513));
    Span4Mux_h I__3220 (
            .O(N__22513),
            .I(N__22510));
    Sp12to4 I__3219 (
            .O(N__22510),
            .I(N__22507));
    Odrv12 I__3218 (
            .O(N__22507),
            .I(\c0.n9493 ));
    CascadeMux I__3217 (
            .O(N__22504),
            .I(\c0.n12_cascade_ ));
    CascadeMux I__3216 (
            .O(N__22501),
            .I(N__22497));
    InMux I__3215 (
            .O(N__22500),
            .I(N__22489));
    InMux I__3214 (
            .O(N__22497),
            .I(N__22486));
    InMux I__3213 (
            .O(N__22496),
            .I(N__22483));
    InMux I__3212 (
            .O(N__22495),
            .I(N__22480));
    InMux I__3211 (
            .O(N__22494),
            .I(N__22477));
    InMux I__3210 (
            .O(N__22493),
            .I(N__22474));
    InMux I__3209 (
            .O(N__22492),
            .I(N__22471));
    LocalMux I__3208 (
            .O(N__22489),
            .I(N__22466));
    LocalMux I__3207 (
            .O(N__22486),
            .I(N__22466));
    LocalMux I__3206 (
            .O(N__22483),
            .I(N__22463));
    LocalMux I__3205 (
            .O(N__22480),
            .I(N__22460));
    LocalMux I__3204 (
            .O(N__22477),
            .I(N__22453));
    LocalMux I__3203 (
            .O(N__22474),
            .I(N__22453));
    LocalMux I__3202 (
            .O(N__22471),
            .I(N__22453));
    Span4Mux_v I__3201 (
            .O(N__22466),
            .I(N__22450));
    Span4Mux_h I__3200 (
            .O(N__22463),
            .I(N__22447));
    Span4Mux_h I__3199 (
            .O(N__22460),
            .I(N__22442));
    Span4Mux_h I__3198 (
            .O(N__22453),
            .I(N__22442));
    Odrv4 I__3197 (
            .O(N__22450),
            .I(\c0.FRAME_MATCHER_i_31 ));
    Odrv4 I__3196 (
            .O(N__22447),
            .I(\c0.FRAME_MATCHER_i_31 ));
    Odrv4 I__3195 (
            .O(N__22442),
            .I(\c0.FRAME_MATCHER_i_31 ));
    CascadeMux I__3194 (
            .O(N__22435),
            .I(n127_adj_2418_cascade_));
    InMux I__3193 (
            .O(N__22432),
            .I(N__22429));
    LocalMux I__3192 (
            .O(N__22429),
            .I(\c0.n17240 ));
    InMux I__3191 (
            .O(N__22426),
            .I(N__22422));
    InMux I__3190 (
            .O(N__22425),
            .I(N__22419));
    LocalMux I__3189 (
            .O(N__22422),
            .I(N__22413));
    LocalMux I__3188 (
            .O(N__22419),
            .I(N__22413));
    CascadeMux I__3187 (
            .O(N__22418),
            .I(N__22410));
    Span4Mux_v I__3186 (
            .O(N__22413),
            .I(N__22405));
    InMux I__3185 (
            .O(N__22410),
            .I(N__22400));
    InMux I__3184 (
            .O(N__22409),
            .I(N__22400));
    InMux I__3183 (
            .O(N__22408),
            .I(N__22397));
    Sp12to4 I__3182 (
            .O(N__22405),
            .I(N__22392));
    LocalMux I__3181 (
            .O(N__22400),
            .I(N__22392));
    LocalMux I__3180 (
            .O(N__22397),
            .I(data_in_1_1));
    Odrv12 I__3179 (
            .O(N__22392),
            .I(data_in_1_1));
    CascadeMux I__3178 (
            .O(N__22387),
            .I(N__22384));
    InMux I__3177 (
            .O(N__22384),
            .I(N__22378));
    InMux I__3176 (
            .O(N__22383),
            .I(N__22378));
    LocalMux I__3175 (
            .O(N__22378),
            .I(\c0.n9482 ));
    InMux I__3174 (
            .O(N__22375),
            .I(N__22372));
    LocalMux I__3173 (
            .O(N__22372),
            .I(N__22368));
    InMux I__3172 (
            .O(N__22371),
            .I(N__22365));
    Span4Mux_h I__3171 (
            .O(N__22368),
            .I(N__22362));
    LocalMux I__3170 (
            .O(N__22365),
            .I(N__22359));
    Odrv4 I__3169 (
            .O(N__22362),
            .I(\c0.n9490 ));
    Odrv4 I__3168 (
            .O(N__22359),
            .I(\c0.n9490 ));
    InMux I__3167 (
            .O(N__22354),
            .I(N__22350));
    InMux I__3166 (
            .O(N__22353),
            .I(N__22346));
    LocalMux I__3165 (
            .O(N__22350),
            .I(N__22343));
    InMux I__3164 (
            .O(N__22349),
            .I(N__22340));
    LocalMux I__3163 (
            .O(N__22346),
            .I(N__22337));
    Span4Mux_h I__3162 (
            .O(N__22343),
            .I(N__22332));
    LocalMux I__3161 (
            .O(N__22340),
            .I(N__22332));
    Odrv12 I__3160 (
            .O(N__22337),
            .I(n16795));
    Odrv4 I__3159 (
            .O(N__22332),
            .I(n16795));
    CascadeMux I__3158 (
            .O(N__22327),
            .I(n127_cascade_));
    InMux I__3157 (
            .O(N__22324),
            .I(N__22321));
    LocalMux I__3156 (
            .O(N__22321),
            .I(N__22318));
    Span4Mux_h I__3155 (
            .O(N__22318),
            .I(N__22315));
    Odrv4 I__3154 (
            .O(N__22315),
            .I(\c0.n2 ));
    CascadeMux I__3153 (
            .O(N__22312),
            .I(\c0.n2_cascade_ ));
    CascadeMux I__3152 (
            .O(N__22309),
            .I(N__22306));
    InMux I__3151 (
            .O(N__22306),
            .I(N__22303));
    LocalMux I__3150 (
            .O(N__22303),
            .I(N__22300));
    Span4Mux_h I__3149 (
            .O(N__22300),
            .I(N__22296));
    InMux I__3148 (
            .O(N__22299),
            .I(N__22293));
    Odrv4 I__3147 (
            .O(N__22296),
            .I(n9435));
    LocalMux I__3146 (
            .O(N__22293),
            .I(n9435));
    CascadeMux I__3145 (
            .O(N__22288),
            .I(N__22284));
    CascadeMux I__3144 (
            .O(N__22287),
            .I(N__22281));
    InMux I__3143 (
            .O(N__22284),
            .I(N__22270));
    InMux I__3142 (
            .O(N__22281),
            .I(N__22270));
    InMux I__3141 (
            .O(N__22280),
            .I(N__22270));
    InMux I__3140 (
            .O(N__22279),
            .I(N__22270));
    LocalMux I__3139 (
            .O(N__22270),
            .I(N__22267));
    Span4Mux_s3_h I__3138 (
            .O(N__22267),
            .I(N__22264));
    Span4Mux_v I__3137 (
            .O(N__22264),
            .I(N__22261));
    Odrv4 I__3136 (
            .O(N__22261),
            .I(n7198));
    InMux I__3135 (
            .O(N__22258),
            .I(N__22255));
    LocalMux I__3134 (
            .O(N__22255),
            .I(N__22252));
    Odrv4 I__3133 (
            .O(N__22252),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_18 ));
    InMux I__3132 (
            .O(N__22249),
            .I(N__22246));
    LocalMux I__3131 (
            .O(N__22246),
            .I(N__22243));
    Odrv4 I__3130 (
            .O(N__22243),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_18 ));
    InMux I__3129 (
            .O(N__22240),
            .I(N__22237));
    LocalMux I__3128 (
            .O(N__22237),
            .I(N__22234));
    Span4Mux_h I__3127 (
            .O(N__22234),
            .I(N__22231));
    Odrv4 I__3126 (
            .O(N__22231),
            .I(\c0.n12_adj_2158 ));
    CascadeMux I__3125 (
            .O(N__22228),
            .I(\c0.n9488_cascade_ ));
    InMux I__3124 (
            .O(N__22225),
            .I(N__22222));
    LocalMux I__3123 (
            .O(N__22222),
            .I(N__22219));
    Span4Mux_h I__3122 (
            .O(N__22219),
            .I(N__22216));
    Odrv4 I__3121 (
            .O(N__22216),
            .I(\c0.n17262 ));
    InMux I__3120 (
            .O(N__22213),
            .I(N__22210));
    LocalMux I__3119 (
            .O(N__22210),
            .I(\c0.n17256 ));
    InMux I__3118 (
            .O(N__22207),
            .I(N__22200));
    InMux I__3117 (
            .O(N__22206),
            .I(N__22200));
    CascadeMux I__3116 (
            .O(N__22205),
            .I(N__22197));
    LocalMux I__3115 (
            .O(N__22200),
            .I(N__22194));
    InMux I__3114 (
            .O(N__22197),
            .I(N__22191));
    Span4Mux_v I__3113 (
            .O(N__22194),
            .I(N__22188));
    LocalMux I__3112 (
            .O(N__22191),
            .I(data_in_0_0));
    Odrv4 I__3111 (
            .O(N__22188),
            .I(data_in_0_0));
    InMux I__3110 (
            .O(N__22183),
            .I(N__22179));
    InMux I__3109 (
            .O(N__22182),
            .I(N__22176));
    LocalMux I__3108 (
            .O(N__22179),
            .I(\c0.n9485 ));
    LocalMux I__3107 (
            .O(N__22176),
            .I(\c0.n9485 ));
    CascadeMux I__3106 (
            .O(N__22171),
            .I(\c0.n10_adj_2149_cascade_ ));
    InMux I__3105 (
            .O(N__22168),
            .I(N__22165));
    LocalMux I__3104 (
            .O(N__22165),
            .I(N__22159));
    InMux I__3103 (
            .O(N__22164),
            .I(N__22156));
    CascadeMux I__3102 (
            .O(N__22163),
            .I(N__22153));
    InMux I__3101 (
            .O(N__22162),
            .I(N__22150));
    Span4Mux_h I__3100 (
            .O(N__22159),
            .I(N__22147));
    LocalMux I__3099 (
            .O(N__22156),
            .I(N__22144));
    InMux I__3098 (
            .O(N__22153),
            .I(N__22141));
    LocalMux I__3097 (
            .O(N__22150),
            .I(N__22138));
    Span4Mux_v I__3096 (
            .O(N__22147),
            .I(N__22135));
    Span4Mux_h I__3095 (
            .O(N__22144),
            .I(N__22132));
    LocalMux I__3094 (
            .O(N__22141),
            .I(\c0.FRAME_MATCHER_i_29 ));
    Odrv12 I__3093 (
            .O(N__22138),
            .I(\c0.FRAME_MATCHER_i_29 ));
    Odrv4 I__3092 (
            .O(N__22135),
            .I(\c0.FRAME_MATCHER_i_29 ));
    Odrv4 I__3091 (
            .O(N__22132),
            .I(\c0.FRAME_MATCHER_i_29 ));
    InMux I__3090 (
            .O(N__22123),
            .I(N__22120));
    LocalMux I__3089 (
            .O(N__22120),
            .I(N__22117));
    Span4Mux_h I__3088 (
            .O(N__22117),
            .I(N__22114));
    Odrv4 I__3087 (
            .O(N__22114),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_29 ));
    InMux I__3086 (
            .O(N__22111),
            .I(N__22107));
    InMux I__3085 (
            .O(N__22110),
            .I(N__22103));
    LocalMux I__3084 (
            .O(N__22107),
            .I(N__22100));
    InMux I__3083 (
            .O(N__22106),
            .I(N__22096));
    LocalMux I__3082 (
            .O(N__22103),
            .I(N__22091));
    Span4Mux_h I__3081 (
            .O(N__22100),
            .I(N__22091));
    InMux I__3080 (
            .O(N__22099),
            .I(N__22088));
    LocalMux I__3079 (
            .O(N__22096),
            .I(data_in_3_0));
    Odrv4 I__3078 (
            .O(N__22091),
            .I(data_in_3_0));
    LocalMux I__3077 (
            .O(N__22088),
            .I(data_in_3_0));
    InMux I__3076 (
            .O(N__22081),
            .I(N__22078));
    LocalMux I__3075 (
            .O(N__22078),
            .I(N__22074));
    InMux I__3074 (
            .O(N__22077),
            .I(N__22070));
    Span4Mux_h I__3073 (
            .O(N__22074),
            .I(N__22067));
    InMux I__3072 (
            .O(N__22073),
            .I(N__22064));
    LocalMux I__3071 (
            .O(N__22070),
            .I(data_in_0_5));
    Odrv4 I__3070 (
            .O(N__22067),
            .I(data_in_0_5));
    LocalMux I__3069 (
            .O(N__22064),
            .I(data_in_0_5));
    CascadeMux I__3068 (
            .O(N__22057),
            .I(N__22054));
    InMux I__3067 (
            .O(N__22054),
            .I(N__22050));
    InMux I__3066 (
            .O(N__22053),
            .I(N__22045));
    LocalMux I__3065 (
            .O(N__22050),
            .I(N__22042));
    InMux I__3064 (
            .O(N__22049),
            .I(N__22037));
    InMux I__3063 (
            .O(N__22048),
            .I(N__22037));
    LocalMux I__3062 (
            .O(N__22045),
            .I(data_in_3_4));
    Odrv4 I__3061 (
            .O(N__22042),
            .I(data_in_3_4));
    LocalMux I__3060 (
            .O(N__22037),
            .I(data_in_3_4));
    CascadeMux I__3059 (
            .O(N__22030),
            .I(\c0.n9451_cascade_ ));
    CascadeMux I__3058 (
            .O(N__22027),
            .I(n12933_cascade_));
    InMux I__3057 (
            .O(N__22024),
            .I(N__22021));
    LocalMux I__3056 (
            .O(N__22021),
            .I(N__22016));
    InMux I__3055 (
            .O(N__22020),
            .I(N__22010));
    InMux I__3054 (
            .O(N__22019),
            .I(N__22010));
    Span4Mux_h I__3053 (
            .O(N__22016),
            .I(N__22005));
    InMux I__3052 (
            .O(N__22015),
            .I(N__22002));
    LocalMux I__3051 (
            .O(N__22010),
            .I(N__21999));
    InMux I__3050 (
            .O(N__22009),
            .I(N__21994));
    InMux I__3049 (
            .O(N__22008),
            .I(N__21994));
    Odrv4 I__3048 (
            .O(N__22005),
            .I(\c0.n9451 ));
    LocalMux I__3047 (
            .O(N__22002),
            .I(\c0.n9451 ));
    Odrv12 I__3046 (
            .O(N__21999),
            .I(\c0.n9451 ));
    LocalMux I__3045 (
            .O(N__21994),
            .I(\c0.n9451 ));
    InMux I__3044 (
            .O(N__21985),
            .I(N__21982));
    LocalMux I__3043 (
            .O(N__21982),
            .I(N__21979));
    Span4Mux_v I__3042 (
            .O(N__21979),
            .I(N__21976));
    Odrv4 I__3041 (
            .O(N__21976),
            .I(\c0.n9 ));
    InMux I__3040 (
            .O(N__21973),
            .I(N__21970));
    LocalMux I__3039 (
            .O(N__21970),
            .I(\c0.n17258 ));
    CascadeMux I__3038 (
            .O(N__21967),
            .I(\c0.n28_cascade_ ));
    InMux I__3037 (
            .O(N__21964),
            .I(N__21961));
    LocalMux I__3036 (
            .O(N__21961),
            .I(\c0.n60 ));
    InMux I__3035 (
            .O(N__21958),
            .I(N__21955));
    LocalMux I__3034 (
            .O(N__21955),
            .I(\c0.n16879 ));
    InMux I__3033 (
            .O(N__21952),
            .I(N__21949));
    LocalMux I__3032 (
            .O(N__21949),
            .I(N__21945));
    InMux I__3031 (
            .O(N__21948),
            .I(N__21942));
    Span4Mux_v I__3030 (
            .O(N__21945),
            .I(N__21939));
    LocalMux I__3029 (
            .O(N__21942),
            .I(N__21936));
    Span4Mux_h I__3028 (
            .O(N__21939),
            .I(N__21931));
    Span4Mux_h I__3027 (
            .O(N__21936),
            .I(N__21931));
    Odrv4 I__3026 (
            .O(N__21931),
            .I(\c0.n33 ));
    CascadeMux I__3025 (
            .O(N__21928),
            .I(\c0.n16879_cascade_ ));
    CascadeMux I__3024 (
            .O(N__21925),
            .I(N__21922));
    InMux I__3023 (
            .O(N__21922),
            .I(N__21919));
    LocalMux I__3022 (
            .O(N__21919),
            .I(N__21915));
    InMux I__3021 (
            .O(N__21918),
            .I(N__21912));
    Span4Mux_v I__3020 (
            .O(N__21915),
            .I(N__21907));
    LocalMux I__3019 (
            .O(N__21912),
            .I(N__21907));
    Span4Mux_h I__3018 (
            .O(N__21907),
            .I(N__21902));
    InMux I__3017 (
            .O(N__21906),
            .I(N__21899));
    InMux I__3016 (
            .O(N__21905),
            .I(N__21896));
    Span4Mux_s3_h I__3015 (
            .O(N__21902),
            .I(N__21893));
    LocalMux I__3014 (
            .O(N__21899),
            .I(\c0.FRAME_MATCHER_i_6 ));
    LocalMux I__3013 (
            .O(N__21896),
            .I(\c0.FRAME_MATCHER_i_6 ));
    Odrv4 I__3012 (
            .O(N__21893),
            .I(\c0.FRAME_MATCHER_i_6 ));
    CascadeMux I__3011 (
            .O(N__21886),
            .I(N__21881));
    InMux I__3010 (
            .O(N__21885),
            .I(N__21877));
    InMux I__3009 (
            .O(N__21884),
            .I(N__21874));
    InMux I__3008 (
            .O(N__21881),
            .I(N__21871));
    InMux I__3007 (
            .O(N__21880),
            .I(N__21868));
    LocalMux I__3006 (
            .O(N__21877),
            .I(N__21865));
    LocalMux I__3005 (
            .O(N__21874),
            .I(\c0.FRAME_MATCHER_i_7 ));
    LocalMux I__3004 (
            .O(N__21871),
            .I(\c0.FRAME_MATCHER_i_7 ));
    LocalMux I__3003 (
            .O(N__21868),
            .I(\c0.FRAME_MATCHER_i_7 ));
    Odrv4 I__3002 (
            .O(N__21865),
            .I(\c0.FRAME_MATCHER_i_7 ));
    CascadeMux I__3001 (
            .O(N__21856),
            .I(N__21852));
    CascadeMux I__3000 (
            .O(N__21855),
            .I(N__21848));
    InMux I__2999 (
            .O(N__21852),
            .I(N__21842));
    InMux I__2998 (
            .O(N__21851),
            .I(N__21842));
    InMux I__2997 (
            .O(N__21848),
            .I(N__21839));
    CascadeMux I__2996 (
            .O(N__21847),
            .I(N__21836));
    LocalMux I__2995 (
            .O(N__21842),
            .I(N__21831));
    LocalMux I__2994 (
            .O(N__21839),
            .I(N__21831));
    InMux I__2993 (
            .O(N__21836),
            .I(N__21828));
    Span4Mux_v I__2992 (
            .O(N__21831),
            .I(N__21825));
    LocalMux I__2991 (
            .O(N__21828),
            .I(N__21822));
    Span4Mux_h I__2990 (
            .O(N__21825),
            .I(N__21819));
    Span4Mux_h I__2989 (
            .O(N__21822),
            .I(N__21816));
    Odrv4 I__2988 (
            .O(N__21819),
            .I(\c0.FRAME_MATCHER_i_9 ));
    Odrv4 I__2987 (
            .O(N__21816),
            .I(\c0.FRAME_MATCHER_i_9 ));
    InMux I__2986 (
            .O(N__21811),
            .I(N__21807));
    InMux I__2985 (
            .O(N__21810),
            .I(N__21804));
    LocalMux I__2984 (
            .O(N__21807),
            .I(n9445));
    LocalMux I__2983 (
            .O(N__21804),
            .I(n9445));
    CascadeMux I__2982 (
            .O(N__21799),
            .I(N__21796));
    InMux I__2981 (
            .O(N__21796),
            .I(N__21793));
    LocalMux I__2980 (
            .O(N__21793),
            .I(N__21790));
    Odrv4 I__2979 (
            .O(N__21790),
            .I(\c0.n9488 ));
    InMux I__2978 (
            .O(N__21787),
            .I(N__21778));
    InMux I__2977 (
            .O(N__21786),
            .I(N__21778));
    InMux I__2976 (
            .O(N__21785),
            .I(N__21778));
    LocalMux I__2975 (
            .O(N__21778),
            .I(\c0.FRAME_MATCHER_state_5 ));
    InMux I__2974 (
            .O(N__21775),
            .I(N__21771));
    InMux I__2973 (
            .O(N__21774),
            .I(N__21767));
    LocalMux I__2972 (
            .O(N__21771),
            .I(N__21764));
    InMux I__2971 (
            .O(N__21770),
            .I(N__21761));
    LocalMux I__2970 (
            .O(N__21767),
            .I(\c0.FRAME_MATCHER_state_6 ));
    Odrv12 I__2969 (
            .O(N__21764),
            .I(\c0.FRAME_MATCHER_state_6 ));
    LocalMux I__2968 (
            .O(N__21761),
            .I(\c0.FRAME_MATCHER_state_6 ));
    InMux I__2967 (
            .O(N__21754),
            .I(N__21749));
    InMux I__2966 (
            .O(N__21753),
            .I(N__21746));
    InMux I__2965 (
            .O(N__21752),
            .I(N__21743));
    LocalMux I__2964 (
            .O(N__21749),
            .I(N__21738));
    LocalMux I__2963 (
            .O(N__21746),
            .I(N__21738));
    LocalMux I__2962 (
            .O(N__21743),
            .I(\c0.FRAME_MATCHER_state_29 ));
    Odrv12 I__2961 (
            .O(N__21738),
            .I(\c0.FRAME_MATCHER_state_29 ));
    CascadeMux I__2960 (
            .O(N__21733),
            .I(\c0.n59_cascade_ ));
    CascadeMux I__2959 (
            .O(N__21730),
            .I(\c0.n5_adj_2262_cascade_ ));
    CascadeMux I__2958 (
            .O(N__21727),
            .I(\c0.n16876_cascade_ ));
    CascadeMux I__2957 (
            .O(N__21724),
            .I(\c0.n60_cascade_ ));
    SRMux I__2956 (
            .O(N__21721),
            .I(N__21718));
    LocalMux I__2955 (
            .O(N__21718),
            .I(N__21715));
    Odrv4 I__2954 (
            .O(N__21715),
            .I(\c0.n16363 ));
    InMux I__2953 (
            .O(N__21712),
            .I(N__21707));
    InMux I__2952 (
            .O(N__21711),
            .I(N__21704));
    InMux I__2951 (
            .O(N__21710),
            .I(N__21701));
    LocalMux I__2950 (
            .O(N__21707),
            .I(N__21698));
    LocalMux I__2949 (
            .O(N__21704),
            .I(N__21695));
    LocalMux I__2948 (
            .O(N__21701),
            .I(\c0.FRAME_MATCHER_state_30 ));
    Odrv4 I__2947 (
            .O(N__21698),
            .I(\c0.FRAME_MATCHER_state_30 ));
    Odrv12 I__2946 (
            .O(N__21695),
            .I(\c0.FRAME_MATCHER_state_30 ));
    InMux I__2945 (
            .O(N__21688),
            .I(N__21679));
    InMux I__2944 (
            .O(N__21687),
            .I(N__21679));
    InMux I__2943 (
            .O(N__21686),
            .I(N__21679));
    LocalMux I__2942 (
            .O(N__21679),
            .I(\c0.FRAME_MATCHER_state_23 ));
    InMux I__2941 (
            .O(N__21676),
            .I(N__21673));
    LocalMux I__2940 (
            .O(N__21673),
            .I(N__21669));
    InMux I__2939 (
            .O(N__21672),
            .I(N__21666));
    Span4Mux_h I__2938 (
            .O(N__21669),
            .I(N__21663));
    LocalMux I__2937 (
            .O(N__21666),
            .I(n9453));
    Odrv4 I__2936 (
            .O(N__21663),
            .I(n9453));
    CascadeMux I__2935 (
            .O(N__21658),
            .I(N__21654));
    CascadeMux I__2934 (
            .O(N__21657),
            .I(N__21649));
    InMux I__2933 (
            .O(N__21654),
            .I(N__21646));
    InMux I__2932 (
            .O(N__21653),
            .I(N__21643));
    CascadeMux I__2931 (
            .O(N__21652),
            .I(N__21637));
    InMux I__2930 (
            .O(N__21649),
            .I(N__21634));
    LocalMux I__2929 (
            .O(N__21646),
            .I(N__21628));
    LocalMux I__2928 (
            .O(N__21643),
            .I(N__21628));
    InMux I__2927 (
            .O(N__21642),
            .I(N__21625));
    InMux I__2926 (
            .O(N__21641),
            .I(N__21618));
    InMux I__2925 (
            .O(N__21640),
            .I(N__21618));
    InMux I__2924 (
            .O(N__21637),
            .I(N__21618));
    LocalMux I__2923 (
            .O(N__21634),
            .I(N__21615));
    InMux I__2922 (
            .O(N__21633),
            .I(N__21612));
    Span4Mux_v I__2921 (
            .O(N__21628),
            .I(N__21607));
    LocalMux I__2920 (
            .O(N__21625),
            .I(N__21607));
    LocalMux I__2919 (
            .O(N__21618),
            .I(N__21602));
    Span4Mux_v I__2918 (
            .O(N__21615),
            .I(N__21602));
    LocalMux I__2917 (
            .O(N__21612),
            .I(N__21597));
    Span4Mux_v I__2916 (
            .O(N__21607),
            .I(N__21597));
    Span4Mux_h I__2915 (
            .O(N__21602),
            .I(N__21594));
    Span4Mux_h I__2914 (
            .O(N__21597),
            .I(N__21591));
    Span4Mux_s1_h I__2913 (
            .O(N__21594),
            .I(N__21588));
    Odrv4 I__2912 (
            .O(N__21591),
            .I(\c0.FRAME_MATCHER_i_1 ));
    Odrv4 I__2911 (
            .O(N__21588),
            .I(\c0.FRAME_MATCHER_i_1 ));
    InMux I__2910 (
            .O(N__21583),
            .I(N__21579));
    CascadeMux I__2909 (
            .O(N__21582),
            .I(N__21576));
    LocalMux I__2908 (
            .O(N__21579),
            .I(N__21573));
    InMux I__2907 (
            .O(N__21576),
            .I(N__21570));
    Span4Mux_s3_h I__2906 (
            .O(N__21573),
            .I(N__21567));
    LocalMux I__2905 (
            .O(N__21570),
            .I(N__21564));
    Odrv4 I__2904 (
            .O(N__21567),
            .I(n2275));
    Odrv4 I__2903 (
            .O(N__21564),
            .I(n2275));
    CascadeMux I__2902 (
            .O(N__21559),
            .I(n2275_cascade_));
    CascadeMux I__2901 (
            .O(N__21556),
            .I(\c0.n7212_cascade_ ));
    CascadeMux I__2900 (
            .O(N__21553),
            .I(\c0.n17452_cascade_ ));
    InMux I__2899 (
            .O(N__21550),
            .I(N__21547));
    LocalMux I__2898 (
            .O(N__21547),
            .I(\c0.n17454 ));
    CascadeMux I__2897 (
            .O(N__21544),
            .I(\c0.n7_cascade_ ));
    SRMux I__2896 (
            .O(N__21541),
            .I(N__21538));
    LocalMux I__2895 (
            .O(N__21538),
            .I(N__21535));
    Odrv4 I__2894 (
            .O(N__21535),
            .I(\c0.n16335 ));
    SRMux I__2893 (
            .O(N__21532),
            .I(N__21529));
    LocalMux I__2892 (
            .O(N__21529),
            .I(N__21526));
    Span4Mux_h I__2891 (
            .O(N__21526),
            .I(N__21523));
    Odrv4 I__2890 (
            .O(N__21523),
            .I(\c0.n16381 ));
    InMux I__2889 (
            .O(N__21520),
            .I(N__21515));
    CascadeMux I__2888 (
            .O(N__21519),
            .I(N__21511));
    InMux I__2887 (
            .O(N__21518),
            .I(N__21508));
    LocalMux I__2886 (
            .O(N__21515),
            .I(N__21505));
    InMux I__2885 (
            .O(N__21514),
            .I(N__21502));
    InMux I__2884 (
            .O(N__21511),
            .I(N__21499));
    LocalMux I__2883 (
            .O(N__21508),
            .I(N__21496));
    Span4Mux_v I__2882 (
            .O(N__21505),
            .I(N__21493));
    LocalMux I__2881 (
            .O(N__21502),
            .I(N__21488));
    LocalMux I__2880 (
            .O(N__21499),
            .I(N__21488));
    Span4Mux_v I__2879 (
            .O(N__21496),
            .I(N__21485));
    Span4Mux_h I__2878 (
            .O(N__21493),
            .I(N__21480));
    Span4Mux_v I__2877 (
            .O(N__21488),
            .I(N__21480));
    Span4Mux_h I__2876 (
            .O(N__21485),
            .I(N__21477));
    Odrv4 I__2875 (
            .O(N__21480),
            .I(\c0.FRAME_MATCHER_i_19 ));
    Odrv4 I__2874 (
            .O(N__21477),
            .I(\c0.FRAME_MATCHER_i_19 ));
    CascadeMux I__2873 (
            .O(N__21472),
            .I(N__21467));
    InMux I__2872 (
            .O(N__21471),
            .I(N__21463));
    CascadeMux I__2871 (
            .O(N__21470),
            .I(N__21460));
    InMux I__2870 (
            .O(N__21467),
            .I(N__21457));
    InMux I__2869 (
            .O(N__21466),
            .I(N__21454));
    LocalMux I__2868 (
            .O(N__21463),
            .I(N__21451));
    InMux I__2867 (
            .O(N__21460),
            .I(N__21448));
    LocalMux I__2866 (
            .O(N__21457),
            .I(N__21445));
    LocalMux I__2865 (
            .O(N__21454),
            .I(N__21442));
    Span4Mux_v I__2864 (
            .O(N__21451),
            .I(N__21439));
    LocalMux I__2863 (
            .O(N__21448),
            .I(N__21436));
    Span12Mux_s9_v I__2862 (
            .O(N__21445),
            .I(N__21433));
    Span4Mux_v I__2861 (
            .O(N__21442),
            .I(N__21426));
    Span4Mux_v I__2860 (
            .O(N__21439),
            .I(N__21426));
    Span4Mux_h I__2859 (
            .O(N__21436),
            .I(N__21426));
    Odrv12 I__2858 (
            .O(N__21433),
            .I(\c0.FRAME_MATCHER_i_24 ));
    Odrv4 I__2857 (
            .O(N__21426),
            .I(\c0.FRAME_MATCHER_i_24 ));
    InMux I__2856 (
            .O(N__21421),
            .I(N__21418));
    LocalMux I__2855 (
            .O(N__21418),
            .I(N__21415));
    Span4Mux_h I__2854 (
            .O(N__21415),
            .I(N__21412));
    Span4Mux_v I__2853 (
            .O(N__21412),
            .I(N__21409));
    Odrv4 I__2852 (
            .O(N__21409),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_16 ));
    CascadeMux I__2851 (
            .O(N__21406),
            .I(n1716_cascade_));
    InMux I__2850 (
            .O(N__21403),
            .I(N__21400));
    LocalMux I__2849 (
            .O(N__21400),
            .I(n14));
    InMux I__2848 (
            .O(N__21397),
            .I(N__21394));
    LocalMux I__2847 (
            .O(N__21394),
            .I(N__21391));
    Odrv4 I__2846 (
            .O(N__21391),
            .I(n16775));
    InMux I__2845 (
            .O(N__21388),
            .I(N__21384));
    InMux I__2844 (
            .O(N__21387),
            .I(N__21381));
    LocalMux I__2843 (
            .O(N__21384),
            .I(N__21378));
    LocalMux I__2842 (
            .O(N__21381),
            .I(N__21375));
    Span4Mux_h I__2841 (
            .O(N__21378),
            .I(N__21372));
    Odrv4 I__2840 (
            .O(N__21375),
            .I(n3977));
    Odrv4 I__2839 (
            .O(N__21372),
            .I(n3977));
    CascadeMux I__2838 (
            .O(N__21367),
            .I(n16775_cascade_));
    InMux I__2837 (
            .O(N__21364),
            .I(N__21360));
    InMux I__2836 (
            .O(N__21363),
            .I(N__21356));
    LocalMux I__2835 (
            .O(N__21360),
            .I(N__21353));
    InMux I__2834 (
            .O(N__21359),
            .I(N__21350));
    LocalMux I__2833 (
            .O(N__21356),
            .I(\c0.delay_counter_10 ));
    Odrv4 I__2832 (
            .O(N__21353),
            .I(\c0.delay_counter_10 ));
    LocalMux I__2831 (
            .O(N__21350),
            .I(\c0.delay_counter_10 ));
    InMux I__2830 (
            .O(N__21343),
            .I(N__21340));
    LocalMux I__2829 (
            .O(N__21340),
            .I(N__21337));
    Odrv12 I__2828 (
            .O(N__21337),
            .I(\c0.n6522 ));
    InMux I__2827 (
            .O(N__21334),
            .I(\c0.n15523 ));
    InMux I__2826 (
            .O(N__21331),
            .I(N__21328));
    LocalMux I__2825 (
            .O(N__21328),
            .I(N__21323));
    InMux I__2824 (
            .O(N__21327),
            .I(N__21318));
    InMux I__2823 (
            .O(N__21326),
            .I(N__21318));
    Odrv4 I__2822 (
            .O(N__21323),
            .I(\c0.delay_counter_11 ));
    LocalMux I__2821 (
            .O(N__21318),
            .I(\c0.delay_counter_11 ));
    CascadeMux I__2820 (
            .O(N__21313),
            .I(N__21310));
    InMux I__2819 (
            .O(N__21310),
            .I(N__21307));
    LocalMux I__2818 (
            .O(N__21307),
            .I(N__21304));
    Span4Mux_v I__2817 (
            .O(N__21304),
            .I(N__21301));
    Odrv4 I__2816 (
            .O(N__21301),
            .I(\c0.n6521 ));
    InMux I__2815 (
            .O(N__21298),
            .I(\c0.n15524 ));
    CascadeMux I__2814 (
            .O(N__21295),
            .I(N__21292));
    InMux I__2813 (
            .O(N__21292),
            .I(N__21286));
    InMux I__2812 (
            .O(N__21291),
            .I(N__21283));
    CascadeMux I__2811 (
            .O(N__21290),
            .I(N__21280));
    InMux I__2810 (
            .O(N__21289),
            .I(N__21277));
    LocalMux I__2809 (
            .O(N__21286),
            .I(N__21274));
    LocalMux I__2808 (
            .O(N__21283),
            .I(N__21271));
    InMux I__2807 (
            .O(N__21280),
            .I(N__21268));
    LocalMux I__2806 (
            .O(N__21277),
            .I(\c0.delay_counter_12 ));
    Odrv4 I__2805 (
            .O(N__21274),
            .I(\c0.delay_counter_12 ));
    Odrv4 I__2804 (
            .O(N__21271),
            .I(\c0.delay_counter_12 ));
    LocalMux I__2803 (
            .O(N__21268),
            .I(\c0.delay_counter_12 ));
    InMux I__2802 (
            .O(N__21259),
            .I(N__21256));
    LocalMux I__2801 (
            .O(N__21256),
            .I(N__21253));
    Odrv4 I__2800 (
            .O(N__21253),
            .I(\c0.n17575 ));
    InMux I__2799 (
            .O(N__21250),
            .I(\c0.n15525 ));
    InMux I__2798 (
            .O(N__21247),
            .I(N__21244));
    LocalMux I__2797 (
            .O(N__21244),
            .I(N__21241));
    Odrv4 I__2796 (
            .O(N__21241),
            .I(\c0.n17639 ));
    InMux I__2795 (
            .O(N__21238),
            .I(\c0.n15526 ));
    InMux I__2794 (
            .O(N__21235),
            .I(N__21230));
    InMux I__2793 (
            .O(N__21234),
            .I(N__21227));
    InMux I__2792 (
            .O(N__21233),
            .I(N__21224));
    LocalMux I__2791 (
            .O(N__21230),
            .I(N__21221));
    LocalMux I__2790 (
            .O(N__21227),
            .I(N__21217));
    LocalMux I__2789 (
            .O(N__21224),
            .I(N__21212));
    Span4Mux_s2_v I__2788 (
            .O(N__21221),
            .I(N__21212));
    InMux I__2787 (
            .O(N__21220),
            .I(N__21209));
    Odrv4 I__2786 (
            .O(N__21217),
            .I(\c0.delay_counter_14 ));
    Odrv4 I__2785 (
            .O(N__21212),
            .I(\c0.delay_counter_14 ));
    LocalMux I__2784 (
            .O(N__21209),
            .I(\c0.delay_counter_14 ));
    InMux I__2783 (
            .O(N__21202),
            .I(\c0.n15527 ));
    CascadeMux I__2782 (
            .O(N__21199),
            .I(N__21196));
    InMux I__2781 (
            .O(N__21196),
            .I(N__21193));
    LocalMux I__2780 (
            .O(N__21193),
            .I(N__21190));
    Odrv4 I__2779 (
            .O(N__21190),
            .I(\c0.n17635 ));
    SRMux I__2778 (
            .O(N__21187),
            .I(N__21184));
    LocalMux I__2777 (
            .O(N__21184),
            .I(N__21181));
    Odrv4 I__2776 (
            .O(N__21181),
            .I(\c0.n16331 ));
    InMux I__2775 (
            .O(N__21178),
            .I(N__21175));
    LocalMux I__2774 (
            .O(N__21175),
            .I(\c0.n6530 ));
    InMux I__2773 (
            .O(N__21172),
            .I(\c0.n15515 ));
    InMux I__2772 (
            .O(N__21169),
            .I(N__21164));
    InMux I__2771 (
            .O(N__21168),
            .I(N__21159));
    InMux I__2770 (
            .O(N__21167),
            .I(N__21159));
    LocalMux I__2769 (
            .O(N__21164),
            .I(\c0.delay_counter_3 ));
    LocalMux I__2768 (
            .O(N__21159),
            .I(\c0.delay_counter_3 ));
    CascadeMux I__2767 (
            .O(N__21154),
            .I(N__21151));
    InMux I__2766 (
            .O(N__21151),
            .I(N__21148));
    LocalMux I__2765 (
            .O(N__21148),
            .I(\c0.n6529 ));
    InMux I__2764 (
            .O(N__21145),
            .I(\c0.n15516 ));
    CascadeMux I__2763 (
            .O(N__21142),
            .I(N__21139));
    InMux I__2762 (
            .O(N__21139),
            .I(N__21136));
    LocalMux I__2761 (
            .O(N__21136),
            .I(\c0.n6528 ));
    InMux I__2760 (
            .O(N__21133),
            .I(\c0.n15517 ));
    InMux I__2759 (
            .O(N__21130),
            .I(N__21124));
    InMux I__2758 (
            .O(N__21129),
            .I(N__21121));
    InMux I__2757 (
            .O(N__21128),
            .I(N__21118));
    InMux I__2756 (
            .O(N__21127),
            .I(N__21115));
    LocalMux I__2755 (
            .O(N__21124),
            .I(\c0.delay_counter_5 ));
    LocalMux I__2754 (
            .O(N__21121),
            .I(\c0.delay_counter_5 ));
    LocalMux I__2753 (
            .O(N__21118),
            .I(\c0.delay_counter_5 ));
    LocalMux I__2752 (
            .O(N__21115),
            .I(\c0.delay_counter_5 ));
    InMux I__2751 (
            .O(N__21106),
            .I(N__21103));
    LocalMux I__2750 (
            .O(N__21103),
            .I(\c0.n17574 ));
    InMux I__2749 (
            .O(N__21100),
            .I(\c0.n15518 ));
    InMux I__2748 (
            .O(N__21097),
            .I(N__21092));
    InMux I__2747 (
            .O(N__21096),
            .I(N__21089));
    InMux I__2746 (
            .O(N__21095),
            .I(N__21086));
    LocalMux I__2745 (
            .O(N__21092),
            .I(N__21083));
    LocalMux I__2744 (
            .O(N__21089),
            .I(\c0.delay_counter_6 ));
    LocalMux I__2743 (
            .O(N__21086),
            .I(\c0.delay_counter_6 ));
    Odrv4 I__2742 (
            .O(N__21083),
            .I(\c0.delay_counter_6 ));
    InMux I__2741 (
            .O(N__21076),
            .I(N__21073));
    LocalMux I__2740 (
            .O(N__21073),
            .I(\c0.n6526 ));
    InMux I__2739 (
            .O(N__21070),
            .I(\c0.n15519 ));
    InMux I__2738 (
            .O(N__21067),
            .I(N__21061));
    InMux I__2737 (
            .O(N__21066),
            .I(N__21058));
    InMux I__2736 (
            .O(N__21065),
            .I(N__21055));
    InMux I__2735 (
            .O(N__21064),
            .I(N__21052));
    LocalMux I__2734 (
            .O(N__21061),
            .I(\c0.delay_counter_7 ));
    LocalMux I__2733 (
            .O(N__21058),
            .I(\c0.delay_counter_7 ));
    LocalMux I__2732 (
            .O(N__21055),
            .I(\c0.delay_counter_7 ));
    LocalMux I__2731 (
            .O(N__21052),
            .I(\c0.delay_counter_7 ));
    InMux I__2730 (
            .O(N__21043),
            .I(N__21040));
    LocalMux I__2729 (
            .O(N__21040),
            .I(\c0.n17638 ));
    InMux I__2728 (
            .O(N__21037),
            .I(\c0.n15520 ));
    CascadeMux I__2727 (
            .O(N__21034),
            .I(N__21031));
    InMux I__2726 (
            .O(N__21031),
            .I(N__21028));
    LocalMux I__2725 (
            .O(N__21028),
            .I(N__21025));
    Odrv4 I__2724 (
            .O(N__21025),
            .I(\c0.n6524 ));
    InMux I__2723 (
            .O(N__21022),
            .I(bfn_5_32_0_));
    InMux I__2722 (
            .O(N__21019),
            .I(N__21014));
    InMux I__2721 (
            .O(N__21018),
            .I(N__21011));
    InMux I__2720 (
            .O(N__21017),
            .I(N__21008));
    LocalMux I__2719 (
            .O(N__21014),
            .I(\c0.delay_counter_9 ));
    LocalMux I__2718 (
            .O(N__21011),
            .I(\c0.delay_counter_9 ));
    LocalMux I__2717 (
            .O(N__21008),
            .I(\c0.delay_counter_9 ));
    InMux I__2716 (
            .O(N__21001),
            .I(N__20998));
    LocalMux I__2715 (
            .O(N__20998),
            .I(\c0.n6523 ));
    InMux I__2714 (
            .O(N__20995),
            .I(\c0.n15522 ));
    CascadeMux I__2713 (
            .O(N__20992),
            .I(\c0.n1419_cascade_ ));
    InMux I__2712 (
            .O(N__20989),
            .I(N__20971));
    InMux I__2711 (
            .O(N__20988),
            .I(N__20971));
    InMux I__2710 (
            .O(N__20987),
            .I(N__20964));
    InMux I__2709 (
            .O(N__20986),
            .I(N__20964));
    InMux I__2708 (
            .O(N__20985),
            .I(N__20964));
    InMux I__2707 (
            .O(N__20984),
            .I(N__20957));
    InMux I__2706 (
            .O(N__20983),
            .I(N__20957));
    InMux I__2705 (
            .O(N__20982),
            .I(N__20957));
    InMux I__2704 (
            .O(N__20981),
            .I(N__20944));
    InMux I__2703 (
            .O(N__20980),
            .I(N__20944));
    InMux I__2702 (
            .O(N__20979),
            .I(N__20944));
    InMux I__2701 (
            .O(N__20978),
            .I(N__20944));
    InMux I__2700 (
            .O(N__20977),
            .I(N__20944));
    InMux I__2699 (
            .O(N__20976),
            .I(N__20944));
    LocalMux I__2698 (
            .O(N__20971),
            .I(\c0.n1419 ));
    LocalMux I__2697 (
            .O(N__20964),
            .I(\c0.n1419 ));
    LocalMux I__2696 (
            .O(N__20957),
            .I(\c0.n1419 ));
    LocalMux I__2695 (
            .O(N__20944),
            .I(\c0.n1419 ));
    InMux I__2694 (
            .O(N__20935),
            .I(N__20932));
    LocalMux I__2693 (
            .O(N__20932),
            .I(n53));
    InMux I__2692 (
            .O(N__20929),
            .I(N__20925));
    InMux I__2691 (
            .O(N__20928),
            .I(N__20920));
    LocalMux I__2690 (
            .O(N__20925),
            .I(N__20917));
    InMux I__2689 (
            .O(N__20924),
            .I(N__20914));
    CascadeMux I__2688 (
            .O(N__20923),
            .I(N__20911));
    LocalMux I__2687 (
            .O(N__20920),
            .I(N__20906));
    Span4Mux_s3_v I__2686 (
            .O(N__20917),
            .I(N__20906));
    LocalMux I__2685 (
            .O(N__20914),
            .I(N__20903));
    InMux I__2684 (
            .O(N__20911),
            .I(N__20900));
    Odrv4 I__2683 (
            .O(N__20906),
            .I(\c0.delay_counter_0 ));
    Odrv4 I__2682 (
            .O(N__20903),
            .I(\c0.delay_counter_0 ));
    LocalMux I__2681 (
            .O(N__20900),
            .I(\c0.delay_counter_0 ));
    InMux I__2680 (
            .O(N__20893),
            .I(N__20890));
    LocalMux I__2679 (
            .O(N__20890),
            .I(N__20887));
    Odrv4 I__2678 (
            .O(N__20887),
            .I(\c0.n17637 ));
    InMux I__2677 (
            .O(N__20884),
            .I(bfn_5_31_0_));
    CascadeMux I__2676 (
            .O(N__20881),
            .I(N__20878));
    InMux I__2675 (
            .O(N__20878),
            .I(N__20873));
    InMux I__2674 (
            .O(N__20877),
            .I(N__20870));
    InMux I__2673 (
            .O(N__20876),
            .I(N__20867));
    LocalMux I__2672 (
            .O(N__20873),
            .I(\c0.delay_counter_1 ));
    LocalMux I__2671 (
            .O(N__20870),
            .I(\c0.delay_counter_1 ));
    LocalMux I__2670 (
            .O(N__20867),
            .I(\c0.delay_counter_1 ));
    InMux I__2669 (
            .O(N__20860),
            .I(N__20857));
    LocalMux I__2668 (
            .O(N__20857),
            .I(\c0.n6531 ));
    InMux I__2667 (
            .O(N__20854),
            .I(\c0.n15514 ));
    InMux I__2666 (
            .O(N__20851),
            .I(N__20842));
    InMux I__2665 (
            .O(N__20850),
            .I(N__20839));
    InMux I__2664 (
            .O(N__20849),
            .I(N__20830));
    InMux I__2663 (
            .O(N__20848),
            .I(N__20830));
    InMux I__2662 (
            .O(N__20847),
            .I(N__20830));
    InMux I__2661 (
            .O(N__20846),
            .I(N__20830));
    InMux I__2660 (
            .O(N__20845),
            .I(N__20827));
    LocalMux I__2659 (
            .O(N__20842),
            .I(n16893));
    LocalMux I__2658 (
            .O(N__20839),
            .I(n16893));
    LocalMux I__2657 (
            .O(N__20830),
            .I(n16893));
    LocalMux I__2656 (
            .O(N__20827),
            .I(n16893));
    InMux I__2655 (
            .O(N__20818),
            .I(N__20815));
    LocalMux I__2654 (
            .O(N__20815),
            .I(\c0.tx.n17462 ));
    InMux I__2653 (
            .O(N__20812),
            .I(N__20805));
    InMux I__2652 (
            .O(N__20811),
            .I(N__20802));
    InMux I__2651 (
            .O(N__20810),
            .I(N__20799));
    InMux I__2650 (
            .O(N__20809),
            .I(N__20796));
    InMux I__2649 (
            .O(N__20808),
            .I(N__20793));
    LocalMux I__2648 (
            .O(N__20805),
            .I(N__20790));
    LocalMux I__2647 (
            .O(N__20802),
            .I(N__20783));
    LocalMux I__2646 (
            .O(N__20799),
            .I(N__20783));
    LocalMux I__2645 (
            .O(N__20796),
            .I(N__20783));
    LocalMux I__2644 (
            .O(N__20793),
            .I(\c0.tx.r_Bit_Index_0 ));
    Odrv12 I__2643 (
            .O(N__20790),
            .I(\c0.tx.r_Bit_Index_0 ));
    Odrv4 I__2642 (
            .O(N__20783),
            .I(\c0.tx.r_Bit_Index_0 ));
    InMux I__2641 (
            .O(N__20776),
            .I(N__20773));
    LocalMux I__2640 (
            .O(N__20773),
            .I(N__20770));
    Span4Mux_h I__2639 (
            .O(N__20770),
            .I(N__20767));
    Odrv4 I__2638 (
            .O(N__20767),
            .I(n17397));
    CascadeMux I__2637 (
            .O(N__20764),
            .I(N__20758));
    InMux I__2636 (
            .O(N__20763),
            .I(N__20755));
    InMux I__2635 (
            .O(N__20762),
            .I(N__20750));
    InMux I__2634 (
            .O(N__20761),
            .I(N__20750));
    InMux I__2633 (
            .O(N__20758),
            .I(N__20747));
    LocalMux I__2632 (
            .O(N__20755),
            .I(\c0.tx.r_Bit_Index_2 ));
    LocalMux I__2631 (
            .O(N__20750),
            .I(\c0.tx.r_Bit_Index_2 ));
    LocalMux I__2630 (
            .O(N__20747),
            .I(\c0.tx.r_Bit_Index_2 ));
    CascadeMux I__2629 (
            .O(N__20740),
            .I(\c0.tx.n17975_cascade_ ));
    CascadeMux I__2628 (
            .O(N__20737),
            .I(\c0.tx.o_Tx_Serial_N_2064_cascade_ ));
    InMux I__2627 (
            .O(N__20734),
            .I(N__20731));
    LocalMux I__2626 (
            .O(N__20731),
            .I(N__20728));
    Odrv4 I__2625 (
            .O(N__20728),
            .I(n3_adj_2406));
    InMux I__2624 (
            .O(N__20725),
            .I(N__20722));
    LocalMux I__2623 (
            .O(N__20722),
            .I(N__20719));
    Span4Mux_h I__2622 (
            .O(N__20719),
            .I(N__20715));
    InMux I__2621 (
            .O(N__20718),
            .I(N__20712));
    Span4Mux_v I__2620 (
            .O(N__20715),
            .I(N__20709));
    LocalMux I__2619 (
            .O(N__20712),
            .I(N__20706));
    Odrv4 I__2618 (
            .O(N__20709),
            .I(n13082));
    Odrv4 I__2617 (
            .O(N__20706),
            .I(n13082));
    CascadeMux I__2616 (
            .O(N__20701),
            .I(\c0.n16891_cascade_ ));
    InMux I__2615 (
            .O(N__20698),
            .I(N__20694));
    InMux I__2614 (
            .O(N__20697),
            .I(N__20690));
    LocalMux I__2613 (
            .O(N__20694),
            .I(N__20687));
    InMux I__2612 (
            .O(N__20693),
            .I(N__20682));
    LocalMux I__2611 (
            .O(N__20690),
            .I(N__20679));
    Span4Mux_v I__2610 (
            .O(N__20687),
            .I(N__20676));
    InMux I__2609 (
            .O(N__20686),
            .I(N__20671));
    InMux I__2608 (
            .O(N__20685),
            .I(N__20671));
    LocalMux I__2607 (
            .O(N__20682),
            .I(r_Bit_Index_0));
    Odrv12 I__2606 (
            .O(N__20679),
            .I(r_Bit_Index_0));
    Odrv4 I__2605 (
            .O(N__20676),
            .I(r_Bit_Index_0));
    LocalMux I__2604 (
            .O(N__20671),
            .I(r_Bit_Index_0));
    InMux I__2603 (
            .O(N__20662),
            .I(N__20659));
    LocalMux I__2602 (
            .O(N__20659),
            .I(N__20655));
    InMux I__2601 (
            .O(N__20658),
            .I(N__20652));
    Odrv4 I__2600 (
            .O(N__20655),
            .I(\c0.rx.n9323 ));
    LocalMux I__2599 (
            .O(N__20652),
            .I(\c0.rx.n9323 ));
    InMux I__2598 (
            .O(N__20647),
            .I(N__20641));
    InMux I__2597 (
            .O(N__20646),
            .I(N__20641));
    LocalMux I__2596 (
            .O(N__20641),
            .I(N__20637));
    InMux I__2595 (
            .O(N__20640),
            .I(N__20634));
    Odrv12 I__2594 (
            .O(N__20637),
            .I(n9477));
    LocalMux I__2593 (
            .O(N__20634),
            .I(n9477));
    InMux I__2592 (
            .O(N__20629),
            .I(N__20626));
    LocalMux I__2591 (
            .O(N__20626),
            .I(N__20622));
    InMux I__2590 (
            .O(N__20625),
            .I(N__20619));
    Odrv4 I__2589 (
            .O(N__20622),
            .I(n4_adj_2409));
    LocalMux I__2588 (
            .O(N__20619),
            .I(n4_adj_2409));
    CascadeMux I__2587 (
            .O(N__20614),
            .I(n9477_cascade_));
    InMux I__2586 (
            .O(N__20611),
            .I(N__20607));
    InMux I__2585 (
            .O(N__20610),
            .I(N__20604));
    LocalMux I__2584 (
            .O(N__20607),
            .I(data_in_0_2));
    LocalMux I__2583 (
            .O(N__20604),
            .I(data_in_0_2));
    InMux I__2582 (
            .O(N__20599),
            .I(N__20596));
    LocalMux I__2581 (
            .O(N__20596),
            .I(N__20591));
    InMux I__2580 (
            .O(N__20595),
            .I(N__20586));
    InMux I__2579 (
            .O(N__20594),
            .I(N__20586));
    Odrv4 I__2578 (
            .O(N__20591),
            .I(data_in_1_3));
    LocalMux I__2577 (
            .O(N__20586),
            .I(data_in_1_3));
    InMux I__2576 (
            .O(N__20581),
            .I(N__20578));
    LocalMux I__2575 (
            .O(N__20578),
            .I(N__20575));
    Odrv4 I__2574 (
            .O(N__20575),
            .I(\c0.n12_adj_2200 ));
    CascadeMux I__2573 (
            .O(N__20572),
            .I(N__20569));
    InMux I__2572 (
            .O(N__20569),
            .I(N__20566));
    LocalMux I__2571 (
            .O(N__20566),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_31 ));
    InMux I__2570 (
            .O(N__20563),
            .I(N__20559));
    InMux I__2569 (
            .O(N__20562),
            .I(N__20556));
    LocalMux I__2568 (
            .O(N__20559),
            .I(N__20553));
    LocalMux I__2567 (
            .O(N__20556),
            .I(N__20550));
    Span4Mux_h I__2566 (
            .O(N__20553),
            .I(N__20547));
    Span4Mux_h I__2565 (
            .O(N__20550),
            .I(N__20544));
    Odrv4 I__2564 (
            .O(N__20547),
            .I(n4_adj_2460));
    Odrv4 I__2563 (
            .O(N__20544),
            .I(n4_adj_2460));
    InMux I__2562 (
            .O(N__20539),
            .I(N__20536));
    LocalMux I__2561 (
            .O(N__20536),
            .I(N__20532));
    InMux I__2560 (
            .O(N__20535),
            .I(N__20529));
    Span4Mux_h I__2559 (
            .O(N__20532),
            .I(N__20524));
    LocalMux I__2558 (
            .O(N__20529),
            .I(N__20524));
    Odrv4 I__2557 (
            .O(N__20524),
            .I(n4_adj_2417));
    CascadeMux I__2556 (
            .O(N__20521),
            .I(\c0.n127_adj_2136_cascade_ ));
    InMux I__2555 (
            .O(N__20518),
            .I(N__20515));
    LocalMux I__2554 (
            .O(N__20515),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_27 ));
    InMux I__2553 (
            .O(N__20512),
            .I(N__20509));
    LocalMux I__2552 (
            .O(N__20509),
            .I(N__20504));
    InMux I__2551 (
            .O(N__20508),
            .I(N__20499));
    InMux I__2550 (
            .O(N__20507),
            .I(N__20499));
    Span4Mux_v I__2549 (
            .O(N__20504),
            .I(N__20496));
    LocalMux I__2548 (
            .O(N__20499),
            .I(N__20493));
    Odrv4 I__2547 (
            .O(N__20496),
            .I(n9472));
    Odrv4 I__2546 (
            .O(N__20493),
            .I(n9472));
    InMux I__2545 (
            .O(N__20488),
            .I(N__20485));
    LocalMux I__2544 (
            .O(N__20485),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_30 ));
    InMux I__2543 (
            .O(N__20482),
            .I(N__20479));
    LocalMux I__2542 (
            .O(N__20479),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_25 ));
    InMux I__2541 (
            .O(N__20476),
            .I(N__20473));
    LocalMux I__2540 (
            .O(N__20473),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_28 ));
    InMux I__2539 (
            .O(N__20470),
            .I(N__20467));
    LocalMux I__2538 (
            .O(N__20467),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_24 ));
    InMux I__2537 (
            .O(N__20464),
            .I(N__20461));
    LocalMux I__2536 (
            .O(N__20461),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_26 ));
    InMux I__2535 (
            .O(N__20458),
            .I(N__20455));
    LocalMux I__2534 (
            .O(N__20455),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_22 ));
    InMux I__2533 (
            .O(N__20452),
            .I(N__20449));
    LocalMux I__2532 (
            .O(N__20449),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_9 ));
    SRMux I__2531 (
            .O(N__20446),
            .I(N__20443));
    LocalMux I__2530 (
            .O(N__20443),
            .I(N__20440));
    Span4Mux_h I__2529 (
            .O(N__20440),
            .I(N__20437));
    Odrv4 I__2528 (
            .O(N__20437),
            .I(\c0.n3_adj_2248 ));
    InMux I__2527 (
            .O(N__20434),
            .I(N__20431));
    LocalMux I__2526 (
            .O(N__20431),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_8 ));
    InMux I__2525 (
            .O(N__20428),
            .I(N__20425));
    LocalMux I__2524 (
            .O(N__20425),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_19 ));
    InMux I__2523 (
            .O(N__20422),
            .I(N__20419));
    LocalMux I__2522 (
            .O(N__20419),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_20 ));
    InMux I__2521 (
            .O(N__20416),
            .I(N__20413));
    LocalMux I__2520 (
            .O(N__20413),
            .I(N__20410));
    Odrv4 I__2519 (
            .O(N__20410),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_21 ));
    InMux I__2518 (
            .O(N__20407),
            .I(N__20404));
    LocalMux I__2517 (
            .O(N__20404),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_23 ));
    CascadeMux I__2516 (
            .O(N__20401),
            .I(\c0.n18_adj_2198_cascade_ ));
    InMux I__2515 (
            .O(N__20398),
            .I(N__20395));
    LocalMux I__2514 (
            .O(N__20395),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_6 ));
    SRMux I__2513 (
            .O(N__20392),
            .I(N__20389));
    LocalMux I__2512 (
            .O(N__20389),
            .I(\c0.n3_adj_2253 ));
    SRMux I__2511 (
            .O(N__20386),
            .I(N__20383));
    LocalMux I__2510 (
            .O(N__20383),
            .I(N__20380));
    Span4Mux_h I__2509 (
            .O(N__20380),
            .I(N__20377));
    Odrv4 I__2508 (
            .O(N__20377),
            .I(\c0.n3_adj_2237 ));
    SRMux I__2507 (
            .O(N__20374),
            .I(N__20371));
    LocalMux I__2506 (
            .O(N__20371),
            .I(N__20368));
    Span4Mux_s1_h I__2505 (
            .O(N__20368),
            .I(N__20365));
    Span4Mux_v I__2504 (
            .O(N__20365),
            .I(N__20362));
    Odrv4 I__2503 (
            .O(N__20362),
            .I(\c0.n3_adj_2235 ));
    InMux I__2502 (
            .O(N__20359),
            .I(N__20356));
    LocalMux I__2501 (
            .O(N__20356),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_11 ));
    InMux I__2500 (
            .O(N__20353),
            .I(N__20350));
    LocalMux I__2499 (
            .O(N__20350),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_11 ));
    SRMux I__2498 (
            .O(N__20347),
            .I(N__20344));
    LocalMux I__2497 (
            .O(N__20344),
            .I(N__20341));
    Odrv4 I__2496 (
            .O(N__20341),
            .I(\c0.n3_adj_2246 ));
    InMux I__2495 (
            .O(N__20338),
            .I(N__20335));
    LocalMux I__2494 (
            .O(N__20335),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_10 ));
    SRMux I__2493 (
            .O(N__20332),
            .I(N__20329));
    LocalMux I__2492 (
            .O(N__20329),
            .I(N__20326));
    Span4Mux_v I__2491 (
            .O(N__20326),
            .I(N__20323));
    Span4Mux_s1_h I__2490 (
            .O(N__20323),
            .I(N__20320));
    Odrv4 I__2489 (
            .O(N__20320),
            .I(\c0.n3_adj_2231 ));
    SRMux I__2488 (
            .O(N__20317),
            .I(N__20314));
    LocalMux I__2487 (
            .O(N__20314),
            .I(N__20311));
    Span4Mux_h I__2486 (
            .O(N__20311),
            .I(N__20308));
    Span4Mux_v I__2485 (
            .O(N__20308),
            .I(N__20305));
    Odrv4 I__2484 (
            .O(N__20305),
            .I(\c0.n3_adj_2227 ));
    SRMux I__2483 (
            .O(N__20302),
            .I(N__20299));
    LocalMux I__2482 (
            .O(N__20299),
            .I(N__20296));
    Span4Mux_v I__2481 (
            .O(N__20296),
            .I(N__20293));
    Odrv4 I__2480 (
            .O(N__20293),
            .I(\c0.n3_adj_2223 ));
    SRMux I__2479 (
            .O(N__20290),
            .I(N__20287));
    LocalMux I__2478 (
            .O(N__20287),
            .I(N__20284));
    Span4Mux_v I__2477 (
            .O(N__20284),
            .I(N__20281));
    Span4Mux_s2_h I__2476 (
            .O(N__20281),
            .I(N__20278));
    Odrv4 I__2475 (
            .O(N__20278),
            .I(\c0.n3_adj_2225 ));
    CascadeMux I__2474 (
            .O(N__20275),
            .I(\c0.n1439_cascade_ ));
    SRMux I__2473 (
            .O(N__20272),
            .I(N__20269));
    LocalMux I__2472 (
            .O(N__20269),
            .I(N__20266));
    Span4Mux_v I__2471 (
            .O(N__20266),
            .I(N__20263));
    Span4Mux_h I__2470 (
            .O(N__20263),
            .I(N__20260));
    Odrv4 I__2469 (
            .O(N__20260),
            .I(\c0.n3_adj_2221 ));
    InMux I__2468 (
            .O(N__20257),
            .I(N__20254));
    LocalMux I__2467 (
            .O(N__20254),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_7 ));
    InMux I__2466 (
            .O(N__20251),
            .I(N__20248));
    LocalMux I__2465 (
            .O(N__20248),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_7 ));
    SRMux I__2464 (
            .O(N__20245),
            .I(N__20242));
    LocalMux I__2463 (
            .O(N__20242),
            .I(N__20239));
    Odrv4 I__2462 (
            .O(N__20239),
            .I(\c0.n3_adj_2250 ));
    CascadeMux I__2461 (
            .O(N__20236),
            .I(n3977_cascade_));
    SRMux I__2460 (
            .O(N__20233),
            .I(N__20230));
    LocalMux I__2459 (
            .O(N__20230),
            .I(\c0.n3_adj_2233 ));
    SRMux I__2458 (
            .O(N__20227),
            .I(N__20224));
    LocalMux I__2457 (
            .O(N__20224),
            .I(N__20221));
    Odrv4 I__2456 (
            .O(N__20221),
            .I(\c0.n3_adj_2219 ));
    SRMux I__2455 (
            .O(N__20218),
            .I(N__20215));
    LocalMux I__2454 (
            .O(N__20215),
            .I(N__20212));
    Span4Mux_h I__2453 (
            .O(N__20212),
            .I(N__20209));
    Odrv4 I__2452 (
            .O(N__20209),
            .I(\c0.n16441 ));
    SRMux I__2451 (
            .O(N__20206),
            .I(N__20203));
    LocalMux I__2450 (
            .O(N__20203),
            .I(N__20200));
    Span4Mux_s2_h I__2449 (
            .O(N__20200),
            .I(N__20197));
    Odrv4 I__2448 (
            .O(N__20197),
            .I(\c0.n3_adj_2229 ));
    CascadeMux I__2447 (
            .O(N__20194),
            .I(n29_cascade_));
    IoInMux I__2446 (
            .O(N__20191),
            .I(N__20188));
    LocalMux I__2445 (
            .O(N__20188),
            .I(tx_enable));
    CascadeMux I__2444 (
            .O(N__20185),
            .I(N__20182));
    InMux I__2443 (
            .O(N__20182),
            .I(N__20179));
    LocalMux I__2442 (
            .O(N__20179),
            .I(\c0.n12991 ));
    CascadeMux I__2441 (
            .O(N__20176),
            .I(\c0.n12991_cascade_ ));
    InMux I__2440 (
            .O(N__20173),
            .I(N__20170));
    LocalMux I__2439 (
            .O(N__20170),
            .I(\c0.n19_adj_2270 ));
    InMux I__2438 (
            .O(N__20167),
            .I(N__20164));
    LocalMux I__2437 (
            .O(N__20164),
            .I(N__20161));
    Odrv4 I__2436 (
            .O(N__20161),
            .I(n16859));
    InMux I__2435 (
            .O(N__20158),
            .I(N__20155));
    LocalMux I__2434 (
            .O(N__20155),
            .I(N__20151));
    InMux I__2433 (
            .O(N__20154),
            .I(N__20148));
    Span4Mux_v I__2432 (
            .O(N__20151),
            .I(N__20142));
    LocalMux I__2431 (
            .O(N__20148),
            .I(N__20142));
    InMux I__2430 (
            .O(N__20147),
            .I(N__20134));
    Span4Mux_s2_v I__2429 (
            .O(N__20142),
            .I(N__20131));
    InMux I__2428 (
            .O(N__20141),
            .I(N__20126));
    InMux I__2427 (
            .O(N__20140),
            .I(N__20126));
    InMux I__2426 (
            .O(N__20139),
            .I(N__20123));
    InMux I__2425 (
            .O(N__20138),
            .I(N__20120));
    InMux I__2424 (
            .O(N__20137),
            .I(N__20117));
    LocalMux I__2423 (
            .O(N__20134),
            .I(N__20114));
    Odrv4 I__2422 (
            .O(N__20131),
            .I(n17_adj_2416));
    LocalMux I__2421 (
            .O(N__20126),
            .I(n17_adj_2416));
    LocalMux I__2420 (
            .O(N__20123),
            .I(n17_adj_2416));
    LocalMux I__2419 (
            .O(N__20120),
            .I(n17_adj_2416));
    LocalMux I__2418 (
            .O(N__20117),
            .I(n17_adj_2416));
    Odrv4 I__2417 (
            .O(N__20114),
            .I(n17_adj_2416));
    InMux I__2416 (
            .O(N__20101),
            .I(N__20097));
    InMux I__2415 (
            .O(N__20100),
            .I(N__20093));
    LocalMux I__2414 (
            .O(N__20097),
            .I(N__20090));
    InMux I__2413 (
            .O(N__20096),
            .I(N__20087));
    LocalMux I__2412 (
            .O(N__20093),
            .I(N__20084));
    Span4Mux_s3_h I__2411 (
            .O(N__20090),
            .I(N__20081));
    LocalMux I__2410 (
            .O(N__20087),
            .I(r_Clock_Count_0_adj_2437));
    Odrv4 I__2409 (
            .O(N__20084),
            .I(r_Clock_Count_0_adj_2437));
    Odrv4 I__2408 (
            .O(N__20081),
            .I(r_Clock_Count_0_adj_2437));
    IoInMux I__2407 (
            .O(N__20074),
            .I(N__20069));
    InMux I__2406 (
            .O(N__20073),
            .I(N__20064));
    InMux I__2405 (
            .O(N__20072),
            .I(N__20064));
    LocalMux I__2404 (
            .O(N__20069),
            .I(tx_o));
    LocalMux I__2403 (
            .O(N__20064),
            .I(tx_o));
    InMux I__2402 (
            .O(N__20059),
            .I(N__20056));
    LocalMux I__2401 (
            .O(N__20056),
            .I(N__20053));
    Span4Mux_h I__2400 (
            .O(N__20053),
            .I(N__20049));
    InMux I__2399 (
            .O(N__20052),
            .I(N__20045));
    Sp12to4 I__2398 (
            .O(N__20049),
            .I(N__20042));
    InMux I__2397 (
            .O(N__20048),
            .I(N__20039));
    LocalMux I__2396 (
            .O(N__20045),
            .I(data_in_1_0));
    Odrv12 I__2395 (
            .O(N__20042),
            .I(data_in_1_0));
    LocalMux I__2394 (
            .O(N__20039),
            .I(data_in_1_0));
    InMux I__2393 (
            .O(N__20032),
            .I(N__20029));
    LocalMux I__2392 (
            .O(N__20029),
            .I(\c0.n12993 ));
    InMux I__2391 (
            .O(N__20026),
            .I(N__20022));
    InMux I__2390 (
            .O(N__20025),
            .I(N__20019));
    LocalMux I__2389 (
            .O(N__20022),
            .I(\c0.n13298 ));
    LocalMux I__2388 (
            .O(N__20019),
            .I(\c0.n13298 ));
    InMux I__2387 (
            .O(N__20014),
            .I(N__20011));
    LocalMux I__2386 (
            .O(N__20011),
            .I(\c0.n20_adj_2267 ));
    CascadeMux I__2385 (
            .O(N__20008),
            .I(\c0.n21_adj_2271_cascade_ ));
    InMux I__2384 (
            .O(N__20005),
            .I(N__19998));
    InMux I__2383 (
            .O(N__20004),
            .I(N__19995));
    InMux I__2382 (
            .O(N__20003),
            .I(N__19990));
    InMux I__2381 (
            .O(N__20002),
            .I(N__19990));
    InMux I__2380 (
            .O(N__20001),
            .I(N__19987));
    LocalMux I__2379 (
            .O(N__19998),
            .I(N__19984));
    LocalMux I__2378 (
            .O(N__19995),
            .I(r_SM_Main_2_N_2033_1));
    LocalMux I__2377 (
            .O(N__19990),
            .I(r_SM_Main_2_N_2033_1));
    LocalMux I__2376 (
            .O(N__19987),
            .I(r_SM_Main_2_N_2033_1));
    Odrv4 I__2375 (
            .O(N__19984),
            .I(r_SM_Main_2_N_2033_1));
    InMux I__2374 (
            .O(N__19975),
            .I(N__19972));
    LocalMux I__2373 (
            .O(N__19972),
            .I(N__19966));
    InMux I__2372 (
            .O(N__19971),
            .I(N__19963));
    CascadeMux I__2371 (
            .O(N__19970),
            .I(N__19958));
    CascadeMux I__2370 (
            .O(N__19969),
            .I(N__19954));
    Sp12to4 I__2369 (
            .O(N__19966),
            .I(N__19949));
    LocalMux I__2368 (
            .O(N__19963),
            .I(N__19949));
    InMux I__2367 (
            .O(N__19962),
            .I(N__19946));
    InMux I__2366 (
            .O(N__19961),
            .I(N__19941));
    InMux I__2365 (
            .O(N__19958),
            .I(N__19941));
    InMux I__2364 (
            .O(N__19957),
            .I(N__19936));
    InMux I__2363 (
            .O(N__19954),
            .I(N__19936));
    Odrv12 I__2362 (
            .O(N__19949),
            .I(r_Bit_Index_2));
    LocalMux I__2361 (
            .O(N__19946),
            .I(r_Bit_Index_2));
    LocalMux I__2360 (
            .O(N__19941),
            .I(r_Bit_Index_2));
    LocalMux I__2359 (
            .O(N__19936),
            .I(r_Bit_Index_2));
    InMux I__2358 (
            .O(N__19927),
            .I(N__19922));
    InMux I__2357 (
            .O(N__19926),
            .I(N__19919));
    CascadeMux I__2356 (
            .O(N__19925),
            .I(N__19914));
    LocalMux I__2355 (
            .O(N__19922),
            .I(N__19910));
    LocalMux I__2354 (
            .O(N__19919),
            .I(N__19907));
    InMux I__2353 (
            .O(N__19918),
            .I(N__19904));
    InMux I__2352 (
            .O(N__19917),
            .I(N__19901));
    InMux I__2351 (
            .O(N__19914),
            .I(N__19896));
    InMux I__2350 (
            .O(N__19913),
            .I(N__19896));
    Span12Mux_v I__2349 (
            .O(N__19910),
            .I(N__19893));
    Span4Mux_v I__2348 (
            .O(N__19907),
            .I(N__19890));
    LocalMux I__2347 (
            .O(N__19904),
            .I(N__19885));
    LocalMux I__2346 (
            .O(N__19901),
            .I(N__19885));
    LocalMux I__2345 (
            .O(N__19896),
            .I(N__19882));
    Odrv12 I__2344 (
            .O(N__19893),
            .I(r_Bit_Index_1_adj_2438));
    Odrv4 I__2343 (
            .O(N__19890),
            .I(r_Bit_Index_1_adj_2438));
    Odrv12 I__2342 (
            .O(N__19885),
            .I(r_Bit_Index_1_adj_2438));
    Odrv4 I__2341 (
            .O(N__19882),
            .I(r_Bit_Index_1_adj_2438));
    InMux I__2340 (
            .O(N__19873),
            .I(N__19869));
    CascadeMux I__2339 (
            .O(N__19872),
            .I(N__19866));
    LocalMux I__2338 (
            .O(N__19869),
            .I(N__19860));
    InMux I__2337 (
            .O(N__19866),
            .I(N__19855));
    InMux I__2336 (
            .O(N__19865),
            .I(N__19855));
    InMux I__2335 (
            .O(N__19864),
            .I(N__19852));
    InMux I__2334 (
            .O(N__19863),
            .I(N__19849));
    Span4Mux_h I__2333 (
            .O(N__19860),
            .I(N__19846));
    LocalMux I__2332 (
            .O(N__19855),
            .I(N__19843));
    LocalMux I__2331 (
            .O(N__19852),
            .I(r_Clock_Count_7));
    LocalMux I__2330 (
            .O(N__19849),
            .I(r_Clock_Count_7));
    Odrv4 I__2329 (
            .O(N__19846),
            .I(r_Clock_Count_7));
    Odrv4 I__2328 (
            .O(N__19843),
            .I(r_Clock_Count_7));
    InMux I__2327 (
            .O(N__19834),
            .I(N__19831));
    LocalMux I__2326 (
            .O(N__19831),
            .I(N__19828));
    Span4Mux_s3_h I__2325 (
            .O(N__19828),
            .I(N__19821));
    InMux I__2324 (
            .O(N__19827),
            .I(N__19816));
    InMux I__2323 (
            .O(N__19826),
            .I(N__19816));
    InMux I__2322 (
            .O(N__19825),
            .I(N__19811));
    InMux I__2321 (
            .O(N__19824),
            .I(N__19811));
    Odrv4 I__2320 (
            .O(N__19821),
            .I(r_Clock_Count_6));
    LocalMux I__2319 (
            .O(N__19816),
            .I(r_Clock_Count_6));
    LocalMux I__2318 (
            .O(N__19811),
            .I(r_Clock_Count_6));
    InMux I__2317 (
            .O(N__19804),
            .I(N__19797));
    InMux I__2316 (
            .O(N__19803),
            .I(N__19797));
    InMux I__2315 (
            .O(N__19802),
            .I(N__19794));
    LocalMux I__2314 (
            .O(N__19797),
            .I(N__19787));
    LocalMux I__2313 (
            .O(N__19794),
            .I(N__19787));
    InMux I__2312 (
            .O(N__19793),
            .I(N__19782));
    InMux I__2311 (
            .O(N__19792),
            .I(N__19782));
    Span4Mux_h I__2310 (
            .O(N__19787),
            .I(N__19779));
    LocalMux I__2309 (
            .O(N__19782),
            .I(r_Clock_Count_8));
    Odrv4 I__2308 (
            .O(N__19779),
            .I(r_Clock_Count_8));
    InMux I__2307 (
            .O(N__19774),
            .I(N__19771));
    LocalMux I__2306 (
            .O(N__19771),
            .I(N__19768));
    Span4Mux_s3_h I__2305 (
            .O(N__19768),
            .I(N__19764));
    InMux I__2304 (
            .O(N__19767),
            .I(N__19761));
    Odrv4 I__2303 (
            .O(N__19764),
            .I(n9937));
    LocalMux I__2302 (
            .O(N__19761),
            .I(n9937));
    CascadeMux I__2301 (
            .O(N__19756),
            .I(\c0.tx.n15683_cascade_ ));
    InMux I__2300 (
            .O(N__19753),
            .I(N__19749));
    InMux I__2299 (
            .O(N__19752),
            .I(N__19745));
    LocalMux I__2298 (
            .O(N__19749),
            .I(N__19742));
    InMux I__2297 (
            .O(N__19748),
            .I(N__19739));
    LocalMux I__2296 (
            .O(N__19745),
            .I(\c0.tx.n14082 ));
    Odrv4 I__2295 (
            .O(N__19742),
            .I(\c0.tx.n14082 ));
    LocalMux I__2294 (
            .O(N__19739),
            .I(\c0.tx.n14082 ));
    InMux I__2293 (
            .O(N__19732),
            .I(N__19729));
    LocalMux I__2292 (
            .O(N__19729),
            .I(N__19726));
    Odrv4 I__2291 (
            .O(N__19726),
            .I(n17573));
    InMux I__2290 (
            .O(N__19723),
            .I(N__19718));
    InMux I__2289 (
            .O(N__19722),
            .I(N__19715));
    InMux I__2288 (
            .O(N__19721),
            .I(N__19712));
    LocalMux I__2287 (
            .O(N__19718),
            .I(N__19709));
    LocalMux I__2286 (
            .O(N__19715),
            .I(N__19706));
    LocalMux I__2285 (
            .O(N__19712),
            .I(r_Clock_Count_4));
    Odrv12 I__2284 (
            .O(N__19709),
            .I(r_Clock_Count_4));
    Odrv4 I__2283 (
            .O(N__19706),
            .I(r_Clock_Count_4));
    CascadeMux I__2282 (
            .O(N__19699),
            .I(\c0.n12993_cascade_ ));
    InMux I__2281 (
            .O(N__19696),
            .I(N__19693));
    LocalMux I__2280 (
            .O(N__19693),
            .I(N__19690));
    Span12Mux_v I__2279 (
            .O(N__19690),
            .I(N__19687));
    Odrv12 I__2278 (
            .O(N__19687),
            .I(n16856));
    CascadeMux I__2277 (
            .O(N__19684),
            .I(N__19681));
    InMux I__2276 (
            .O(N__19681),
            .I(N__19673));
    InMux I__2275 (
            .O(N__19680),
            .I(N__19673));
    InMux I__2274 (
            .O(N__19679),
            .I(N__19669));
    InMux I__2273 (
            .O(N__19678),
            .I(N__19666));
    LocalMux I__2272 (
            .O(N__19673),
            .I(N__19663));
    InMux I__2271 (
            .O(N__19672),
            .I(N__19660));
    LocalMux I__2270 (
            .O(N__19669),
            .I(N__19656));
    LocalMux I__2269 (
            .O(N__19666),
            .I(N__19649));
    Span4Mux_s2_h I__2268 (
            .O(N__19663),
            .I(N__19649));
    LocalMux I__2267 (
            .O(N__19660),
            .I(N__19649));
    InMux I__2266 (
            .O(N__19659),
            .I(N__19646));
    Span4Mux_v I__2265 (
            .O(N__19656),
            .I(N__19643));
    Span4Mux_v I__2264 (
            .O(N__19649),
            .I(N__19640));
    LocalMux I__2263 (
            .O(N__19646),
            .I(r_Clock_Count_6_adj_2431));
    Odrv4 I__2262 (
            .O(N__19643),
            .I(r_Clock_Count_6_adj_2431));
    Odrv4 I__2261 (
            .O(N__19640),
            .I(r_Clock_Count_6_adj_2431));
    CascadeMux I__2260 (
            .O(N__19633),
            .I(n16893_cascade_));
    InMux I__2259 (
            .O(N__19630),
            .I(N__19627));
    LocalMux I__2258 (
            .O(N__19627),
            .I(n5));
    InMux I__2257 (
            .O(N__19624),
            .I(N__19621));
    LocalMux I__2256 (
            .O(N__19621),
            .I(N__19618));
    Span4Mux_h I__2255 (
            .O(N__19618),
            .I(N__19615));
    Odrv4 I__2254 (
            .O(N__19615),
            .I(n17636));
    InMux I__2253 (
            .O(N__19612),
            .I(N__19603));
    InMux I__2252 (
            .O(N__19611),
            .I(N__19603));
    InMux I__2251 (
            .O(N__19610),
            .I(N__19603));
    LocalMux I__2250 (
            .O(N__19603),
            .I(data_in_2_4));
    InMux I__2249 (
            .O(N__19600),
            .I(N__19592));
    InMux I__2248 (
            .O(N__19599),
            .I(N__19592));
    InMux I__2247 (
            .O(N__19598),
            .I(N__19587));
    InMux I__2246 (
            .O(N__19597),
            .I(N__19587));
    LocalMux I__2245 (
            .O(N__19592),
            .I(data_in_1_4));
    LocalMux I__2244 (
            .O(N__19587),
            .I(data_in_1_4));
    InMux I__2243 (
            .O(N__19582),
            .I(N__19579));
    LocalMux I__2242 (
            .O(N__19579),
            .I(N__19576));
    Span4Mux_h I__2241 (
            .O(N__19576),
            .I(N__19573));
    Odrv4 I__2240 (
            .O(N__19573),
            .I(n17567));
    InMux I__2239 (
            .O(N__19570),
            .I(N__19566));
    InMux I__2238 (
            .O(N__19569),
            .I(N__19563));
    LocalMux I__2237 (
            .O(N__19566),
            .I(N__19559));
    LocalMux I__2236 (
            .O(N__19563),
            .I(N__19556));
    InMux I__2235 (
            .O(N__19562),
            .I(N__19553));
    Span4Mux_s3_h I__2234 (
            .O(N__19559),
            .I(N__19548));
    Span4Mux_s3_h I__2233 (
            .O(N__19556),
            .I(N__19548));
    LocalMux I__2232 (
            .O(N__19553),
            .I(r_Clock_Count_4_adj_2450));
    Odrv4 I__2231 (
            .O(N__19548),
            .I(r_Clock_Count_4_adj_2450));
    InMux I__2230 (
            .O(N__19543),
            .I(N__19537));
    InMux I__2229 (
            .O(N__19542),
            .I(N__19532));
    InMux I__2228 (
            .O(N__19541),
            .I(N__19532));
    InMux I__2227 (
            .O(N__19540),
            .I(N__19529));
    LocalMux I__2226 (
            .O(N__19537),
            .I(data_in_2_3));
    LocalMux I__2225 (
            .O(N__19532),
            .I(data_in_2_3));
    LocalMux I__2224 (
            .O(N__19529),
            .I(data_in_2_3));
    InMux I__2223 (
            .O(N__19522),
            .I(N__19519));
    LocalMux I__2222 (
            .O(N__19519),
            .I(N__19516));
    Odrv12 I__2221 (
            .O(N__19516),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_29 ));
    InMux I__2220 (
            .O(N__19513),
            .I(\c0.n15650 ));
    InMux I__2219 (
            .O(N__19510),
            .I(N__19507));
    LocalMux I__2218 (
            .O(N__19507),
            .I(N__19504));
    Sp12to4 I__2217 (
            .O(N__19504),
            .I(N__19501));
    Odrv12 I__2216 (
            .O(N__19501),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_30 ));
    InMux I__2215 (
            .O(N__19498),
            .I(\c0.n15651 ));
    InMux I__2214 (
            .O(N__19495),
            .I(\c0.n15652 ));
    InMux I__2213 (
            .O(N__19492),
            .I(N__19489));
    LocalMux I__2212 (
            .O(N__19489),
            .I(N__19486));
    Span4Mux_s2_h I__2211 (
            .O(N__19486),
            .I(N__19483));
    Span4Mux_v I__2210 (
            .O(N__19483),
            .I(N__19480));
    Odrv4 I__2209 (
            .O(N__19480),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_31 ));
    InMux I__2208 (
            .O(N__19477),
            .I(N__19472));
    InMux I__2207 (
            .O(N__19476),
            .I(N__19469));
    InMux I__2206 (
            .O(N__19475),
            .I(N__19466));
    LocalMux I__2205 (
            .O(N__19472),
            .I(data_in_0_6));
    LocalMux I__2204 (
            .O(N__19469),
            .I(data_in_0_6));
    LocalMux I__2203 (
            .O(N__19466),
            .I(data_in_0_6));
    CascadeMux I__2202 (
            .O(N__19459),
            .I(\c0.n17274_cascade_ ));
    CascadeMux I__2201 (
            .O(N__19456),
            .I(N__19433));
    CascadeMux I__2200 (
            .O(N__19455),
            .I(N__19430));
    CascadeMux I__2199 (
            .O(N__19454),
            .I(N__19427));
    CascadeMux I__2198 (
            .O(N__19453),
            .I(N__19424));
    CascadeMux I__2197 (
            .O(N__19452),
            .I(N__19421));
    CascadeMux I__2196 (
            .O(N__19451),
            .I(N__19417));
    CascadeMux I__2195 (
            .O(N__19450),
            .I(N__19414));
    CascadeMux I__2194 (
            .O(N__19449),
            .I(N__19410));
    CascadeMux I__2193 (
            .O(N__19448),
            .I(N__19407));
    CascadeMux I__2192 (
            .O(N__19447),
            .I(N__19404));
    CascadeMux I__2191 (
            .O(N__19446),
            .I(N__19399));
    CascadeMux I__2190 (
            .O(N__19445),
            .I(N__19395));
    CascadeMux I__2189 (
            .O(N__19444),
            .I(N__19391));
    CascadeMux I__2188 (
            .O(N__19443),
            .I(N__19387));
    CascadeMux I__2187 (
            .O(N__19442),
            .I(N__19384));
    CascadeMux I__2186 (
            .O(N__19441),
            .I(N__19380));
    CascadeMux I__2185 (
            .O(N__19440),
            .I(N__19376));
    CascadeMux I__2184 (
            .O(N__19439),
            .I(N__19372));
    CascadeMux I__2183 (
            .O(N__19438),
            .I(N__19368));
    CascadeMux I__2182 (
            .O(N__19437),
            .I(N__19365));
    CascadeMux I__2181 (
            .O(N__19436),
            .I(N__19362));
    InMux I__2180 (
            .O(N__19433),
            .I(N__19355));
    InMux I__2179 (
            .O(N__19430),
            .I(N__19355));
    InMux I__2178 (
            .O(N__19427),
            .I(N__19355));
    InMux I__2177 (
            .O(N__19424),
            .I(N__19344));
    InMux I__2176 (
            .O(N__19421),
            .I(N__19344));
    InMux I__2175 (
            .O(N__19420),
            .I(N__19344));
    InMux I__2174 (
            .O(N__19417),
            .I(N__19344));
    InMux I__2173 (
            .O(N__19414),
            .I(N__19344));
    InMux I__2172 (
            .O(N__19413),
            .I(N__19333));
    InMux I__2171 (
            .O(N__19410),
            .I(N__19333));
    InMux I__2170 (
            .O(N__19407),
            .I(N__19333));
    InMux I__2169 (
            .O(N__19404),
            .I(N__19333));
    InMux I__2168 (
            .O(N__19403),
            .I(N__19333));
    InMux I__2167 (
            .O(N__19402),
            .I(N__19316));
    InMux I__2166 (
            .O(N__19399),
            .I(N__19316));
    InMux I__2165 (
            .O(N__19398),
            .I(N__19316));
    InMux I__2164 (
            .O(N__19395),
            .I(N__19316));
    InMux I__2163 (
            .O(N__19394),
            .I(N__19316));
    InMux I__2162 (
            .O(N__19391),
            .I(N__19316));
    InMux I__2161 (
            .O(N__19390),
            .I(N__19316));
    InMux I__2160 (
            .O(N__19387),
            .I(N__19316));
    InMux I__2159 (
            .O(N__19384),
            .I(N__19299));
    InMux I__2158 (
            .O(N__19383),
            .I(N__19299));
    InMux I__2157 (
            .O(N__19380),
            .I(N__19299));
    InMux I__2156 (
            .O(N__19379),
            .I(N__19299));
    InMux I__2155 (
            .O(N__19376),
            .I(N__19299));
    InMux I__2154 (
            .O(N__19375),
            .I(N__19299));
    InMux I__2153 (
            .O(N__19372),
            .I(N__19299));
    InMux I__2152 (
            .O(N__19371),
            .I(N__19299));
    InMux I__2151 (
            .O(N__19368),
            .I(N__19292));
    InMux I__2150 (
            .O(N__19365),
            .I(N__19292));
    InMux I__2149 (
            .O(N__19362),
            .I(N__19292));
    LocalMux I__2148 (
            .O(N__19355),
            .I(N__19287));
    LocalMux I__2147 (
            .O(N__19344),
            .I(N__19287));
    LocalMux I__2146 (
            .O(N__19333),
            .I(N__19280));
    LocalMux I__2145 (
            .O(N__19316),
            .I(N__19280));
    LocalMux I__2144 (
            .O(N__19299),
            .I(N__19280));
    LocalMux I__2143 (
            .O(N__19292),
            .I(\c0.n17889 ));
    Odrv4 I__2142 (
            .O(N__19287),
            .I(\c0.n17889 ));
    Odrv12 I__2141 (
            .O(N__19280),
            .I(\c0.n17889 ));
    InMux I__2140 (
            .O(N__19273),
            .I(N__19268));
    InMux I__2139 (
            .O(N__19272),
            .I(N__19265));
    InMux I__2138 (
            .O(N__19271),
            .I(N__19262));
    LocalMux I__2137 (
            .O(N__19268),
            .I(N__19259));
    LocalMux I__2136 (
            .O(N__19265),
            .I(data_in_3_1));
    LocalMux I__2135 (
            .O(N__19262),
            .I(data_in_3_1));
    Odrv4 I__2134 (
            .O(N__19259),
            .I(data_in_3_1));
    InMux I__2133 (
            .O(N__19252),
            .I(N__19247));
    CascadeMux I__2132 (
            .O(N__19251),
            .I(N__19244));
    CascadeMux I__2131 (
            .O(N__19250),
            .I(N__19241));
    LocalMux I__2130 (
            .O(N__19247),
            .I(N__19238));
    InMux I__2129 (
            .O(N__19244),
            .I(N__19233));
    InMux I__2128 (
            .O(N__19241),
            .I(N__19233));
    Odrv4 I__2127 (
            .O(N__19238),
            .I(data_in_2_1));
    LocalMux I__2126 (
            .O(N__19233),
            .I(data_in_2_1));
    InMux I__2125 (
            .O(N__19228),
            .I(N__19225));
    LocalMux I__2124 (
            .O(N__19225),
            .I(N__19222));
    Span4Mux_v I__2123 (
            .O(N__19222),
            .I(N__19219));
    Odrv4 I__2122 (
            .O(N__19219),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_20 ));
    InMux I__2121 (
            .O(N__19216),
            .I(\c0.n15641 ));
    InMux I__2120 (
            .O(N__19213),
            .I(N__19210));
    LocalMux I__2119 (
            .O(N__19210),
            .I(N__19207));
    Span4Mux_h I__2118 (
            .O(N__19207),
            .I(N__19204));
    Span4Mux_v I__2117 (
            .O(N__19204),
            .I(N__19201));
    Odrv4 I__2116 (
            .O(N__19201),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_21 ));
    InMux I__2115 (
            .O(N__19198),
            .I(\c0.n15642 ));
    InMux I__2114 (
            .O(N__19195),
            .I(N__19192));
    LocalMux I__2113 (
            .O(N__19192),
            .I(N__19189));
    Span4Mux_s3_h I__2112 (
            .O(N__19189),
            .I(N__19186));
    Odrv4 I__2111 (
            .O(N__19186),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_22 ));
    InMux I__2110 (
            .O(N__19183),
            .I(\c0.n15643 ));
    InMux I__2109 (
            .O(N__19180),
            .I(N__19177));
    LocalMux I__2108 (
            .O(N__19177),
            .I(N__19174));
    Span4Mux_s1_h I__2107 (
            .O(N__19174),
            .I(N__19171));
    Span4Mux_v I__2106 (
            .O(N__19171),
            .I(N__19168));
    Odrv4 I__2105 (
            .O(N__19168),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_23 ));
    InMux I__2104 (
            .O(N__19165),
            .I(\c0.n15644 ));
    InMux I__2103 (
            .O(N__19162),
            .I(N__19159));
    LocalMux I__2102 (
            .O(N__19159),
            .I(N__19156));
    Odrv12 I__2101 (
            .O(N__19156),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_24 ));
    InMux I__2100 (
            .O(N__19153),
            .I(bfn_4_25_0_));
    InMux I__2099 (
            .O(N__19150),
            .I(N__19147));
    LocalMux I__2098 (
            .O(N__19147),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_25 ));
    InMux I__2097 (
            .O(N__19144),
            .I(\c0.n15646 ));
    InMux I__2096 (
            .O(N__19141),
            .I(N__19138));
    LocalMux I__2095 (
            .O(N__19138),
            .I(N__19135));
    Span4Mux_s3_h I__2094 (
            .O(N__19135),
            .I(N__19132));
    Odrv4 I__2093 (
            .O(N__19132),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_26 ));
    InMux I__2092 (
            .O(N__19129),
            .I(\c0.n15647 ));
    InMux I__2091 (
            .O(N__19126),
            .I(N__19123));
    LocalMux I__2090 (
            .O(N__19123),
            .I(N__19120));
    Span4Mux_s3_h I__2089 (
            .O(N__19120),
            .I(N__19117));
    Odrv4 I__2088 (
            .O(N__19117),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_27 ));
    InMux I__2087 (
            .O(N__19114),
            .I(\c0.n15648 ));
    InMux I__2086 (
            .O(N__19111),
            .I(N__19108));
    LocalMux I__2085 (
            .O(N__19108),
            .I(N__19105));
    Sp12to4 I__2084 (
            .O(N__19105),
            .I(N__19102));
    Odrv12 I__2083 (
            .O(N__19102),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_28 ));
    InMux I__2082 (
            .O(N__19099),
            .I(\c0.n15649 ));
    InMux I__2081 (
            .O(N__19096),
            .I(N__19093));
    LocalMux I__2080 (
            .O(N__19093),
            .I(N__19090));
    Odrv4 I__2079 (
            .O(N__19090),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_12 ));
    InMux I__2078 (
            .O(N__19087),
            .I(\c0.n15633 ));
    InMux I__2077 (
            .O(N__19084),
            .I(N__19081));
    LocalMux I__2076 (
            .O(N__19081),
            .I(N__19078));
    Odrv4 I__2075 (
            .O(N__19078),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_13 ));
    InMux I__2074 (
            .O(N__19075),
            .I(N__19072));
    LocalMux I__2073 (
            .O(N__19072),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_13 ));
    InMux I__2072 (
            .O(N__19069),
            .I(\c0.n15634 ));
    InMux I__2071 (
            .O(N__19066),
            .I(N__19063));
    LocalMux I__2070 (
            .O(N__19063),
            .I(N__19060));
    Odrv12 I__2069 (
            .O(N__19060),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_14 ));
    InMux I__2068 (
            .O(N__19057),
            .I(N__19054));
    LocalMux I__2067 (
            .O(N__19054),
            .I(N__19051));
    Odrv4 I__2066 (
            .O(N__19051),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_14 ));
    InMux I__2065 (
            .O(N__19048),
            .I(\c0.n15635 ));
    InMux I__2064 (
            .O(N__19045),
            .I(N__19042));
    LocalMux I__2063 (
            .O(N__19042),
            .I(N__19039));
    Odrv4 I__2062 (
            .O(N__19039),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_15 ));
    InMux I__2061 (
            .O(N__19036),
            .I(N__19033));
    LocalMux I__2060 (
            .O(N__19033),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_15 ));
    InMux I__2059 (
            .O(N__19030),
            .I(\c0.n15636 ));
    InMux I__2058 (
            .O(N__19027),
            .I(bfn_4_24_0_));
    InMux I__2057 (
            .O(N__19024),
            .I(\c0.n15638 ));
    InMux I__2056 (
            .O(N__19021),
            .I(\c0.n15639 ));
    InMux I__2055 (
            .O(N__19018),
            .I(N__19015));
    LocalMux I__2054 (
            .O(N__19015),
            .I(N__19012));
    Odrv4 I__2053 (
            .O(N__19012),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_19 ));
    InMux I__2052 (
            .O(N__19009),
            .I(\c0.n15640 ));
    InMux I__2051 (
            .O(N__19006),
            .I(\c0.n15624 ));
    InMux I__2050 (
            .O(N__19003),
            .I(N__19000));
    LocalMux I__2049 (
            .O(N__19000),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_4 ));
    InMux I__2048 (
            .O(N__18997),
            .I(\c0.n15625 ));
    InMux I__2047 (
            .O(N__18994),
            .I(N__18991));
    LocalMux I__2046 (
            .O(N__18991),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_5 ));
    InMux I__2045 (
            .O(N__18988),
            .I(N__18985));
    LocalMux I__2044 (
            .O(N__18985),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_5 ));
    InMux I__2043 (
            .O(N__18982),
            .I(\c0.n15626 ));
    InMux I__2042 (
            .O(N__18979),
            .I(N__18976));
    LocalMux I__2041 (
            .O(N__18976),
            .I(N__18973));
    Odrv4 I__2040 (
            .O(N__18973),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_6 ));
    InMux I__2039 (
            .O(N__18970),
            .I(\c0.n15627 ));
    InMux I__2038 (
            .O(N__18967),
            .I(\c0.n15628 ));
    InMux I__2037 (
            .O(N__18964),
            .I(N__18961));
    LocalMux I__2036 (
            .O(N__18961),
            .I(N__18958));
    Odrv12 I__2035 (
            .O(N__18958),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_8 ));
    InMux I__2034 (
            .O(N__18955),
            .I(bfn_4_23_0_));
    InMux I__2033 (
            .O(N__18952),
            .I(N__18949));
    LocalMux I__2032 (
            .O(N__18949),
            .I(N__18946));
    Span4Mux_s3_h I__2031 (
            .O(N__18946),
            .I(N__18943));
    Odrv4 I__2030 (
            .O(N__18943),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_9 ));
    InMux I__2029 (
            .O(N__18940),
            .I(\c0.n15630 ));
    InMux I__2028 (
            .O(N__18937),
            .I(\c0.n15631 ));
    InMux I__2027 (
            .O(N__18934),
            .I(\c0.n15632 ));
    SRMux I__2026 (
            .O(N__18931),
            .I(N__18928));
    LocalMux I__2025 (
            .O(N__18928),
            .I(N__18925));
    Span4Mux_h I__2024 (
            .O(N__18925),
            .I(N__18922));
    Odrv4 I__2023 (
            .O(N__18922),
            .I(\c0.n3_adj_2259 ));
    InMux I__2022 (
            .O(N__18919),
            .I(N__18916));
    LocalMux I__2021 (
            .O(N__18916),
            .I(\c0.n10_adj_2329 ));
    InMux I__2020 (
            .O(N__18913),
            .I(N__18910));
    LocalMux I__2019 (
            .O(N__18910),
            .I(\c0.n16895 ));
    CascadeMux I__2018 (
            .O(N__18907),
            .I(\c0.n16895_cascade_ ));
    CascadeMux I__2017 (
            .O(N__18904),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_1_cascade_ ));
    SRMux I__2016 (
            .O(N__18901),
            .I(N__18898));
    LocalMux I__2015 (
            .O(N__18898),
            .I(N__18895));
    Span4Mux_v I__2014 (
            .O(N__18895),
            .I(N__18892));
    Odrv4 I__2013 (
            .O(N__18892),
            .I(\c0.n3_adj_2260 ));
    InMux I__2012 (
            .O(N__18889),
            .I(bfn_4_22_0_));
    InMux I__2011 (
            .O(N__18886),
            .I(N__18883));
    LocalMux I__2010 (
            .O(N__18883),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_1 ));
    CascadeMux I__2009 (
            .O(N__18880),
            .I(N__18877));
    InMux I__2008 (
            .O(N__18877),
            .I(N__18874));
    LocalMux I__2007 (
            .O(N__18874),
            .I(N__18871));
    Span4Mux_v I__2006 (
            .O(N__18871),
            .I(N__18868));
    Odrv4 I__2005 (
            .O(N__18868),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_1 ));
    InMux I__2004 (
            .O(N__18865),
            .I(\c0.n15622 ));
    InMux I__2003 (
            .O(N__18862),
            .I(N__18859));
    LocalMux I__2002 (
            .O(N__18859),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_2 ));
    InMux I__2001 (
            .O(N__18856),
            .I(N__18853));
    LocalMux I__2000 (
            .O(N__18853),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_2 ));
    InMux I__1999 (
            .O(N__18850),
            .I(\c0.n15623 ));
    InMux I__1998 (
            .O(N__18847),
            .I(N__18844));
    LocalMux I__1997 (
            .O(N__18844),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_3 ));
    InMux I__1996 (
            .O(N__18841),
            .I(N__18838));
    LocalMux I__1995 (
            .O(N__18838),
            .I(N__18835));
    Odrv4 I__1994 (
            .O(N__18835),
            .I(\c0.FRAME_MATCHER_i_31_N_1280_3 ));
    SRMux I__1993 (
            .O(N__18832),
            .I(N__18829));
    LocalMux I__1992 (
            .O(N__18829),
            .I(N__18826));
    Odrv4 I__1991 (
            .O(N__18826),
            .I(\c0.n3_adj_2217 ));
    SRMux I__1990 (
            .O(N__18823),
            .I(N__18820));
    LocalMux I__1989 (
            .O(N__18820),
            .I(\c0.n3_adj_2215 ));
    SRMux I__1988 (
            .O(N__18817),
            .I(N__18814));
    LocalMux I__1987 (
            .O(N__18814),
            .I(N__18811));
    Span4Mux_s3_h I__1986 (
            .O(N__18811),
            .I(N__18808));
    Span4Mux_h I__1985 (
            .O(N__18808),
            .I(N__18805));
    Odrv4 I__1984 (
            .O(N__18805),
            .I(\c0.n3_adj_2210 ));
    SRMux I__1983 (
            .O(N__18802),
            .I(N__18799));
    LocalMux I__1982 (
            .O(N__18799),
            .I(N__18796));
    Span4Mux_v I__1981 (
            .O(N__18796),
            .I(N__18793));
    Span4Mux_s0_h I__1980 (
            .O(N__18793),
            .I(N__18790));
    Odrv4 I__1979 (
            .O(N__18790),
            .I(\c0.n3_adj_2249 ));
    InMux I__1978 (
            .O(N__18787),
            .I(N__18784));
    LocalMux I__1977 (
            .O(N__18784),
            .I(\c0.n9393 ));
    CascadeMux I__1976 (
            .O(N__18781),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_2_cascade_ ));
    InMux I__1975 (
            .O(N__18778),
            .I(N__18775));
    LocalMux I__1974 (
            .O(N__18775),
            .I(n16857));
    CascadeMux I__1973 (
            .O(N__18772),
            .I(N__18766));
    InMux I__1972 (
            .O(N__18771),
            .I(N__18763));
    InMux I__1971 (
            .O(N__18770),
            .I(N__18758));
    InMux I__1970 (
            .O(N__18769),
            .I(N__18758));
    InMux I__1969 (
            .O(N__18766),
            .I(N__18753));
    LocalMux I__1968 (
            .O(N__18763),
            .I(N__18748));
    LocalMux I__1967 (
            .O(N__18758),
            .I(N__18748));
    InMux I__1966 (
            .O(N__18757),
            .I(N__18744));
    InMux I__1965 (
            .O(N__18756),
            .I(N__18741));
    LocalMux I__1964 (
            .O(N__18753),
            .I(N__18736));
    Span4Mux_s1_v I__1963 (
            .O(N__18748),
            .I(N__18736));
    InMux I__1962 (
            .O(N__18747),
            .I(N__18733));
    LocalMux I__1961 (
            .O(N__18744),
            .I(r_Clock_Count_5_adj_2432));
    LocalMux I__1960 (
            .O(N__18741),
            .I(r_Clock_Count_5_adj_2432));
    Odrv4 I__1959 (
            .O(N__18736),
            .I(r_Clock_Count_5_adj_2432));
    LocalMux I__1958 (
            .O(N__18733),
            .I(r_Clock_Count_5_adj_2432));
    InMux I__1957 (
            .O(N__18724),
            .I(N__18721));
    LocalMux I__1956 (
            .O(N__18721),
            .I(n16858));
    InMux I__1955 (
            .O(N__18718),
            .I(N__18714));
    CascadeMux I__1954 (
            .O(N__18717),
            .I(N__18710));
    LocalMux I__1953 (
            .O(N__18714),
            .I(N__18707));
    InMux I__1952 (
            .O(N__18713),
            .I(N__18704));
    InMux I__1951 (
            .O(N__18710),
            .I(N__18701));
    Odrv4 I__1950 (
            .O(N__18707),
            .I(r_Clock_Count_3_adj_2434));
    LocalMux I__1949 (
            .O(N__18704),
            .I(r_Clock_Count_3_adj_2434));
    LocalMux I__1948 (
            .O(N__18701),
            .I(r_Clock_Count_3_adj_2434));
    InMux I__1947 (
            .O(N__18694),
            .I(N__18691));
    LocalMux I__1946 (
            .O(N__18691),
            .I(N__18688));
    Odrv4 I__1945 (
            .O(N__18688),
            .I(n9406));
    InMux I__1944 (
            .O(N__18685),
            .I(N__18682));
    LocalMux I__1943 (
            .O(N__18682),
            .I(N__18679));
    Odrv4 I__1942 (
            .O(N__18679),
            .I(n17461));
    InMux I__1941 (
            .O(N__18676),
            .I(N__18672));
    InMux I__1940 (
            .O(N__18675),
            .I(N__18668));
    LocalMux I__1939 (
            .O(N__18672),
            .I(N__18665));
    InMux I__1938 (
            .O(N__18671),
            .I(N__18662));
    LocalMux I__1937 (
            .O(N__18668),
            .I(r_Clock_Count_1));
    Odrv4 I__1936 (
            .O(N__18665),
            .I(r_Clock_Count_1));
    LocalMux I__1935 (
            .O(N__18662),
            .I(r_Clock_Count_1));
    InMux I__1934 (
            .O(N__18655),
            .I(N__18652));
    LocalMux I__1933 (
            .O(N__18652),
            .I(N__18649));
    Span4Mux_h I__1932 (
            .O(N__18649),
            .I(N__18646));
    Odrv4 I__1931 (
            .O(N__18646),
            .I(n17601));
    InMux I__1930 (
            .O(N__18643),
            .I(N__18640));
    LocalMux I__1929 (
            .O(N__18640),
            .I(N__18637));
    Span4Mux_h I__1928 (
            .O(N__18637),
            .I(N__18634));
    Odrv4 I__1927 (
            .O(N__18634),
            .I(n17602));
    InMux I__1926 (
            .O(N__18631),
            .I(N__18627));
    InMux I__1925 (
            .O(N__18630),
            .I(N__18623));
    LocalMux I__1924 (
            .O(N__18627),
            .I(N__18620));
    InMux I__1923 (
            .O(N__18626),
            .I(N__18617));
    LocalMux I__1922 (
            .O(N__18623),
            .I(r_Clock_Count_4_adj_2433));
    Odrv4 I__1921 (
            .O(N__18620),
            .I(r_Clock_Count_4_adj_2433));
    LocalMux I__1920 (
            .O(N__18617),
            .I(r_Clock_Count_4_adj_2433));
    InMux I__1919 (
            .O(N__18610),
            .I(N__18607));
    LocalMux I__1918 (
            .O(N__18607),
            .I(\c0.rx.n6 ));
    InMux I__1917 (
            .O(N__18604),
            .I(N__18601));
    LocalMux I__1916 (
            .O(N__18601),
            .I(N__18598));
    Odrv4 I__1915 (
            .O(N__18598),
            .I(n16853));
    CascadeMux I__1914 (
            .O(N__18595),
            .I(N__18592));
    InMux I__1913 (
            .O(N__18592),
            .I(N__18589));
    LocalMux I__1912 (
            .O(N__18589),
            .I(N__18584));
    InMux I__1911 (
            .O(N__18588),
            .I(N__18579));
    InMux I__1910 (
            .O(N__18587),
            .I(N__18579));
    Odrv4 I__1909 (
            .O(N__18584),
            .I(r_Clock_Count_1_adj_2436));
    LocalMux I__1908 (
            .O(N__18579),
            .I(r_Clock_Count_1_adj_2436));
    InMux I__1907 (
            .O(N__18574),
            .I(N__18569));
    InMux I__1906 (
            .O(N__18573),
            .I(N__18564));
    InMux I__1905 (
            .O(N__18572),
            .I(N__18564));
    LocalMux I__1904 (
            .O(N__18569),
            .I(N__18561));
    LocalMux I__1903 (
            .O(N__18564),
            .I(N__18558));
    Odrv12 I__1902 (
            .O(N__18561),
            .I(n4_adj_2411));
    Odrv4 I__1901 (
            .O(N__18558),
            .I(n4_adj_2411));
    InMux I__1900 (
            .O(N__18553),
            .I(N__18547));
    InMux I__1899 (
            .O(N__18552),
            .I(N__18544));
    InMux I__1898 (
            .O(N__18551),
            .I(N__18539));
    InMux I__1897 (
            .O(N__18550),
            .I(N__18539));
    LocalMux I__1896 (
            .O(N__18547),
            .I(N__18534));
    LocalMux I__1895 (
            .O(N__18544),
            .I(N__18534));
    LocalMux I__1894 (
            .O(N__18539),
            .I(N__18531));
    Span4Mux_v I__1893 (
            .O(N__18534),
            .I(N__18528));
    Span4Mux_h I__1892 (
            .O(N__18531),
            .I(N__18525));
    Odrv4 I__1891 (
            .O(N__18528),
            .I(n17260));
    Odrv4 I__1890 (
            .O(N__18525),
            .I(n17260));
    InMux I__1889 (
            .O(N__18520),
            .I(N__18516));
    InMux I__1888 (
            .O(N__18519),
            .I(N__18513));
    LocalMux I__1887 (
            .O(N__18516),
            .I(N__18508));
    LocalMux I__1886 (
            .O(N__18513),
            .I(N__18508));
    Odrv4 I__1885 (
            .O(N__18508),
            .I(n10425));
    CascadeMux I__1884 (
            .O(N__18505),
            .I(n7866_cascade_));
    CascadeMux I__1883 (
            .O(N__18502),
            .I(n10425_cascade_));
    InMux I__1882 (
            .O(N__18499),
            .I(N__18494));
    InMux I__1881 (
            .O(N__18498),
            .I(N__18489));
    InMux I__1880 (
            .O(N__18497),
            .I(N__18489));
    LocalMux I__1879 (
            .O(N__18494),
            .I(N__18486));
    LocalMux I__1878 (
            .O(N__18489),
            .I(n12));
    Odrv4 I__1877 (
            .O(N__18486),
            .I(n12));
    InMux I__1876 (
            .O(N__18481),
            .I(N__18478));
    LocalMux I__1875 (
            .O(N__18478),
            .I(n13276));
    CascadeMux I__1874 (
            .O(N__18475),
            .I(n10_adj_2415_cascade_));
    InMux I__1873 (
            .O(N__18472),
            .I(N__18467));
    InMux I__1872 (
            .O(N__18471),
            .I(N__18464));
    InMux I__1871 (
            .O(N__18470),
            .I(N__18461));
    LocalMux I__1870 (
            .O(N__18467),
            .I(n15701));
    LocalMux I__1869 (
            .O(N__18464),
            .I(n15701));
    LocalMux I__1868 (
            .O(N__18461),
            .I(n15701));
    InMux I__1867 (
            .O(N__18454),
            .I(N__18451));
    LocalMux I__1866 (
            .O(N__18451),
            .I(N__18446));
    InMux I__1865 (
            .O(N__18450),
            .I(N__18443));
    InMux I__1864 (
            .O(N__18449),
            .I(N__18440));
    Span4Mux_s3_h I__1863 (
            .O(N__18446),
            .I(N__18437));
    LocalMux I__1862 (
            .O(N__18443),
            .I(N__18432));
    LocalMux I__1861 (
            .O(N__18440),
            .I(N__18432));
    Odrv4 I__1860 (
            .O(N__18437),
            .I(n16844));
    Odrv4 I__1859 (
            .O(N__18432),
            .I(n16844));
    CascadeMux I__1858 (
            .O(N__18427),
            .I(n9472_cascade_));
    CascadeMux I__1857 (
            .O(N__18424),
            .I(\c0.rx.n10086_cascade_ ));
    InMux I__1856 (
            .O(N__18421),
            .I(N__18417));
    InMux I__1855 (
            .O(N__18420),
            .I(N__18414));
    LocalMux I__1854 (
            .O(N__18417),
            .I(N__18409));
    LocalMux I__1853 (
            .O(N__18414),
            .I(N__18406));
    InMux I__1852 (
            .O(N__18413),
            .I(N__18403));
    InMux I__1851 (
            .O(N__18412),
            .I(N__18400));
    Span4Mux_v I__1850 (
            .O(N__18409),
            .I(N__18397));
    Span4Mux_h I__1849 (
            .O(N__18406),
            .I(N__18392));
    LocalMux I__1848 (
            .O(N__18403),
            .I(N__18392));
    LocalMux I__1847 (
            .O(N__18400),
            .I(N__18389));
    Odrv4 I__1846 (
            .O(N__18397),
            .I(\c0.rx.r_SM_Main_2_N_2090_2 ));
    Odrv4 I__1845 (
            .O(N__18392),
            .I(\c0.rx.r_SM_Main_2_N_2090_2 ));
    Odrv12 I__1844 (
            .O(N__18389),
            .I(\c0.rx.r_SM_Main_2_N_2090_2 ));
    CascadeMux I__1843 (
            .O(N__18382),
            .I(n14060_cascade_));
    InMux I__1842 (
            .O(N__18379),
            .I(N__18375));
    InMux I__1841 (
            .O(N__18378),
            .I(N__18372));
    LocalMux I__1840 (
            .O(N__18375),
            .I(data_in_0_7));
    LocalMux I__1839 (
            .O(N__18372),
            .I(data_in_0_7));
    InMux I__1838 (
            .O(N__18367),
            .I(N__18362));
    InMux I__1837 (
            .O(N__18366),
            .I(N__18359));
    InMux I__1836 (
            .O(N__18365),
            .I(N__18356));
    LocalMux I__1835 (
            .O(N__18362),
            .I(data_in_1_5));
    LocalMux I__1834 (
            .O(N__18359),
            .I(data_in_1_5));
    LocalMux I__1833 (
            .O(N__18356),
            .I(data_in_1_5));
    InMux I__1832 (
            .O(N__18349),
            .I(N__18343));
    InMux I__1831 (
            .O(N__18348),
            .I(N__18343));
    LocalMux I__1830 (
            .O(N__18343),
            .I(data_in_0_4));
    CascadeMux I__1829 (
            .O(N__18340),
            .I(\c0.n17172_cascade_ ));
    SRMux I__1828 (
            .O(N__18337),
            .I(N__18334));
    LocalMux I__1827 (
            .O(N__18334),
            .I(N__18331));
    Odrv4 I__1826 (
            .O(N__18331),
            .I(\c0.n3_adj_2242 ));
    SRMux I__1825 (
            .O(N__18328),
            .I(N__18325));
    LocalMux I__1824 (
            .O(N__18325),
            .I(\c0.n3_adj_2243 ));
    SRMux I__1823 (
            .O(N__18322),
            .I(N__18319));
    LocalMux I__1822 (
            .O(N__18319),
            .I(N__18316));
    Span4Mux_s3_h I__1821 (
            .O(N__18316),
            .I(N__18313));
    Odrv4 I__1820 (
            .O(N__18313),
            .I(\c0.n3_adj_2244 ));
    SRMux I__1819 (
            .O(N__18310),
            .I(N__18307));
    LocalMux I__1818 (
            .O(N__18307),
            .I(N__18304));
    Span4Mux_s3_h I__1817 (
            .O(N__18304),
            .I(N__18301));
    Odrv4 I__1816 (
            .O(N__18301),
            .I(\c0.n3_adj_2256 ));
    CascadeMux I__1815 (
            .O(N__18298),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_4_cascade_ ));
    CascadeMux I__1814 (
            .O(N__18295),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_3_cascade_ ));
    SRMux I__1813 (
            .O(N__18292),
            .I(N__18289));
    LocalMux I__1812 (
            .O(N__18289),
            .I(N__18286));
    Span4Mux_s2_h I__1811 (
            .O(N__18286),
            .I(N__18283));
    Odrv4 I__1810 (
            .O(N__18283),
            .I(\c0.n3_adj_2258 ));
    SRMux I__1809 (
            .O(N__18280),
            .I(N__18277));
    LocalMux I__1808 (
            .O(N__18277),
            .I(N__18274));
    Span4Mux_s3_h I__1807 (
            .O(N__18274),
            .I(N__18271));
    Odrv4 I__1806 (
            .O(N__18271),
            .I(\c0.n16379 ));
    InMux I__1805 (
            .O(N__18268),
            .I(N__18265));
    LocalMux I__1804 (
            .O(N__18265),
            .I(n1651));
    CascadeMux I__1803 (
            .O(N__18262),
            .I(n6_cascade_));
    InMux I__1802 (
            .O(N__18259),
            .I(N__18256));
    LocalMux I__1801 (
            .O(N__18256),
            .I(n4));
    CascadeMux I__1800 (
            .O(N__18253),
            .I(n8_adj_2459_cascade_));
    InMux I__1799 (
            .O(N__18250),
            .I(N__18247));
    LocalMux I__1798 (
            .O(N__18247),
            .I(FRAME_MATCHER_state_31_N_1440_1));
    InMux I__1797 (
            .O(N__18244),
            .I(N__18241));
    LocalMux I__1796 (
            .O(N__18241),
            .I(n3_adj_2408));
    CascadeMux I__1795 (
            .O(N__18238),
            .I(\c0.FRAME_MATCHER_i_31_N_1312_5_cascade_ ));
    InMux I__1794 (
            .O(N__18235),
            .I(N__18232));
    LocalMux I__1793 (
            .O(N__18232),
            .I(N__18229));
    Odrv4 I__1792 (
            .O(N__18229),
            .I(n16854));
    InMux I__1791 (
            .O(N__18226),
            .I(\c0.rx.n15671 ));
    InMux I__1790 (
            .O(N__18223),
            .I(\c0.rx.n15672 ));
    InMux I__1789 (
            .O(N__18220),
            .I(\c0.rx.n15673 ));
    InMux I__1788 (
            .O(N__18217),
            .I(N__18214));
    LocalMux I__1787 (
            .O(N__18214),
            .I(N__18206));
    InMux I__1786 (
            .O(N__18213),
            .I(N__18203));
    InMux I__1785 (
            .O(N__18212),
            .I(N__18200));
    InMux I__1784 (
            .O(N__18211),
            .I(N__18197));
    InMux I__1783 (
            .O(N__18210),
            .I(N__18192));
    InMux I__1782 (
            .O(N__18209),
            .I(N__18192));
    Odrv4 I__1781 (
            .O(N__18206),
            .I(r_Clock_Count_7_adj_2430));
    LocalMux I__1780 (
            .O(N__18203),
            .I(r_Clock_Count_7_adj_2430));
    LocalMux I__1779 (
            .O(N__18200),
            .I(r_Clock_Count_7_adj_2430));
    LocalMux I__1778 (
            .O(N__18197),
            .I(r_Clock_Count_7_adj_2430));
    LocalMux I__1777 (
            .O(N__18192),
            .I(r_Clock_Count_7_adj_2430));
    InMux I__1776 (
            .O(N__18181),
            .I(N__18167));
    InMux I__1775 (
            .O(N__18180),
            .I(N__18167));
    InMux I__1774 (
            .O(N__18179),
            .I(N__18167));
    InMux I__1773 (
            .O(N__18178),
            .I(N__18156));
    InMux I__1772 (
            .O(N__18177),
            .I(N__18156));
    InMux I__1771 (
            .O(N__18176),
            .I(N__18156));
    InMux I__1770 (
            .O(N__18175),
            .I(N__18156));
    InMux I__1769 (
            .O(N__18174),
            .I(N__18156));
    LocalMux I__1768 (
            .O(N__18167),
            .I(n16852));
    LocalMux I__1767 (
            .O(N__18156),
            .I(n16852));
    InMux I__1766 (
            .O(N__18151),
            .I(\c0.rx.n15674 ));
    InMux I__1765 (
            .O(N__18148),
            .I(N__18145));
    LocalMux I__1764 (
            .O(N__18145),
            .I(n16855));
    InMux I__1763 (
            .O(N__18142),
            .I(N__18137));
    InMux I__1762 (
            .O(N__18141),
            .I(N__18132));
    InMux I__1761 (
            .O(N__18140),
            .I(N__18132));
    LocalMux I__1760 (
            .O(N__18137),
            .I(\c0.FRAME_MATCHER_state_15 ));
    LocalMux I__1759 (
            .O(N__18132),
            .I(\c0.FRAME_MATCHER_state_15 ));
    SRMux I__1758 (
            .O(N__18127),
            .I(N__18124));
    LocalMux I__1757 (
            .O(N__18124),
            .I(\c0.n16349 ));
    CascadeMux I__1756 (
            .O(N__18121),
            .I(n1651_cascade_));
    CascadeMux I__1755 (
            .O(N__18118),
            .I(\c0.rx.r_SM_Main_2_N_2096_0_cascade_ ));
    InMux I__1754 (
            .O(N__18115),
            .I(N__18112));
    LocalMux I__1753 (
            .O(N__18112),
            .I(n6_adj_2461));
    InMux I__1752 (
            .O(N__18109),
            .I(N__18106));
    LocalMux I__1751 (
            .O(N__18106),
            .I(n17641));
    CascadeMux I__1750 (
            .O(N__18103),
            .I(n17144_cascade_));
    InMux I__1749 (
            .O(N__18100),
            .I(N__18088));
    InMux I__1748 (
            .O(N__18099),
            .I(N__18088));
    InMux I__1747 (
            .O(N__18098),
            .I(N__18088));
    InMux I__1746 (
            .O(N__18097),
            .I(N__18081));
    InMux I__1745 (
            .O(N__18096),
            .I(N__18081));
    InMux I__1744 (
            .O(N__18095),
            .I(N__18081));
    LocalMux I__1743 (
            .O(N__18088),
            .I(n16828));
    LocalMux I__1742 (
            .O(N__18081),
            .I(n16828));
    InMux I__1741 (
            .O(N__18076),
            .I(bfn_2_32_0_));
    InMux I__1740 (
            .O(N__18073),
            .I(\c0.rx.n15668 ));
    InMux I__1739 (
            .O(N__18070),
            .I(N__18066));
    InMux I__1738 (
            .O(N__18069),
            .I(N__18062));
    LocalMux I__1737 (
            .O(N__18066),
            .I(N__18059));
    InMux I__1736 (
            .O(N__18065),
            .I(N__18056));
    LocalMux I__1735 (
            .O(N__18062),
            .I(r_Clock_Count_2_adj_2435));
    Odrv4 I__1734 (
            .O(N__18059),
            .I(r_Clock_Count_2_adj_2435));
    LocalMux I__1733 (
            .O(N__18056),
            .I(r_Clock_Count_2_adj_2435));
    InMux I__1732 (
            .O(N__18049),
            .I(N__18046));
    LocalMux I__1731 (
            .O(N__18046),
            .I(N__18043));
    Odrv4 I__1730 (
            .O(N__18043),
            .I(n16860));
    InMux I__1729 (
            .O(N__18040),
            .I(\c0.rx.n15669 ));
    InMux I__1728 (
            .O(N__18037),
            .I(\c0.rx.n15670 ));
    InMux I__1727 (
            .O(N__18034),
            .I(N__18031));
    LocalMux I__1726 (
            .O(N__18031),
            .I(n17494));
    InMux I__1725 (
            .O(N__18028),
            .I(N__18025));
    LocalMux I__1724 (
            .O(N__18025),
            .I(n17542));
    CascadeMux I__1723 (
            .O(N__18022),
            .I(N__18019));
    InMux I__1722 (
            .O(N__18019),
            .I(N__18016));
    LocalMux I__1721 (
            .O(N__18016),
            .I(n17484));
    CascadeMux I__1720 (
            .O(N__18013),
            .I(n17_adj_2416_cascade_));
    InMux I__1719 (
            .O(N__18010),
            .I(N__18005));
    InMux I__1718 (
            .O(N__18009),
            .I(N__18000));
    InMux I__1717 (
            .O(N__18008),
            .I(N__18000));
    LocalMux I__1716 (
            .O(N__18005),
            .I(r_Clock_Count_2));
    LocalMux I__1715 (
            .O(N__18000),
            .I(r_Clock_Count_2));
    CascadeMux I__1714 (
            .O(N__17995),
            .I(N__17990));
    InMux I__1713 (
            .O(N__17994),
            .I(N__17987));
    InMux I__1712 (
            .O(N__17993),
            .I(N__17982));
    InMux I__1711 (
            .O(N__17990),
            .I(N__17982));
    LocalMux I__1710 (
            .O(N__17987),
            .I(r_Clock_Count_3));
    LocalMux I__1709 (
            .O(N__17982),
            .I(r_Clock_Count_3));
    InMux I__1708 (
            .O(N__17977),
            .I(N__17972));
    InMux I__1707 (
            .O(N__17976),
            .I(N__17967));
    InMux I__1706 (
            .O(N__17975),
            .I(N__17967));
    LocalMux I__1705 (
            .O(N__17972),
            .I(r_Clock_Count_0));
    LocalMux I__1704 (
            .O(N__17967),
            .I(r_Clock_Count_0));
    InMux I__1703 (
            .O(N__17962),
            .I(N__17957));
    InMux I__1702 (
            .O(N__17961),
            .I(N__17954));
    InMux I__1701 (
            .O(N__17960),
            .I(N__17951));
    LocalMux I__1700 (
            .O(N__17957),
            .I(r_Clock_Count_5));
    LocalMux I__1699 (
            .O(N__17954),
            .I(r_Clock_Count_5));
    LocalMux I__1698 (
            .O(N__17951),
            .I(r_Clock_Count_5));
    CascadeMux I__1697 (
            .O(N__17944),
            .I(\c0.tx.n10_cascade_ ));
    InMux I__1696 (
            .O(N__17941),
            .I(N__17935));
    InMux I__1695 (
            .O(N__17940),
            .I(N__17928));
    InMux I__1694 (
            .O(N__17939),
            .I(N__17928));
    InMux I__1693 (
            .O(N__17938),
            .I(N__17928));
    LocalMux I__1692 (
            .O(N__17935),
            .I(n16863));
    LocalMux I__1691 (
            .O(N__17928),
            .I(n16863));
    CascadeMux I__1690 (
            .O(N__17923),
            .I(n16863_cascade_));
    InMux I__1689 (
            .O(N__17920),
            .I(N__17917));
    LocalMux I__1688 (
            .O(N__17917),
            .I(n9403));
    CascadeMux I__1687 (
            .O(N__17914),
            .I(n17140_cascade_));
    InMux I__1686 (
            .O(N__17911),
            .I(N__17899));
    InMux I__1685 (
            .O(N__17910),
            .I(N__17899));
    InMux I__1684 (
            .O(N__17909),
            .I(N__17899));
    InMux I__1683 (
            .O(N__17908),
            .I(N__17892));
    InMux I__1682 (
            .O(N__17907),
            .I(N__17892));
    InMux I__1681 (
            .O(N__17906),
            .I(N__17892));
    LocalMux I__1680 (
            .O(N__17899),
            .I(n16817));
    LocalMux I__1679 (
            .O(N__17892),
            .I(n16817));
    InMux I__1678 (
            .O(N__17887),
            .I(N__17882));
    InMux I__1677 (
            .O(N__17886),
            .I(N__17877));
    InMux I__1676 (
            .O(N__17885),
            .I(N__17877));
    LocalMux I__1675 (
            .O(N__17882),
            .I(n12_adj_2410));
    LocalMux I__1674 (
            .O(N__17877),
            .I(n12_adj_2410));
    InMux I__1673 (
            .O(N__17872),
            .I(N__17867));
    InMux I__1672 (
            .O(N__17871),
            .I(N__17864));
    InMux I__1671 (
            .O(N__17870),
            .I(N__17861));
    LocalMux I__1670 (
            .O(N__17867),
            .I(r_Clock_Count_5_adj_2449));
    LocalMux I__1669 (
            .O(N__17864),
            .I(r_Clock_Count_5_adj_2449));
    LocalMux I__1668 (
            .O(N__17861),
            .I(r_Clock_Count_5_adj_2449));
    CascadeMux I__1667 (
            .O(N__17854),
            .I(N__17851));
    InMux I__1666 (
            .O(N__17851),
            .I(N__17846));
    InMux I__1665 (
            .O(N__17850),
            .I(N__17843));
    InMux I__1664 (
            .O(N__17849),
            .I(N__17840));
    LocalMux I__1663 (
            .O(N__17846),
            .I(r_Clock_Count_1_adj_2453));
    LocalMux I__1662 (
            .O(N__17843),
            .I(r_Clock_Count_1_adj_2453));
    LocalMux I__1661 (
            .O(N__17840),
            .I(r_Clock_Count_1_adj_2453));
    InMux I__1660 (
            .O(N__17833),
            .I(N__17830));
    LocalMux I__1659 (
            .O(N__17830),
            .I(\c0.tx2.n10 ));
    CascadeMux I__1658 (
            .O(N__17827),
            .I(N__17824));
    InMux I__1657 (
            .O(N__17824),
            .I(N__17820));
    InMux I__1656 (
            .O(N__17823),
            .I(N__17817));
    LocalMux I__1655 (
            .O(N__17820),
            .I(n15837));
    LocalMux I__1654 (
            .O(N__17817),
            .I(n15837));
    CascadeMux I__1653 (
            .O(N__17812),
            .I(n15837_cascade_));
    CascadeMux I__1652 (
            .O(N__17809),
            .I(r_SM_Main_2_N_2033_1_cascade_));
    InMux I__1651 (
            .O(N__17806),
            .I(N__17799));
    InMux I__1650 (
            .O(N__17805),
            .I(N__17796));
    InMux I__1649 (
            .O(N__17804),
            .I(N__17789));
    InMux I__1648 (
            .O(N__17803),
            .I(N__17789));
    InMux I__1647 (
            .O(N__17802),
            .I(N__17789));
    LocalMux I__1646 (
            .O(N__17799),
            .I(r_Clock_Count_7_adj_2447));
    LocalMux I__1645 (
            .O(N__17796),
            .I(r_Clock_Count_7_adj_2447));
    LocalMux I__1644 (
            .O(N__17789),
            .I(r_Clock_Count_7_adj_2447));
    InMux I__1643 (
            .O(N__17782),
            .I(N__17773));
    InMux I__1642 (
            .O(N__17781),
            .I(N__17773));
    InMux I__1641 (
            .O(N__17780),
            .I(N__17766));
    InMux I__1640 (
            .O(N__17779),
            .I(N__17766));
    InMux I__1639 (
            .O(N__17778),
            .I(N__17766));
    LocalMux I__1638 (
            .O(N__17773),
            .I(r_Clock_Count_8_adj_2446));
    LocalMux I__1637 (
            .O(N__17766),
            .I(r_Clock_Count_8_adj_2446));
    InMux I__1636 (
            .O(N__17761),
            .I(N__17757));
    InMux I__1635 (
            .O(N__17760),
            .I(N__17754));
    LocalMux I__1634 (
            .O(N__17757),
            .I(n9929));
    LocalMux I__1633 (
            .O(N__17754),
            .I(n9929));
    CascadeMux I__1632 (
            .O(N__17749),
            .I(N__17745));
    InMux I__1631 (
            .O(N__17748),
            .I(N__17739));
    InMux I__1630 (
            .O(N__17745),
            .I(N__17739));
    InMux I__1629 (
            .O(N__17744),
            .I(N__17736));
    LocalMux I__1628 (
            .O(N__17739),
            .I(blink_counter_23));
    LocalMux I__1627 (
            .O(N__17736),
            .I(blink_counter_23));
    InMux I__1626 (
            .O(N__17731),
            .I(n15612));
    CascadeMux I__1625 (
            .O(N__17728),
            .I(N__17725));
    InMux I__1624 (
            .O(N__17725),
            .I(N__17718));
    InMux I__1623 (
            .O(N__17724),
            .I(N__17718));
    InMux I__1622 (
            .O(N__17723),
            .I(N__17715));
    LocalMux I__1621 (
            .O(N__17718),
            .I(blink_counter_24));
    LocalMux I__1620 (
            .O(N__17715),
            .I(blink_counter_24));
    InMux I__1619 (
            .O(N__17710),
            .I(bfn_2_28_0_));
    InMux I__1618 (
            .O(N__17707),
            .I(n15614));
    InMux I__1617 (
            .O(N__17704),
            .I(N__17700));
    InMux I__1616 (
            .O(N__17703),
            .I(N__17697));
    LocalMux I__1615 (
            .O(N__17700),
            .I(blink_counter_25));
    LocalMux I__1614 (
            .O(N__17697),
            .I(blink_counter_25));
    InMux I__1613 (
            .O(N__17692),
            .I(N__17689));
    LocalMux I__1612 (
            .O(N__17689),
            .I(n17570));
    InMux I__1611 (
            .O(N__17686),
            .I(N__17683));
    LocalMux I__1610 (
            .O(N__17683),
            .I(n17629));
    InMux I__1609 (
            .O(N__17680),
            .I(N__17677));
    LocalMux I__1608 (
            .O(N__17677),
            .I(n17504));
    InMux I__1607 (
            .O(N__17674),
            .I(N__17669));
    InMux I__1606 (
            .O(N__17673),
            .I(N__17664));
    InMux I__1605 (
            .O(N__17672),
            .I(N__17664));
    LocalMux I__1604 (
            .O(N__17669),
            .I(r_Clock_Count_2_adj_2452));
    LocalMux I__1603 (
            .O(N__17664),
            .I(r_Clock_Count_2_adj_2452));
    InMux I__1602 (
            .O(N__17659),
            .I(N__17654));
    InMux I__1601 (
            .O(N__17658),
            .I(N__17651));
    InMux I__1600 (
            .O(N__17657),
            .I(N__17648));
    LocalMux I__1599 (
            .O(N__17654),
            .I(r_Clock_Count_3_adj_2451));
    LocalMux I__1598 (
            .O(N__17651),
            .I(r_Clock_Count_3_adj_2451));
    LocalMux I__1597 (
            .O(N__17648),
            .I(r_Clock_Count_3_adj_2451));
    InMux I__1596 (
            .O(N__17641),
            .I(n15603));
    InMux I__1595 (
            .O(N__17638),
            .I(N__17635));
    LocalMux I__1594 (
            .O(N__17635),
            .I(n11));
    InMux I__1593 (
            .O(N__17632),
            .I(n15604));
    InMux I__1592 (
            .O(N__17629),
            .I(N__17626));
    LocalMux I__1591 (
            .O(N__17626),
            .I(n10_adj_2420));
    InMux I__1590 (
            .O(N__17623),
            .I(bfn_2_27_0_));
    InMux I__1589 (
            .O(N__17620),
            .I(N__17617));
    LocalMux I__1588 (
            .O(N__17617),
            .I(n9));
    InMux I__1587 (
            .O(N__17614),
            .I(n15606));
    InMux I__1586 (
            .O(N__17611),
            .I(N__17608));
    LocalMux I__1585 (
            .O(N__17608),
            .I(n8));
    InMux I__1584 (
            .O(N__17605),
            .I(n15607));
    InMux I__1583 (
            .O(N__17602),
            .I(N__17599));
    LocalMux I__1582 (
            .O(N__17599),
            .I(n7));
    InMux I__1581 (
            .O(N__17596),
            .I(n15608));
    InMux I__1580 (
            .O(N__17593),
            .I(N__17590));
    LocalMux I__1579 (
            .O(N__17590),
            .I(n6_adj_2421));
    InMux I__1578 (
            .O(N__17587),
            .I(n15609));
    InMux I__1577 (
            .O(N__17584),
            .I(N__17578));
    InMux I__1576 (
            .O(N__17583),
            .I(N__17578));
    LocalMux I__1575 (
            .O(N__17578),
            .I(N__17574));
    InMux I__1574 (
            .O(N__17577),
            .I(N__17571));
    Odrv4 I__1573 (
            .O(N__17574),
            .I(blink_counter_21));
    LocalMux I__1572 (
            .O(N__17571),
            .I(blink_counter_21));
    InMux I__1571 (
            .O(N__17566),
            .I(n15610));
    InMux I__1570 (
            .O(N__17563),
            .I(N__17556));
    InMux I__1569 (
            .O(N__17562),
            .I(N__17556));
    InMux I__1568 (
            .O(N__17561),
            .I(N__17553));
    LocalMux I__1567 (
            .O(N__17556),
            .I(blink_counter_22));
    LocalMux I__1566 (
            .O(N__17553),
            .I(blink_counter_22));
    InMux I__1565 (
            .O(N__17548),
            .I(n15611));
    InMux I__1564 (
            .O(N__17545),
            .I(N__17542));
    LocalMux I__1563 (
            .O(N__17542),
            .I(n20));
    InMux I__1562 (
            .O(N__17539),
            .I(n15595));
    InMux I__1561 (
            .O(N__17536),
            .I(N__17533));
    LocalMux I__1560 (
            .O(N__17533),
            .I(n19));
    InMux I__1559 (
            .O(N__17530),
            .I(n15596));
    InMux I__1558 (
            .O(N__17527),
            .I(N__17524));
    LocalMux I__1557 (
            .O(N__17524),
            .I(n18));
    InMux I__1556 (
            .O(N__17521),
            .I(bfn_2_26_0_));
    InMux I__1555 (
            .O(N__17518),
            .I(N__17515));
    LocalMux I__1554 (
            .O(N__17515),
            .I(n17_adj_2422));
    InMux I__1553 (
            .O(N__17512),
            .I(n15598));
    InMux I__1552 (
            .O(N__17509),
            .I(N__17506));
    LocalMux I__1551 (
            .O(N__17506),
            .I(n16));
    InMux I__1550 (
            .O(N__17503),
            .I(n15599));
    InMux I__1549 (
            .O(N__17500),
            .I(N__17497));
    LocalMux I__1548 (
            .O(N__17497),
            .I(n15));
    InMux I__1547 (
            .O(N__17494),
            .I(n15600));
    InMux I__1546 (
            .O(N__17491),
            .I(N__17488));
    LocalMux I__1545 (
            .O(N__17488),
            .I(n14_adj_2424));
    InMux I__1544 (
            .O(N__17485),
            .I(n15601));
    InMux I__1543 (
            .O(N__17482),
            .I(N__17479));
    LocalMux I__1542 (
            .O(N__17479),
            .I(n13));
    InMux I__1541 (
            .O(N__17476),
            .I(n15602));
    InMux I__1540 (
            .O(N__17473),
            .I(N__17470));
    LocalMux I__1539 (
            .O(N__17470),
            .I(n12_adj_2419));
    InMux I__1538 (
            .O(N__17467),
            .I(N__17464));
    LocalMux I__1537 (
            .O(N__17464),
            .I(n26));
    InMux I__1536 (
            .O(N__17461),
            .I(bfn_2_25_0_));
    InMux I__1535 (
            .O(N__17458),
            .I(N__17455));
    LocalMux I__1534 (
            .O(N__17455),
            .I(n25));
    InMux I__1533 (
            .O(N__17452),
            .I(n15590));
    InMux I__1532 (
            .O(N__17449),
            .I(N__17446));
    LocalMux I__1531 (
            .O(N__17446),
            .I(n24));
    InMux I__1530 (
            .O(N__17443),
            .I(n15591));
    InMux I__1529 (
            .O(N__17440),
            .I(N__17437));
    LocalMux I__1528 (
            .O(N__17437),
            .I(n23));
    InMux I__1527 (
            .O(N__17434),
            .I(n15592));
    InMux I__1526 (
            .O(N__17431),
            .I(N__17428));
    LocalMux I__1525 (
            .O(N__17428),
            .I(n22));
    InMux I__1524 (
            .O(N__17425),
            .I(n15593));
    InMux I__1523 (
            .O(N__17422),
            .I(N__17419));
    LocalMux I__1522 (
            .O(N__17419),
            .I(n21));
    InMux I__1521 (
            .O(N__17416),
            .I(n15594));
    InMux I__1520 (
            .O(N__17413),
            .I(N__17404));
    InMux I__1519 (
            .O(N__17412),
            .I(N__17404));
    InMux I__1518 (
            .O(N__17411),
            .I(N__17404));
    LocalMux I__1517 (
            .O(N__17404),
            .I(\c0.FRAME_MATCHER_state_7 ));
    SRMux I__1516 (
            .O(N__17401),
            .I(N__17398));
    LocalMux I__1515 (
            .O(N__17398),
            .I(N__17395));
    Odrv4 I__1514 (
            .O(N__17395),
            .I(\c0.n16443 ));
    InMux I__1513 (
            .O(N__17392),
            .I(N__17387));
    InMux I__1512 (
            .O(N__17391),
            .I(N__17382));
    InMux I__1511 (
            .O(N__17390),
            .I(N__17382));
    LocalMux I__1510 (
            .O(N__17387),
            .I(\c0.FRAME_MATCHER_state_13 ));
    LocalMux I__1509 (
            .O(N__17382),
            .I(\c0.FRAME_MATCHER_state_13 ));
    SRMux I__1508 (
            .O(N__17377),
            .I(N__17374));
    LocalMux I__1507 (
            .O(N__17374),
            .I(N__17371));
    Span4Mux_s1_h I__1506 (
            .O(N__17371),
            .I(N__17368));
    Span4Mux_h I__1505 (
            .O(N__17368),
            .I(N__17365));
    Odrv4 I__1504 (
            .O(N__17365),
            .I(\c0.n16447 ));
    CascadeMux I__1503 (
            .O(N__17362),
            .I(N__17358));
    InMux I__1502 (
            .O(N__17361),
            .I(N__17353));
    InMux I__1501 (
            .O(N__17358),
            .I(N__17353));
    LocalMux I__1500 (
            .O(N__17353),
            .I(N__17349));
    InMux I__1499 (
            .O(N__17352),
            .I(N__17346));
    Span4Mux_h I__1498 (
            .O(N__17349),
            .I(N__17343));
    LocalMux I__1497 (
            .O(N__17346),
            .I(\c0.FRAME_MATCHER_state_11 ));
    Odrv4 I__1496 (
            .O(N__17343),
            .I(\c0.FRAME_MATCHER_state_11 ));
    SRMux I__1495 (
            .O(N__17338),
            .I(N__17335));
    LocalMux I__1494 (
            .O(N__17335),
            .I(\c0.n16451 ));
    SRMux I__1493 (
            .O(N__17332),
            .I(N__17329));
    LocalMux I__1492 (
            .O(N__17329),
            .I(N__17326));
    Odrv12 I__1491 (
            .O(N__17326),
            .I(\c0.n16445 ));
    CascadeMux I__1490 (
            .O(N__17323),
            .I(\c0.rx.r_SM_Main_2_N_2090_2_cascade_ ));
    InMux I__1489 (
            .O(N__17320),
            .I(N__17317));
    LocalMux I__1488 (
            .O(N__17317),
            .I(n17631));
    CascadeMux I__1487 (
            .O(N__17314),
            .I(n16810_cascade_));
    CascadeMux I__1486 (
            .O(N__17311),
            .I(\c0.rx.n13452_cascade_ ));
    InMux I__1485 (
            .O(N__17308),
            .I(N__17305));
    LocalMux I__1484 (
            .O(N__17305),
            .I(n16867));
    InMux I__1483 (
            .O(N__17302),
            .I(N__17296));
    InMux I__1482 (
            .O(N__17301),
            .I(N__17296));
    LocalMux I__1481 (
            .O(N__17296),
            .I(n17222));
    SRMux I__1480 (
            .O(N__17293),
            .I(N__17290));
    LocalMux I__1479 (
            .O(N__17290),
            .I(N__17287));
    Span4Mux_s3_v I__1478 (
            .O(N__17287),
            .I(N__17284));
    Span4Mux_s1_h I__1477 (
            .O(N__17284),
            .I(N__17281));
    Odrv4 I__1476 (
            .O(N__17281),
            .I(\c0.rx.n16850 ));
    InMux I__1475 (
            .O(N__17278),
            .I(\c0.tx.n15662 ));
    InMux I__1474 (
            .O(N__17275),
            .I(\c0.tx.n15663 ));
    InMux I__1473 (
            .O(N__17272),
            .I(\c0.tx.n15664 ));
    InMux I__1472 (
            .O(N__17269),
            .I(\c0.tx.n15665 ));
    InMux I__1471 (
            .O(N__17266),
            .I(\c0.tx.n15666 ));
    InMux I__1470 (
            .O(N__17263),
            .I(bfn_1_31_0_));
    CascadeMux I__1469 (
            .O(N__17260),
            .I(n17537_cascade_));
    InMux I__1468 (
            .O(N__17257),
            .I(bfn_1_29_0_));
    InMux I__1467 (
            .O(N__17254),
            .I(N__17251));
    LocalMux I__1466 (
            .O(N__17251),
            .I(n17640));
    InMux I__1465 (
            .O(N__17248),
            .I(N__17243));
    InMux I__1464 (
            .O(N__17247),
            .I(N__17240));
    InMux I__1463 (
            .O(N__17246),
            .I(N__17237));
    LocalMux I__1462 (
            .O(N__17243),
            .I(n16824));
    LocalMux I__1461 (
            .O(N__17240),
            .I(n16824));
    LocalMux I__1460 (
            .O(N__17237),
            .I(n16824));
    InMux I__1459 (
            .O(N__17230),
            .I(N__17227));
    LocalMux I__1458 (
            .O(N__17227),
            .I(n10_adj_2412));
    InMux I__1457 (
            .O(N__17224),
            .I(N__17221));
    LocalMux I__1456 (
            .O(N__17221),
            .I(n17458));
    InMux I__1455 (
            .O(N__17218),
            .I(bfn_1_30_0_));
    InMux I__1454 (
            .O(N__17215),
            .I(\c0.tx.n15660 ));
    InMux I__1453 (
            .O(N__17212),
            .I(\c0.tx.n15661 ));
    InMux I__1452 (
            .O(N__17209),
            .I(N__17206));
    LocalMux I__1451 (
            .O(N__17206),
            .I(n17298));
    InMux I__1450 (
            .O(N__17203),
            .I(bfn_1_28_0_));
    InMux I__1449 (
            .O(N__17200),
            .I(\c0.tx2.n15675 ));
    InMux I__1448 (
            .O(N__17197),
            .I(\c0.tx2.n15676 ));
    InMux I__1447 (
            .O(N__17194),
            .I(N__17191));
    LocalMux I__1446 (
            .O(N__17191),
            .I(n17457));
    InMux I__1445 (
            .O(N__17188),
            .I(\c0.tx2.n15677 ));
    InMux I__1444 (
            .O(N__17185),
            .I(\c0.tx2.n15678 ));
    InMux I__1443 (
            .O(N__17182),
            .I(\c0.tx2.n15679 ));
    InMux I__1442 (
            .O(N__17179),
            .I(\c0.tx2.n15680 ));
    InMux I__1441 (
            .O(N__17176),
            .I(\c0.tx2.n15681 ));
    CascadeMux I__1440 (
            .O(N__17173),
            .I(n17299_cascade_));
    IoInMux I__1439 (
            .O(N__17170),
            .I(N__17167));
    LocalMux I__1438 (
            .O(N__17167),
            .I(N__17164));
    Span4Mux_s1_v I__1437 (
            .O(N__17164),
            .I(N__17161));
    Span4Mux_v I__1436 (
            .O(N__17161),
            .I(N__17158));
    Odrv4 I__1435 (
            .O(N__17158),
            .I(LED_c));
    IoInMux I__1434 (
            .O(N__17155),
            .I(N__17152));
    LocalMux I__1433 (
            .O(N__17152),
            .I(tx2_enable));
    IoInMux I__1432 (
            .O(N__17149),
            .I(N__17146));
    LocalMux I__1431 (
            .O(N__17146),
            .I(N__17143));
    IoSpan4Mux I__1430 (
            .O(N__17143),
            .I(N__17140));
    IoSpan4Mux I__1429 (
            .O(N__17140),
            .I(N__17137));
    IoSpan4Mux I__1428 (
            .O(N__17137),
            .I(N__17134));
    Odrv4 I__1427 (
            .O(N__17134),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_13_29_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_29_0_));
    defparam IN_MUX_bfv_13_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_30_0_ (
            .carryinitin(n15566),
            .carryinitout(bfn_13_30_0_));
    defparam IN_MUX_bfv_13_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_31_0_ (
            .carryinitin(n15574),
            .carryinitout(bfn_13_31_0_));
    defparam IN_MUX_bfv_13_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_32_0_ (
            .carryinitin(n15582),
            .carryinitout(bfn_13_32_0_));
    defparam IN_MUX_bfv_13_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_25_0_));
    defparam IN_MUX_bfv_13_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_26_0_ (
            .carryinitin(n15535),
            .carryinitout(bfn_13_26_0_));
    defparam IN_MUX_bfv_13_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_27_0_ (
            .carryinitin(n15543),
            .carryinitout(bfn_13_27_0_));
    defparam IN_MUX_bfv_13_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_28_0_ (
            .carryinitin(n15551),
            .carryinitout(bfn_13_28_0_));
    defparam IN_MUX_bfv_1_28_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_28_0_));
    defparam IN_MUX_bfv_1_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_29_0_ (
            .carryinitin(\c0.tx2.n15682 ),
            .carryinitout(bfn_1_29_0_));
    defparam IN_MUX_bfv_1_30_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_30_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_30_0_));
    defparam IN_MUX_bfv_1_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_31_0_ (
            .carryinitin(\c0.tx.n15667 ),
            .carryinitout(bfn_1_31_0_));
    defparam IN_MUX_bfv_2_32_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_32_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_32_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_4_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_22_0_));
    defparam IN_MUX_bfv_4_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_23_0_ (
            .carryinitin(\c0.n15629 ),
            .carryinitout(bfn_4_23_0_));
    defparam IN_MUX_bfv_4_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_24_0_ (
            .carryinitin(\c0.n15637 ),
            .carryinitout(bfn_4_24_0_));
    defparam IN_MUX_bfv_4_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_25_0_ (
            .carryinitin(\c0.n15645 ),
            .carryinitout(bfn_4_25_0_));
    defparam IN_MUX_bfv_5_31_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_31_0_));
    defparam IN_MUX_bfv_5_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_32_0_ (
            .carryinitin(\c0.n15521 ),
            .carryinitout(bfn_5_32_0_));
    defparam IN_MUX_bfv_6_30_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_30_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_30_0_));
    defparam IN_MUX_bfv_2_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_25_0_));
    defparam IN_MUX_bfv_2_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_26_0_ (
            .carryinitin(n15597),
            .carryinitout(bfn_2_26_0_));
    defparam IN_MUX_bfv_2_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_27_0_ (
            .carryinitin(n15605),
            .carryinitout(bfn_2_27_0_));
    defparam IN_MUX_bfv_2_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_28_0_ (
            .carryinitin(n15613),
            .carryinitout(bfn_2_28_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__17149),
            .GLOBALBUFFEROUTPUT(CLK_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i11_LC_1_17_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i11_LC_1_17_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i11_LC_1_17_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.FRAME_MATCHER_state_i11_LC_1_17_0  (
            .in0(N__34663),
            .in1(N__17352),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_state_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50377),
            .ce(),
            .sr(N__17338));
    defparam \c0.FRAME_MATCHER_state_i8_LC_1_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i8_LC_1_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i8_LC_1_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i8_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(N__34655),
            .in2(_gnd_net_),
            .in3(N__30110),
            .lcout(\c0.FRAME_MATCHER_state_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50378),
            .ce(),
            .sr(N__17332));
    defparam \c0.FRAME_MATCHER_state_i13_LC_1_19_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i13_LC_1_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i13_LC_1_19_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.FRAME_MATCHER_state_i13_LC_1_19_0  (
            .in0(N__34660),
            .in1(N__17392),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_state_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50380),
            .ce(),
            .sr(N__17377));
    defparam \c0.FRAME_MATCHER_i_i23_LC_1_20_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i23_LC_1_20_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i23_LC_1_20_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i23_LC_1_20_0  (
            .in0(N__33226),
            .in1(N__33004),
            .in2(_gnd_net_),
            .in3(N__19180),
            .lcout(\c0.FRAME_MATCHER_i_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50383),
            .ce(),
            .sr(N__20206));
    defparam \c0.FRAME_MATCHER_i_i20_LC_1_21_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i20_LC_1_21_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i20_LC_1_21_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i20_LC_1_21_0  (
            .in0(N__33257),
            .in1(N__32911),
            .in2(_gnd_net_),
            .in3(N__19228),
            .lcout(\c0.FRAME_MATCHER_i_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50387),
            .ce(),
            .sr(N__20374));
    defparam \c0.FRAME_MATCHER_i_i22_LC_1_22_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i22_LC_1_22_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i22_LC_1_22_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i22_LC_1_22_0  (
            .in0(N__33266),
            .in1(N__33003),
            .in2(_gnd_net_),
            .in3(N__19195),
            .lcout(\c0.FRAME_MATCHER_i_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50393),
            .ce(),
            .sr(N__20332));
    defparam \c0.FRAME_MATCHER_i_i8_LC_1_23_5 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i8_LC_1_23_5 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i8_LC_1_23_5 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i8_LC_1_23_5  (
            .in0(N__32999),
            .in1(N__33268),
            .in2(_gnd_net_),
            .in3(N__18964),
            .lcout(\c0.FRAME_MATCHER_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50400),
            .ce(),
            .sr(N__18802));
    defparam \c0.FRAME_MATCHER_i_i26_LC_1_24_7 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i26_LC_1_24_7 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i26_LC_1_24_7 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i26_LC_1_24_7  (
            .in0(N__33000),
            .in1(N__33269),
            .in2(_gnd_net_),
            .in3(N__19141),
            .lcout(\c0.FRAME_MATCHER_i_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50406),
            .ce(),
            .sr(N__20302));
    defparam \c0.FRAME_MATCHER_i_i1_LC_1_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i1_LC_1_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i1_LC_1_25_0 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \c0.FRAME_MATCHER_i_i1_LC_1_25_0  (
            .in0(_gnd_net_),
            .in1(N__33279),
            .in2(N__18880),
            .in3(N__33001),
            .lcout(\c0.FRAME_MATCHER_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50413),
            .ce(),
            .sr(N__18901));
    defparam \c0.FRAME_MATCHER_i_i27_LC_1_26_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i27_LC_1_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i27_LC_1_26_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i27_LC_1_26_0  (
            .in0(N__33280),
            .in1(N__33002),
            .in2(_gnd_net_),
            .in3(N__19126),
            .lcout(\c0.FRAME_MATCHER_i_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50423),
            .ce(),
            .sr(N__20272));
    defparam \c0.tx2.r_Clock_Count__i3_LC_1_27_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i3_LC_1_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i3_LC_1_27_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.tx2.r_Clock_Count__i3_LC_1_27_0  (
            .in0(N__17194),
            .in1(N__31532),
            .in2(_gnd_net_),
            .in3(N__17659),
            .lcout(r_Clock_Count_3_adj_2451),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50431),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i14822_4_lut_LC_1_27_1 .C_ON=1'b0;
    defparam \c0.rx.i14822_4_lut_LC_1_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i14822_4_lut_LC_1_27_1 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \c0.rx.i14822_4_lut_LC_1_27_1  (
            .in0(N__30779),
            .in1(N__30852),
            .in2(N__33874),
            .in3(N__18412),
            .lcout(n17260),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14861_4_lut_LC_1_27_2.C_ON=1'b0;
    defparam i14861_4_lut_LC_1_27_2.SEQ_MODE=4'b0000;
    defparam i14861_4_lut_LC_1_27_2.LUT_INIT=16'b1111111011000100;
    LogicCell40 i14861_4_lut_LC_1_27_2 (
            .in0(N__17563),
            .in1(N__17748),
            .in2(N__17728),
            .in3(N__17584),
            .lcout(),
            .ltout(n17299_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14862_3_lut_LC_1_27_3.C_ON=1'b0;
    defparam i14862_3_lut_LC_1_27_3.SEQ_MODE=4'b0000;
    defparam i14862_3_lut_LC_1_27_3.LUT_INIT=16'b0000101001011111;
    LogicCell40 i14862_3_lut_LC_1_27_3 (
            .in0(N__17704),
            .in1(_gnd_net_),
            .in2(N__17173),
            .in3(N__17209),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i81_LC_1_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i81_LC_1_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i81_LC_1_27_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i81_LC_1_27_4  (
            .in0(N__25602),
            .in1(N__31924),
            .in2(N__23664),
            .in3(N__31137),
            .lcout(\c0.data_in_frame_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50431),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15447_2_lut_3_lut_LC_1_27_5 .C_ON=1'b0;
    defparam \c0.rx.i15447_2_lut_3_lut_LC_1_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15447_2_lut_3_lut_LC_1_27_5 .LUT_INIT=16'b1111111101011111;
    LogicCell40 \c0.rx.i15447_2_lut_3_lut_LC_1_27_5  (
            .in0(N__30780),
            .in1(_gnd_net_),
            .in2(N__33875),
            .in3(N__30853),
            .lcout(\c0.rx.n16850 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_1_27_6 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_1_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_1_27_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_1_27_6  (
            .in0(N__28689),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(tx2_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14860_4_lut_LC_1_27_7.C_ON=1'b0;
    defparam i14860_4_lut_LC_1_27_7.SEQ_MODE=4'b0000;
    defparam i14860_4_lut_LC_1_27_7.LUT_INIT=16'b1011101000100010;
    LogicCell40 i14860_4_lut_LC_1_27_7 (
            .in0(N__17583),
            .in1(N__17724),
            .in2(N__17749),
            .in3(N__17562),
            .lcout(n17298),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_2_lut_LC_1_28_0 .C_ON=1'b1;
    defparam \c0.tx2.add_59_2_lut_LC_1_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_2_lut_LC_1_28_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx2.add_59_2_lut_LC_1_28_0  (
            .in0(N__17906),
            .in1(N__31407),
            .in2(_gnd_net_),
            .in3(N__17203),
            .lcout(n17544),
            .ltout(),
            .carryin(bfn_1_28_0_),
            .carryout(\c0.tx2.n15675 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_3_lut_LC_1_28_1 .C_ON=1'b1;
    defparam \c0.tx2.add_59_3_lut_LC_1_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_3_lut_LC_1_28_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx2.add_59_3_lut_LC_1_28_1  (
            .in0(N__17910),
            .in1(N__17850),
            .in2(_gnd_net_),
            .in3(N__17200),
            .lcout(n17504),
            .ltout(),
            .carryin(\c0.tx2.n15675 ),
            .carryout(\c0.tx2.n15676 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_4_lut_LC_1_28_2 .C_ON=1'b1;
    defparam \c0.tx2.add_59_4_lut_LC_1_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_4_lut_LC_1_28_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx2.add_59_4_lut_LC_1_28_2  (
            .in0(N__17908),
            .in1(N__17674),
            .in2(_gnd_net_),
            .in3(N__17197),
            .lcout(n17570),
            .ltout(),
            .carryin(\c0.tx2.n15676 ),
            .carryout(\c0.tx2.n15677 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_5_lut_LC_1_28_3 .C_ON=1'b1;
    defparam \c0.tx2.add_59_5_lut_LC_1_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_5_lut_LC_1_28_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx2.add_59_5_lut_LC_1_28_3  (
            .in0(N__17909),
            .in1(N__17658),
            .in2(_gnd_net_),
            .in3(N__17188),
            .lcout(n17457),
            .ltout(),
            .carryin(\c0.tx2.n15677 ),
            .carryout(\c0.tx2.n15678 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_6_lut_LC_1_28_4 .C_ON=1'b1;
    defparam \c0.tx2.add_59_6_lut_LC_1_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_6_lut_LC_1_28_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx2.add_59_6_lut_LC_1_28_4  (
            .in0(N__17907),
            .in1(N__19570),
            .in2(_gnd_net_),
            .in3(N__17185),
            .lcout(n17567),
            .ltout(),
            .carryin(\c0.tx2.n15678 ),
            .carryout(\c0.tx2.n15679 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_7_lut_LC_1_28_5 .C_ON=1'b1;
    defparam \c0.tx2.add_59_7_lut_LC_1_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_7_lut_LC_1_28_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx2.add_59_7_lut_LC_1_28_5  (
            .in0(N__17911),
            .in1(N__17871),
            .in2(_gnd_net_),
            .in3(N__17182),
            .lcout(n17629),
            .ltout(),
            .carryin(\c0.tx2.n15679 ),
            .carryout(\c0.tx2.n15680 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_8_lut_LC_1_28_6 .C_ON=1'b1;
    defparam \c0.tx2.add_59_8_lut_LC_1_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_8_lut_LC_1_28_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx2.add_59_8_lut_LC_1_28_6  (
            .in0(N__17246),
            .in1(N__26382),
            .in2(_gnd_net_),
            .in3(N__17179),
            .lcout(n17634),
            .ltout(),
            .carryin(\c0.tx2.n15680 ),
            .carryout(\c0.tx2.n15681 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_9_lut_LC_1_28_7 .C_ON=1'b1;
    defparam \c0.tx2.add_59_9_lut_LC_1_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_9_lut_LC_1_28_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx2.add_59_9_lut_LC_1_28_7  (
            .in0(N__17247),
            .in1(N__17805),
            .in2(_gnd_net_),
            .in3(N__17176),
            .lcout(n17640),
            .ltout(),
            .carryin(\c0.tx2.n15681 ),
            .carryout(\c0.tx2.n15682 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_10_lut_LC_1_29_0 .C_ON=1'b0;
    defparam \c0.tx2.add_59_10_lut_LC_1_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_10_lut_LC_1_29_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx2.add_59_10_lut_LC_1_29_0  (
            .in0(N__17248),
            .in1(N__17781),
            .in2(_gnd_net_),
            .in3(N__17257),
            .lcout(n17458),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i7_LC_1_29_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i7_LC_1_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i7_LC_1_29_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i7_LC_1_29_1  (
            .in0(N__31513),
            .in1(N__17806),
            .in2(_gnd_net_),
            .in3(N__17254),
            .lcout(r_Clock_Count_7_adj_2447),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50447),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_777_LC_1_29_3.C_ON=1'b0;
    defparam i1_4_lut_adj_777_LC_1_29_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_777_LC_1_29_3.LUT_INIT=16'b0000110000001110;
    LogicCell40 i1_4_lut_adj_777_LC_1_29_3 (
            .in0(N__17886),
            .in1(N__17230),
            .in2(N__17827),
            .in3(N__30996),
            .lcout(n16824),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_797_LC_1_29_4.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_797_LC_1_29_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_797_LC_1_29_4.LUT_INIT=16'b0000101000000010;
    LogicCell40 i1_3_lut_4_lut_adj_797_LC_1_29_4 (
            .in0(N__30995),
            .in1(N__17760),
            .in2(N__31514),
            .in3(N__17885),
            .lcout(n10_adj_2412),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_2_lut_LC_1_29_6 .C_ON=1'b0;
    defparam \c0.tx2.i1_2_lut_LC_1_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_2_lut_LC_1_29_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.tx2.i1_2_lut_LC_1_29_6  (
            .in0(N__31481),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30994),
            .lcout(n9403),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_29_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_29_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i8_LC_1_29_7  (
            .in0(N__17782),
            .in1(N__31485),
            .in2(_gnd_net_),
            .in3(N__17224),
            .lcout(r_Clock_Count_8_adj_2446),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50447),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_2_lut_LC_1_30_0 .C_ON=1'b1;
    defparam \c0.tx.add_59_2_lut_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_2_lut_LC_1_30_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_2_lut_LC_1_30_0  (
            .in0(N__18099),
            .in1(N__17977),
            .in2(_gnd_net_),
            .in3(N__17218),
            .lcout(n17542),
            .ltout(),
            .carryin(bfn_1_30_0_),
            .carryout(\c0.tx.n15660 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_3_lut_LC_1_30_1 .C_ON=1'b1;
    defparam \c0.tx.add_59_3_lut_LC_1_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_3_lut_LC_1_30_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_3_lut_LC_1_30_1  (
            .in0(N__18095),
            .in1(N__18676),
            .in2(_gnd_net_),
            .in3(N__17215),
            .lcout(n17461),
            .ltout(),
            .carryin(\c0.tx.n15660 ),
            .carryout(\c0.tx.n15661 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_4_lut_LC_1_30_2 .C_ON=1'b1;
    defparam \c0.tx.add_59_4_lut_LC_1_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_4_lut_LC_1_30_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_4_lut_LC_1_30_2  (
            .in0(N__18100),
            .in1(N__18010),
            .in2(_gnd_net_),
            .in3(N__17212),
            .lcout(n17484),
            .ltout(),
            .carryin(\c0.tx.n15661 ),
            .carryout(\c0.tx.n15662 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_5_lut_LC_1_30_3 .C_ON=1'b1;
    defparam \c0.tx.add_59_5_lut_LC_1_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_5_lut_LC_1_30_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_5_lut_LC_1_30_3  (
            .in0(N__18096),
            .in1(N__17994),
            .in2(_gnd_net_),
            .in3(N__17278),
            .lcout(n17494),
            .ltout(),
            .carryin(\c0.tx.n15662 ),
            .carryout(\c0.tx.n15663 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_6_lut_LC_1_30_4 .C_ON=1'b1;
    defparam \c0.tx.add_59_6_lut_LC_1_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_6_lut_LC_1_30_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_6_lut_LC_1_30_4  (
            .in0(N__18098),
            .in1(N__19723),
            .in2(_gnd_net_),
            .in3(N__17275),
            .lcout(n17573),
            .ltout(),
            .carryin(\c0.tx.n15663 ),
            .carryout(\c0.tx.n15664 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_7_lut_LC_1_30_5 .C_ON=1'b1;
    defparam \c0.tx.add_59_7_lut_LC_1_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_7_lut_LC_1_30_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_7_lut_LC_1_30_5  (
            .in0(N__18097),
            .in1(N__17961),
            .in2(_gnd_net_),
            .in3(N__17272),
            .lcout(n17631),
            .ltout(),
            .carryin(\c0.tx.n15664 ),
            .carryout(\c0.tx.n15665 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_8_lut_LC_1_30_6 .C_ON=1'b1;
    defparam \c0.tx.add_59_8_lut_LC_1_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_8_lut_LC_1_30_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_8_lut_LC_1_30_6  (
            .in0(N__18449),
            .in1(N__19834),
            .in2(_gnd_net_),
            .in3(N__17269),
            .lcout(n17636),
            .ltout(),
            .carryin(\c0.tx.n15665 ),
            .carryout(\c0.tx.n15666 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_9_lut_LC_1_30_7 .C_ON=1'b1;
    defparam \c0.tx.add_59_9_lut_LC_1_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_9_lut_LC_1_30_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_9_lut_LC_1_30_7  (
            .in0(N__18450),
            .in1(N__19863),
            .in2(_gnd_net_),
            .in3(N__17266),
            .lcout(n17641),
            .ltout(),
            .carryin(\c0.tx.n15666 ),
            .carryout(\c0.tx.n15667 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_10_lut_LC_1_31_0 .C_ON=1'b0;
    defparam \c0.tx.add_59_10_lut_LC_1_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_10_lut_LC_1_31_0 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \c0.tx.add_59_10_lut_LC_1_31_0  (
            .in0(N__19792),
            .in1(N__18454),
            .in2(_gnd_net_),
            .in3(N__17263),
            .lcout(),
            .ltout(n17537_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i8_LC_1_31_1 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i8_LC_1_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i8_LC_1_31_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.tx.r_Clock_Count__i8_LC_1_31_1  (
            .in0(N__23969),
            .in1(_gnd_net_),
            .in2(N__17260),
            .in3(N__19793),
            .lcout(r_Clock_Count_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50469),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15303_3_lut_LC_1_31_4 .C_ON=1'b0;
    defparam \c0.rx.i15303_3_lut_LC_1_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15303_3_lut_LC_1_31_4 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \c0.rx.i15303_3_lut_LC_1_31_4  (
            .in0(N__33880),
            .in1(N__33780),
            .in2(_gnd_net_),
            .in3(N__33754),
            .lcout(n17601),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_4_lut_LC_1_31_5 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_4_lut_LC_1_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_4_lut_LC_1_31_5 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \c0.rx.i1_2_lut_4_lut_LC_1_31_5  (
            .in0(N__19679),
            .in1(N__18212),
            .in2(N__18772),
            .in3(N__17941),
            .lcout(\c0.rx.r_SM_Main_2_N_2090_2 ),
            .ltout(\c0.rx.r_SM_Main_2_N_2090_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15361_2_lut_LC_1_31_6 .C_ON=1'b0;
    defparam \c0.rx.i15361_2_lut_LC_1_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15361_2_lut_LC_1_31_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \c0.rx.i15361_2_lut_LC_1_31_6  (
            .in0(N__33881),
            .in1(_gnd_net_),
            .in2(N__17323),
            .in3(_gnd_net_),
            .lcout(n17602),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i5_LC_1_31_7 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i5_LC_1_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i5_LC_1_31_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i5_LC_1_31_7  (
            .in0(N__23968),
            .in1(N__17962),
            .in2(_gnd_net_),
            .in3(N__17320),
            .lcout(r_Clock_Count_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50469),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_796_LC_1_32_0.C_ON=1'b0;
    defparam i1_4_lut_adj_796_LC_1_32_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_796_LC_1_32_0.LUT_INIT=16'b1111000010110000;
    LogicCell40 i1_4_lut_adj_796_LC_1_32_0 (
            .in0(N__17302),
            .in1(N__17939),
            .in2(N__33885),
            .in3(N__18770),
            .lcout(),
            .ltout(n16810_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_LC_1_32_1.C_ON=1'b0;
    defparam i2_4_lut_LC_1_32_1.SEQ_MODE=4'b0000;
    defparam i2_4_lut_LC_1_32_1.LUT_INIT=16'b0101010100010000;
    LogicCell40 i2_4_lut_LC_1_32_1 (
            .in0(N__20147),
            .in1(N__30770),
            .in2(N__17314),
            .in3(N__17308),
            .lcout(n16852),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i11107_2_lut_LC_1_32_2 .C_ON=1'b0;
    defparam \c0.rx.i11107_2_lut_LC_1_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i11107_2_lut_LC_1_32_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i11107_2_lut_LC_1_32_2  (
            .in0(_gnd_net_),
            .in1(N__17938),
            .in2(_gnd_net_),
            .in3(N__18769),
            .lcout(),
            .ltout(\c0.rx.n13452_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_4_lut_adj_398_LC_1_32_3 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_4_lut_adj_398_LC_1_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_4_lut_adj_398_LC_1_32_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.rx.i2_3_lut_4_lut_adj_398_LC_1_32_3  (
            .in0(N__30769),
            .in1(N__30830),
            .in2(N__17311),
            .in3(N__17301),
            .lcout(n16867),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i14784_2_lut_LC_1_32_4 .C_ON=1'b0;
    defparam \c0.rx.i14784_2_lut_LC_1_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i14784_2_lut_LC_1_32_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i14784_2_lut_LC_1_32_4  (
            .in0(_gnd_net_),
            .in1(N__18211),
            .in2(_gnd_net_),
            .in3(N__19680),
            .lcout(n17222),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i2_LC_1_32_5 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i2_LC_1_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i2_LC_1_32_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \c0.rx.r_SM_Main_i2_LC_1_32_5  (
            .in0(N__17940),
            .in1(N__18771),
            .in2(N__19684),
            .in3(N__18217),
            .lcout(r_SM_Main_2_adj_2439),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50482),
            .ce(),
            .sr(N__17293));
    defparam \c0.i3_4_lut_adj_457_LC_2_18_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_457_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_457_LC_2_18_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_457_LC_2_18_0  (
            .in0(N__17390),
            .in1(N__17411),
            .in2(N__17362),
            .in3(N__18140),
            .lcout(\c0.n16772 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i7_LC_2_18_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i7_LC_2_18_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i7_LC_2_18_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i7_LC_2_18_1  (
            .in0(N__17413),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34661),
            .lcout(\c0.FRAME_MATCHER_state_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50381),
            .ce(),
            .sr(N__17401));
    defparam \c0.i1_2_lut_adj_711_LC_2_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_711_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_711_LC_2_18_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_711_LC_2_18_2  (
            .in0(_gnd_net_),
            .in1(N__17412),
            .in2(_gnd_net_),
            .in3(N__32567),
            .lcout(\c0.n16443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_726_LC_2_18_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_726_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_726_LC_2_18_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.i1_2_lut_adj_726_LC_2_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32584),
            .in3(N__17391),
            .lcout(\c0.n16447 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_721_LC_2_18_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_721_LC_2_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_721_LC_2_18_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_721_LC_2_18_4  (
            .in0(N__17361),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32571),
            .lcout(\c0.n16451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_730_LC_2_18_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_730_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_730_LC_2_18_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_730_LC_2_18_5  (
            .in0(N__18141),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29966),
            .lcout(\c0.n16349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_709_LC_2_18_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_709_LC_2_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_709_LC_2_18_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_709_LC_2_18_6  (
            .in0(_gnd_net_),
            .in1(N__21775),
            .in2(_gnd_net_),
            .in3(N__32566),
            .lcout(\c0.n16441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_713_LC_2_18_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_713_LC_2_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_713_LC_2_18_7 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \c0.i1_2_lut_adj_713_LC_2_18_7  (
            .in0(_gnd_net_),
            .in1(N__30109),
            .in2(N__32583),
            .in3(_gnd_net_),
            .lcout(\c0.n16445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i9_LC_2_19_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i9_LC_2_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i9_LC_2_19_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i9_LC_2_19_0  (
            .in0(N__33225),
            .in1(N__33005),
            .in2(_gnd_net_),
            .in3(N__18952),
            .lcout(\c0.FRAME_MATCHER_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50384),
            .ce(),
            .sr(N__20446));
    defparam \c0.FRAME_MATCHER_state_i30_LC_2_20_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i30_LC_2_20_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i30_LC_2_20_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.FRAME_MATCHER_state_i30_LC_2_20_0  (
            .in0(N__34659),
            .in1(N__21710),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_state_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50388),
            .ce(),
            .sr(N__18280));
    defparam \c0.FRAME_MATCHER_i_i31_LC_2_21_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i31_LC_2_21_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i31_LC_2_21_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i31_LC_2_21_0  (
            .in0(N__33256),
            .in1(N__32910),
            .in2(_gnd_net_),
            .in3(N__19492),
            .lcout(\c0.FRAME_MATCHER_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50394),
            .ce(),
            .sr(N__18817));
    defparam \c0.FRAME_MATCHER_i_i3_LC_2_22_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i3_LC_2_22_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i3_LC_2_22_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i3_LC_2_22_0  (
            .in0(N__33260),
            .in1(N__32960),
            .in2(_gnd_net_),
            .in3(N__18841),
            .lcout(\c0.FRAME_MATCHER_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50401),
            .ce(),
            .sr(N__18292));
    defparam \c0.FRAME_MATCHER_i_i14_LC_2_23_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i14_LC_2_23_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i14_LC_2_23_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i14_LC_2_23_0  (
            .in0(N__33265),
            .in1(N__32997),
            .in2(_gnd_net_),
            .in3(N__19057),
            .lcout(\c0.FRAME_MATCHER_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50407),
            .ce(),
            .sr(N__18328));
    defparam \c0.FRAME_MATCHER_i_i19_LC_2_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i19_LC_2_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i19_LC_2_24_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i19_LC_2_24_0  (
            .in0(N__33267),
            .in1(N__32998),
            .in2(_gnd_net_),
            .in3(N__19018),
            .lcout(\c0.FRAME_MATCHER_i_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50414),
            .ce(),
            .sr(N__20386));
    defparam blink_counter_2352__i0_LC_2_25_0.C_ON=1'b1;
    defparam blink_counter_2352__i0_LC_2_25_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i0_LC_2_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i0_LC_2_25_0 (
            .in0(_gnd_net_),
            .in1(N__17467),
            .in2(_gnd_net_),
            .in3(N__17461),
            .lcout(n26),
            .ltout(),
            .carryin(bfn_2_25_0_),
            .carryout(n15590),
            .clk(N__50424),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i1_LC_2_25_1.C_ON=1'b1;
    defparam blink_counter_2352__i1_LC_2_25_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i1_LC_2_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i1_LC_2_25_1 (
            .in0(_gnd_net_),
            .in1(N__17458),
            .in2(_gnd_net_),
            .in3(N__17452),
            .lcout(n25),
            .ltout(),
            .carryin(n15590),
            .carryout(n15591),
            .clk(N__50424),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i2_LC_2_25_2.C_ON=1'b1;
    defparam blink_counter_2352__i2_LC_2_25_2.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i2_LC_2_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i2_LC_2_25_2 (
            .in0(_gnd_net_),
            .in1(N__17449),
            .in2(_gnd_net_),
            .in3(N__17443),
            .lcout(n24),
            .ltout(),
            .carryin(n15591),
            .carryout(n15592),
            .clk(N__50424),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i3_LC_2_25_3.C_ON=1'b1;
    defparam blink_counter_2352__i3_LC_2_25_3.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i3_LC_2_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i3_LC_2_25_3 (
            .in0(_gnd_net_),
            .in1(N__17440),
            .in2(_gnd_net_),
            .in3(N__17434),
            .lcout(n23),
            .ltout(),
            .carryin(n15592),
            .carryout(n15593),
            .clk(N__50424),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i4_LC_2_25_4.C_ON=1'b1;
    defparam blink_counter_2352__i4_LC_2_25_4.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i4_LC_2_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i4_LC_2_25_4 (
            .in0(_gnd_net_),
            .in1(N__17431),
            .in2(_gnd_net_),
            .in3(N__17425),
            .lcout(n22),
            .ltout(),
            .carryin(n15593),
            .carryout(n15594),
            .clk(N__50424),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i5_LC_2_25_5.C_ON=1'b1;
    defparam blink_counter_2352__i5_LC_2_25_5.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i5_LC_2_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i5_LC_2_25_5 (
            .in0(_gnd_net_),
            .in1(N__17422),
            .in2(_gnd_net_),
            .in3(N__17416),
            .lcout(n21),
            .ltout(),
            .carryin(n15594),
            .carryout(n15595),
            .clk(N__50424),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i6_LC_2_25_6.C_ON=1'b1;
    defparam blink_counter_2352__i6_LC_2_25_6.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i6_LC_2_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i6_LC_2_25_6 (
            .in0(_gnd_net_),
            .in1(N__17545),
            .in2(_gnd_net_),
            .in3(N__17539),
            .lcout(n20),
            .ltout(),
            .carryin(n15595),
            .carryout(n15596),
            .clk(N__50424),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i7_LC_2_25_7.C_ON=1'b1;
    defparam blink_counter_2352__i7_LC_2_25_7.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i7_LC_2_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i7_LC_2_25_7 (
            .in0(_gnd_net_),
            .in1(N__17536),
            .in2(_gnd_net_),
            .in3(N__17530),
            .lcout(n19),
            .ltout(),
            .carryin(n15596),
            .carryout(n15597),
            .clk(N__50424),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i8_LC_2_26_0.C_ON=1'b1;
    defparam blink_counter_2352__i8_LC_2_26_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i8_LC_2_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i8_LC_2_26_0 (
            .in0(_gnd_net_),
            .in1(N__17527),
            .in2(_gnd_net_),
            .in3(N__17521),
            .lcout(n18),
            .ltout(),
            .carryin(bfn_2_26_0_),
            .carryout(n15598),
            .clk(N__50432),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i9_LC_2_26_1.C_ON=1'b1;
    defparam blink_counter_2352__i9_LC_2_26_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i9_LC_2_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i9_LC_2_26_1 (
            .in0(_gnd_net_),
            .in1(N__17518),
            .in2(_gnd_net_),
            .in3(N__17512),
            .lcout(n17_adj_2422),
            .ltout(),
            .carryin(n15598),
            .carryout(n15599),
            .clk(N__50432),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i10_LC_2_26_2.C_ON=1'b1;
    defparam blink_counter_2352__i10_LC_2_26_2.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i10_LC_2_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i10_LC_2_26_2 (
            .in0(_gnd_net_),
            .in1(N__17509),
            .in2(_gnd_net_),
            .in3(N__17503),
            .lcout(n16),
            .ltout(),
            .carryin(n15599),
            .carryout(n15600),
            .clk(N__50432),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i11_LC_2_26_3.C_ON=1'b1;
    defparam blink_counter_2352__i11_LC_2_26_3.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i11_LC_2_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i11_LC_2_26_3 (
            .in0(_gnd_net_),
            .in1(N__17500),
            .in2(_gnd_net_),
            .in3(N__17494),
            .lcout(n15),
            .ltout(),
            .carryin(n15600),
            .carryout(n15601),
            .clk(N__50432),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i12_LC_2_26_4.C_ON=1'b1;
    defparam blink_counter_2352__i12_LC_2_26_4.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i12_LC_2_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i12_LC_2_26_4 (
            .in0(_gnd_net_),
            .in1(N__17491),
            .in2(_gnd_net_),
            .in3(N__17485),
            .lcout(n14_adj_2424),
            .ltout(),
            .carryin(n15601),
            .carryout(n15602),
            .clk(N__50432),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i13_LC_2_26_5.C_ON=1'b1;
    defparam blink_counter_2352__i13_LC_2_26_5.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i13_LC_2_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i13_LC_2_26_5 (
            .in0(_gnd_net_),
            .in1(N__17482),
            .in2(_gnd_net_),
            .in3(N__17476),
            .lcout(n13),
            .ltout(),
            .carryin(n15602),
            .carryout(n15603),
            .clk(N__50432),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i14_LC_2_26_6.C_ON=1'b1;
    defparam blink_counter_2352__i14_LC_2_26_6.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i14_LC_2_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i14_LC_2_26_6 (
            .in0(_gnd_net_),
            .in1(N__17473),
            .in2(_gnd_net_),
            .in3(N__17641),
            .lcout(n12_adj_2419),
            .ltout(),
            .carryin(n15603),
            .carryout(n15604),
            .clk(N__50432),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i15_LC_2_26_7.C_ON=1'b1;
    defparam blink_counter_2352__i15_LC_2_26_7.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i15_LC_2_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i15_LC_2_26_7 (
            .in0(_gnd_net_),
            .in1(N__17638),
            .in2(_gnd_net_),
            .in3(N__17632),
            .lcout(n11),
            .ltout(),
            .carryin(n15604),
            .carryout(n15605),
            .clk(N__50432),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i16_LC_2_27_0.C_ON=1'b1;
    defparam blink_counter_2352__i16_LC_2_27_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i16_LC_2_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i16_LC_2_27_0 (
            .in0(_gnd_net_),
            .in1(N__17629),
            .in2(_gnd_net_),
            .in3(N__17623),
            .lcout(n10_adj_2420),
            .ltout(),
            .carryin(bfn_2_27_0_),
            .carryout(n15606),
            .clk(N__50439),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i17_LC_2_27_1.C_ON=1'b1;
    defparam blink_counter_2352__i17_LC_2_27_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i17_LC_2_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i17_LC_2_27_1 (
            .in0(_gnd_net_),
            .in1(N__17620),
            .in2(_gnd_net_),
            .in3(N__17614),
            .lcout(n9),
            .ltout(),
            .carryin(n15606),
            .carryout(n15607),
            .clk(N__50439),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i18_LC_2_27_2.C_ON=1'b1;
    defparam blink_counter_2352__i18_LC_2_27_2.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i18_LC_2_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i18_LC_2_27_2 (
            .in0(_gnd_net_),
            .in1(N__17611),
            .in2(_gnd_net_),
            .in3(N__17605),
            .lcout(n8),
            .ltout(),
            .carryin(n15607),
            .carryout(n15608),
            .clk(N__50439),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i19_LC_2_27_3.C_ON=1'b1;
    defparam blink_counter_2352__i19_LC_2_27_3.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i19_LC_2_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i19_LC_2_27_3 (
            .in0(_gnd_net_),
            .in1(N__17602),
            .in2(_gnd_net_),
            .in3(N__17596),
            .lcout(n7),
            .ltout(),
            .carryin(n15608),
            .carryout(n15609),
            .clk(N__50439),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i20_LC_2_27_4.C_ON=1'b1;
    defparam blink_counter_2352__i20_LC_2_27_4.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i20_LC_2_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i20_LC_2_27_4 (
            .in0(_gnd_net_),
            .in1(N__17593),
            .in2(_gnd_net_),
            .in3(N__17587),
            .lcout(n6_adj_2421),
            .ltout(),
            .carryin(n15609),
            .carryout(n15610),
            .clk(N__50439),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i21_LC_2_27_5.C_ON=1'b1;
    defparam blink_counter_2352__i21_LC_2_27_5.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i21_LC_2_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i21_LC_2_27_5 (
            .in0(_gnd_net_),
            .in1(N__17577),
            .in2(_gnd_net_),
            .in3(N__17566),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n15610),
            .carryout(n15611),
            .clk(N__50439),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i22_LC_2_27_6.C_ON=1'b1;
    defparam blink_counter_2352__i22_LC_2_27_6.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i22_LC_2_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i22_LC_2_27_6 (
            .in0(_gnd_net_),
            .in1(N__17561),
            .in2(_gnd_net_),
            .in3(N__17548),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n15611),
            .carryout(n15612),
            .clk(N__50439),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i23_LC_2_27_7.C_ON=1'b1;
    defparam blink_counter_2352__i23_LC_2_27_7.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i23_LC_2_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i23_LC_2_27_7 (
            .in0(_gnd_net_),
            .in1(N__17744),
            .in2(_gnd_net_),
            .in3(N__17731),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n15612),
            .carryout(n15613),
            .clk(N__50439),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i24_LC_2_28_0.C_ON=1'b1;
    defparam blink_counter_2352__i24_LC_2_28_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i24_LC_2_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i24_LC_2_28_0 (
            .in0(_gnd_net_),
            .in1(N__17723),
            .in2(_gnd_net_),
            .in3(N__17710),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_2_28_0_),
            .carryout(n15614),
            .clk(N__50448),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2352__i25_LC_2_28_1.C_ON=1'b0;
    defparam blink_counter_2352__i25_LC_2_28_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2352__i25_LC_2_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2352__i25_LC_2_28_1 (
            .in0(_gnd_net_),
            .in1(N__17703),
            .in2(_gnd_net_),
            .in3(N__17707),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50448),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_4_lut_LC_2_28_2 .C_ON=1'b0;
    defparam \c0.rx.i2_4_lut_LC_2_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_4_lut_LC_2_28_2 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \c0.rx.i2_4_lut_LC_2_28_2  (
            .in0(N__30759),
            .in1(N__30864),
            .in2(N__33886),
            .in3(N__18413),
            .lcout(\c0.rx.n9323 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i2_LC_2_28_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i2_LC_2_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i2_LC_2_28_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx2.r_Clock_Count__i2_LC_2_28_3  (
            .in0(N__31497),
            .in1(N__17692),
            .in2(_gnd_net_),
            .in3(N__17673),
            .lcout(r_Clock_Count_2_adj_2452),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50448),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i1_LC_2_28_4 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i1_LC_2_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i1_LC_2_28_4 .LUT_INIT=16'b1111000000101000;
    LogicCell40 \c0.tx.r_Bit_Index_i1_LC_2_28_4  (
            .in0(N__24065),
            .in1(N__20812),
            .in2(N__31361),
            .in3(N__19752),
            .lcout(r_Bit_Index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50448),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i5_LC_2_28_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i5_LC_2_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i5_LC_2_28_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i5_LC_2_28_5  (
            .in0(N__31498),
            .in1(N__17872),
            .in2(_gnd_net_),
            .in3(N__17686),
            .lcout(r_Clock_Count_5_adj_2449),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50448),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i1_LC_2_28_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i1_LC_2_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i1_LC_2_28_6 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \c0.tx2.r_Clock_Count__i1_LC_2_28_6  (
            .in0(N__31496),
            .in1(N__17680),
            .in2(N__17854),
            .in3(_gnd_net_),
            .lcout(r_Clock_Count_1_adj_2453),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50448),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i4_4_lut_LC_2_28_7 .C_ON=1'b0;
    defparam \c0.tx2.i4_4_lut_LC_2_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i4_4_lut_LC_2_28_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx2.i4_4_lut_LC_2_28_7  (
            .in0(N__19569),
            .in1(N__17672),
            .in2(N__31408),
            .in3(N__17657),
            .lcout(\c0.tx2.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14702_3_lut_LC_2_29_0.C_ON=1'b0;
    defparam i14702_3_lut_LC_2_29_0.SEQ_MODE=4'b0000;
    defparam i14702_3_lut_LC_2_29_0.LUT_INIT=16'b1000100011111111;
    LogicCell40 i14702_3_lut_LC_2_29_0 (
            .in0(N__31486),
            .in1(N__30997),
            .in2(_gnd_net_),
            .in3(N__17887),
            .lcout(),
            .ltout(n17140_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14847_4_lut_LC_2_29_1.C_ON=1'b0;
    defparam i14847_4_lut_LC_2_29_1.SEQ_MODE=4'b0000;
    defparam i14847_4_lut_LC_2_29_1.LUT_INIT=16'b0000000000101111;
    LogicCell40 i14847_4_lut_LC_2_29_1 (
            .in0(N__17920),
            .in1(N__17761),
            .in2(N__17914),
            .in3(N__17823),
            .lcout(n16817),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_2_lut_4_lut_LC_2_29_2 .C_ON=1'b0;
    defparam \c0.tx2.i1_2_lut_4_lut_LC_2_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_2_lut_4_lut_LC_2_29_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx2.i1_2_lut_4_lut_LC_2_29_2  (
            .in0(N__26390),
            .in1(N__17802),
            .in2(N__29344),
            .in3(N__17778),
            .lcout(n12_adj_2410),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i5_3_lut_LC_2_29_3 .C_ON=1'b0;
    defparam \c0.tx2.i5_3_lut_LC_2_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i5_3_lut_LC_2_29_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx2.i5_3_lut_LC_2_29_3  (
            .in0(N__17870),
            .in1(N__17849),
            .in2(_gnd_net_),
            .in3(N__17833),
            .lcout(n15837),
            .ltout(n15837_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_2_lut_4_lut_adj_399_LC_2_29_4 .C_ON=1'b0;
    defparam \c0.tx2.i1_2_lut_4_lut_adj_399_LC_2_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_2_lut_4_lut_adj_399_LC_2_29_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx2.i1_2_lut_4_lut_adj_399_LC_2_29_4  (
            .in0(N__26392),
            .in1(N__17804),
            .in2(N__17812),
            .in3(N__17780),
            .lcout(r_SM_Main_2_N_2033_1),
            .ltout(r_SM_Main_2_N_2033_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i1_LC_2_29_5 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i1_LC_2_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i1_LC_2_29_5 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \c0.tx2.r_SM_Main_i1_LC_2_29_5  (
            .in0(N__29325),
            .in1(N__31014),
            .in2(N__17809),
            .in3(N__31488),
            .lcout(r_SM_Main_1_adj_2444),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50458),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_2_lut_4_lut_LC_2_29_6 .C_ON=1'b0;
    defparam \c0.tx2.i2_2_lut_4_lut_LC_2_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_2_lut_4_lut_LC_2_29_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx2.i2_2_lut_4_lut_LC_2_29_6  (
            .in0(N__26391),
            .in1(N__17803),
            .in2(N__29343),
            .in3(N__17779),
            .lcout(n9929),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i2_LC_2_29_7 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i2_LC_2_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i2_LC_2_29_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.tx2.r_SM_Main_i2_LC_2_29_7  (
            .in0(N__29326),
            .in1(N__31487),
            .in2(N__31021),
            .in3(N__20004),
            .lcout(r_SM_Main_2_adj_2443),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50458),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i2_LC_2_30_0 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i2_LC_2_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i2_LC_2_30_0 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \c0.rx.r_Clock_Count__i2_LC_2_30_0  (
            .in0(N__18069),
            .in1(N__18049),
            .in2(_gnd_net_),
            .in3(N__20137),
            .lcout(r_Clock_Count_2_adj_2435),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50470),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i3_LC_2_30_1 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i3_LC_2_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i3_LC_2_30_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Clock_Count__i3_LC_2_30_1  (
            .in0(N__23970),
            .in1(N__18034),
            .in2(_gnd_net_),
            .in3(N__17993),
            .lcout(r_Clock_Count_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50470),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i0_LC_2_30_2 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i0_LC_2_30_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i0_LC_2_30_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Clock_Count__i0_LC_2_30_2  (
            .in0(N__23959),
            .in1(N__18028),
            .in2(_gnd_net_),
            .in3(N__17976),
            .lcout(r_Clock_Count_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50470),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i2_LC_2_30_3 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i2_LC_2_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i2_LC_2_30_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.tx.r_Clock_Count__i2_LC_2_30_3  (
            .in0(N__18009),
            .in1(_gnd_net_),
            .in2(N__18022),
            .in3(N__23960),
            .lcout(r_Clock_Count_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50470),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_793_LC_2_30_4.C_ON=1'b0;
    defparam i1_4_lut_adj_793_LC_2_30_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_793_LC_2_30_4.LUT_INIT=16'b1011101010101010;
    LogicCell40 i1_4_lut_adj_793_LC_2_30_4 (
            .in0(N__30848),
            .in1(N__30735),
            .in2(N__33876),
            .in3(N__18115),
            .lcout(n17_adj_2416),
            .ltout(n17_adj_2416_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i4_LC_2_30_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i4_LC_2_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i4_LC_2_30_5 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \c0.rx.r_Clock_Count__i4_LC_2_30_5  (
            .in0(_gnd_net_),
            .in1(N__18630),
            .in2(N__18013),
            .in3(N__18235),
            .lcout(r_Clock_Count_4_adj_2433),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50470),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4_4_lut_LC_2_30_6 .C_ON=1'b0;
    defparam \c0.tx.i4_4_lut_LC_2_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4_4_lut_LC_2_30_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx.i4_4_lut_LC_2_30_6  (
            .in0(N__19722),
            .in1(N__18008),
            .in2(N__17995),
            .in3(N__17975),
            .lcout(),
            .ltout(\c0.tx.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i5_3_lut_LC_2_30_7 .C_ON=1'b0;
    defparam \c0.tx.i5_3_lut_LC_2_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i5_3_lut_LC_2_30_7 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \c0.tx.i5_3_lut_LC_2_30_7  (
            .in0(_gnd_net_),
            .in1(N__17960),
            .in2(N__17944),
            .in3(N__18671),
            .lcout(n15701),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_LC_2_31_1 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_LC_2_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_LC_2_31_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.rx.i1_4_lut_LC_2_31_1  (
            .in0(N__18065),
            .in1(N__20101),
            .in2(N__18717),
            .in3(N__18610),
            .lcout(n16863),
            .ltout(n16863_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_4_lut_LC_2_31_2 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_4_lut_LC_2_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_4_lut_LC_2_31_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.rx.i2_3_lut_4_lut_LC_2_31_2  (
            .in0(N__18747),
            .in1(N__18209),
            .in2(N__17923),
            .in3(N__19672),
            .lcout(\c0.rx.r_SM_Main_2_N_2096_0 ),
            .ltout(\c0.rx.r_SM_Main_2_N_2096_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_2_lut_adj_397_LC_2_31_3 .C_ON=1'b0;
    defparam \c0.rx.i2_2_lut_adj_397_LC_2_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_2_lut_adj_397_LC_2_31_3 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \c0.rx.i2_2_lut_adj_397_LC_2_31_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18118),
            .in3(N__33747),
            .lcout(n6_adj_2461),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i7_LC_2_31_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i7_LC_2_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i7_LC_2_31_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i7_LC_2_31_4  (
            .in0(N__23961),
            .in1(N__19864),
            .in2(_gnd_net_),
            .in3(N__18109),
            .lcout(r_Clock_Count_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50483),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i7_LC_2_31_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i7_LC_2_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i7_LC_2_31_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \c0.rx.r_Clock_Count__i7_LC_2_31_5  (
            .in0(N__18210),
            .in1(N__18148),
            .in2(_gnd_net_),
            .in3(N__20139),
            .lcout(r_Clock_Count_7_adj_2430),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50483),
            .ce(),
            .sr(_gnd_net_));
    defparam i14706_3_lut_LC_2_31_6.C_ON=1'b0;
    defparam i14706_3_lut_LC_2_31_6.SEQ_MODE=4'b0000;
    defparam i14706_3_lut_LC_2_31_6.LUT_INIT=16'b1000100011111111;
    LogicCell40 i14706_3_lut_LC_2_31_6 (
            .in0(N__24066),
            .in1(N__23957),
            .in2(_gnd_net_),
            .in3(N__18499),
            .lcout(),
            .ltout(n17144_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14845_4_lut_LC_2_31_7.C_ON=1'b0;
    defparam i14845_4_lut_LC_2_31_7.SEQ_MODE=4'b0000;
    defparam i14845_4_lut_LC_2_31_7.LUT_INIT=16'b0000010101000101;
    LogicCell40 i14845_4_lut_LC_2_31_7 (
            .in0(N__18471),
            .in1(N__18694),
            .in2(N__18103),
            .in3(N__19774),
            .lcout(n16828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_2_lut_LC_2_32_0 .C_ON=1'b1;
    defparam \c0.rx.add_62_2_lut_LC_2_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_2_lut_LC_2_32_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_2_lut_LC_2_32_0  (
            .in0(N__18175),
            .in1(N__20100),
            .in2(_gnd_net_),
            .in3(N__18076),
            .lcout(n16859),
            .ltout(),
            .carryin(bfn_2_32_0_),
            .carryout(\c0.rx.n15668 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_3_lut_LC_2_32_1 .C_ON=1'b1;
    defparam \c0.rx.add_62_3_lut_LC_2_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_3_lut_LC_2_32_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_3_lut_LC_2_32_1  (
            .in0(N__18179),
            .in1(_gnd_net_),
            .in2(N__18595),
            .in3(N__18073),
            .lcout(n16853),
            .ltout(),
            .carryin(\c0.rx.n15668 ),
            .carryout(\c0.rx.n15669 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_4_lut_LC_2_32_2 .C_ON=1'b1;
    defparam \c0.rx.add_62_4_lut_LC_2_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_4_lut_LC_2_32_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_4_lut_LC_2_32_2  (
            .in0(N__18176),
            .in1(N__18070),
            .in2(_gnd_net_),
            .in3(N__18040),
            .lcout(n16860),
            .ltout(),
            .carryin(\c0.rx.n15669 ),
            .carryout(\c0.rx.n15670 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_5_lut_LC_2_32_3 .C_ON=1'b1;
    defparam \c0.rx.add_62_5_lut_LC_2_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_5_lut_LC_2_32_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_5_lut_LC_2_32_3  (
            .in0(N__18180),
            .in1(N__18713),
            .in2(_gnd_net_),
            .in3(N__18037),
            .lcout(n16858),
            .ltout(),
            .carryin(\c0.rx.n15670 ),
            .carryout(\c0.rx.n15671 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_6_lut_LC_2_32_4 .C_ON=1'b1;
    defparam \c0.rx.add_62_6_lut_LC_2_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_6_lut_LC_2_32_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_6_lut_LC_2_32_4  (
            .in0(N__18177),
            .in1(N__18631),
            .in2(_gnd_net_),
            .in3(N__18226),
            .lcout(n16854),
            .ltout(),
            .carryin(\c0.rx.n15671 ),
            .carryout(\c0.rx.n15672 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_7_lut_LC_2_32_5 .C_ON=1'b1;
    defparam \c0.rx.add_62_7_lut_LC_2_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_7_lut_LC_2_32_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_7_lut_LC_2_32_5  (
            .in0(N__18181),
            .in1(N__18756),
            .in2(_gnd_net_),
            .in3(N__18223),
            .lcout(n16857),
            .ltout(),
            .carryin(\c0.rx.n15672 ),
            .carryout(\c0.rx.n15673 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_8_lut_LC_2_32_6 .C_ON=1'b1;
    defparam \c0.rx.add_62_8_lut_LC_2_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_8_lut_LC_2_32_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_8_lut_LC_2_32_6  (
            .in0(N__18174),
            .in1(N__19678),
            .in2(_gnd_net_),
            .in3(N__18220),
            .lcout(n16856),
            .ltout(),
            .carryin(\c0.rx.n15673 ),
            .carryout(\c0.rx.n15674 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_9_lut_LC_2_32_7 .C_ON=1'b0;
    defparam \c0.rx.add_62_9_lut_LC_2_32_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_9_lut_LC_2_32_7 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \c0.rx.add_62_9_lut_LC_2_32_7  (
            .in0(N__18213),
            .in1(N__18178),
            .in2(_gnd_net_),
            .in3(N__18151),
            .lcout(n16855),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__5__2252_LC_3_17_0 .C_ON=1'b0;
    defparam \c0.data_in_3__5__2252_LC_3_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__5__2252_LC_3_17_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__5__2252_LC_3_17_0  (
            .in0(N__31228),
            .in1(N__27801),
            .in2(_gnd_net_),
            .in3(N__25908),
            .lcout(data_in_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50379),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i15_LC_3_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i15_LC_3_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i15_LC_3_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i15_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(N__18142),
            .in2(_gnd_net_),
            .in3(N__34642),
            .lcout(\c0.FRAME_MATCHER_state_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50385),
            .ce(),
            .sr(N__18127));
    defparam \c0.i10728_2_lut_LC_3_19_0 .C_ON=1'b0;
    defparam \c0.i10728_2_lut_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10728_2_lut_LC_3_19_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i10728_2_lut_LC_3_19_0  (
            .in0(_gnd_net_),
            .in1(N__32260),
            .in2(_gnd_net_),
            .in3(N__23253),
            .lcout(n1651),
            .ltout(n1651_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_776_LC_3_19_1.C_ON=1'b0;
    defparam i1_4_lut_adj_776_LC_3_19_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_776_LC_3_19_1.LUT_INIT=16'b0011001000100010;
    LogicCell40 i1_4_lut_adj_776_LC_3_19_1 (
            .in0(N__21388),
            .in1(N__21676),
            .in2(N__18121),
            .in3(N__22279),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10657_3_lut_4_lut_LC_3_19_2 .C_ON=1'b0;
    defparam \c0.i10657_3_lut_4_lut_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10657_3_lut_4_lut_LC_3_19_2 .LUT_INIT=16'b1110101011111010;
    LogicCell40 \c0.i10657_3_lut_4_lut_LC_3_19_2  (
            .in0(N__21583),
            .in1(N__32261),
            .in2(N__22287),
            .in3(N__23254),
            .lcout(FRAME_MATCHER_state_31_N_1440_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_775_LC_3_19_3.C_ON=1'b0;
    defparam i1_4_lut_adj_775_LC_3_19_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_775_LC_3_19_3.LUT_INIT=16'b1101110001010000;
    LogicCell40 i1_4_lut_adj_775_LC_3_19_3 (
            .in0(N__27907),
            .in1(N__28036),
            .in2(N__22309),
            .in3(N__22280),
            .lcout(),
            .ltout(n6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_3_19_4.C_ON=1'b0;
    defparam i3_4_lut_LC_3_19_4.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_3_19_4.LUT_INIT=16'b1111111111010101;
    LogicCell40 i3_4_lut_LC_3_19_4 (
            .in0(N__32454),
            .in1(N__18268),
            .in2(N__18262),
            .in3(N__18259),
            .lcout(),
            .ltout(n8_adj_2459_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i1_LC_3_19_5 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i1_LC_3_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_state_i1_LC_3_19_5 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \c0.FRAME_MATCHER_state_i1_LC_3_19_5  (
            .in0(N__33278),
            .in1(N__18244),
            .in2(N__18253),
            .in3(N__18250),
            .lcout(FRAME_MATCHER_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50389),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_798_LC_3_19_6.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_798_LC_3_19_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_798_LC_3_19_6.LUT_INIT=16'b0010000000110000;
    LogicCell40 i1_3_lut_4_lut_adj_798_LC_3_19_6 (
            .in0(N__32268),
            .in1(N__22354),
            .in2(N__22288),
            .in3(N__23255),
            .lcout(n3_adj_2408),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_725_LC_3_19_7 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_725_LC_3_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_725_LC_3_19_7 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \c0.i1_4_lut_adj_725_LC_3_19_7  (
            .in0(N__18787),
            .in1(N__32892),
            .in2(N__22702),
            .in3(N__22324),
            .lcout(\c0.n4_adj_2360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i27_LC_3_20_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i27_LC_3_20_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i27_LC_3_20_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i27_LC_3_20_0  (
            .in0(_gnd_net_),
            .in1(N__25328),
            .in2(_gnd_net_),
            .in3(N__34643),
            .lcout(\c0.FRAME_MATCHER_state_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50395),
            .ce(),
            .sr(N__25309));
    defparam \c0.i10765_2_lut_3_lut_4_lut_LC_3_21_0 .C_ON=1'b0;
    defparam \c0.i10765_2_lut_3_lut_4_lut_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10765_2_lut_3_lut_4_lut_LC_3_21_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10765_2_lut_3_lut_4_lut_LC_3_21_0  (
            .in0(N__23428),
            .in1(N__23258),
            .in2(N__24440),
            .in3(N__23049),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_5 ),
            .ltout(\c0.FRAME_MATCHER_i_31_N_1312_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_5_i3_2_lut_LC_3_21_1 .C_ON=1'b0;
    defparam \c0.select_238_Select_5_i3_2_lut_LC_3_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_5_i3_2_lut_LC_3_21_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \c0.select_238_Select_5_i3_2_lut_LC_3_21_1  (
            .in0(N__29728),
            .in1(_gnd_net_),
            .in2(N__18238),
            .in3(_gnd_net_),
            .lcout(\c0.n3_adj_2256 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i5_LC_3_21_2 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i5_LC_3_21_2 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i5_LC_3_21_2 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i5_LC_3_21_2  (
            .in0(N__33255),
            .in1(N__32896),
            .in2(_gnd_net_),
            .in3(N__18988),
            .lcout(\c0.FRAME_MATCHER_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50402),
            .ce(),
            .sr(N__18310));
    defparam \c0.i10766_2_lut_3_lut_4_lut_LC_3_21_3 .C_ON=1'b0;
    defparam \c0.i10766_2_lut_3_lut_4_lut_LC_3_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10766_2_lut_3_lut_4_lut_LC_3_21_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10766_2_lut_3_lut_4_lut_LC_3_21_3  (
            .in0(N__23259),
            .in1(N__24491),
            .in2(N__23064),
            .in3(N__23426),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_4 ),
            .ltout(\c0.FRAME_MATCHER_i_31_N_1312_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_4_i3_2_lut_LC_3_21_4 .C_ON=1'b0;
    defparam \c0.select_238_Select_4_i3_2_lut_LC_3_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_4_i3_2_lut_LC_3_21_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.select_238_Select_4_i3_2_lut_LC_3_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18298),
            .in3(N__29727),
            .lcout(\c0.n3_adj_2257 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10767_2_lut_3_lut_4_lut_LC_3_21_5 .C_ON=1'b0;
    defparam \c0.i10767_2_lut_3_lut_4_lut_LC_3_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10767_2_lut_3_lut_4_lut_LC_3_21_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10767_2_lut_3_lut_4_lut_LC_3_21_5  (
            .in0(N__23260),
            .in1(N__25120),
            .in2(N__23065),
            .in3(N__23427),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_3 ),
            .ltout(\c0.FRAME_MATCHER_i_31_N_1312_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_3_i3_2_lut_LC_3_21_6 .C_ON=1'b0;
    defparam \c0.select_238_Select_3_i3_2_lut_LC_3_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_3_i3_2_lut_LC_3_21_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.select_238_Select_3_i3_2_lut_LC_3_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18295),
            .in3(N__29726),
            .lcout(\c0.n3_adj_2258 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_42_i10_2_lut_3_lut_LC_3_21_7 .C_ON=1'b0;
    defparam \c0.equal_42_i10_2_lut_3_lut_LC_3_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.equal_42_i10_2_lut_3_lut_LC_3_21_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.equal_42_i10_2_lut_3_lut_LC_3_21_7  (
            .in0(N__25116),
            .in1(N__24490),
            .in2(_gnd_net_),
            .in3(N__24429),
            .lcout(\c0.n10_adj_2329 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i13_LC_3_22_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i13_LC_3_22_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i13_LC_3_22_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i13_LC_3_22_0  (
            .in0(N__32912),
            .in1(N__33258),
            .in2(_gnd_net_),
            .in3(N__19075),
            .lcout(\c0.FRAME_MATCHER_i_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50408),
            .ce(),
            .sr(N__18322));
    defparam \c0.i1_2_lut_adj_762_LC_3_22_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_762_LC_3_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_762_LC_3_22_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_762_LC_3_22_1  (
            .in0(_gnd_net_),
            .in1(N__21712),
            .in2(_gnd_net_),
            .in3(N__29941),
            .lcout(\c0.n16379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_LC_3_22_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_LC_3_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_LC_3_22_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i2_2_lut_LC_3_22_2  (
            .in0(_gnd_net_),
            .in1(N__30027),
            .in2(_gnd_net_),
            .in3(N__30117),
            .lcout(\c0.n33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i10739_2_lut_LC_3_22_3 .C_ON=1'b0;
    defparam \c0.rx.i10739_2_lut_LC_3_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i10739_2_lut_LC_3_22_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.rx.i10739_2_lut_LC_3_22_3  (
            .in0(N__19927),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19975),
            .lcout(n13082),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_400_LC_3_22_5 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_400_LC_3_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_400_LC_3_22_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.i1_2_lut_adj_400_LC_3_22_5  (
            .in0(_gnd_net_),
            .in1(N__31728),
            .in2(_gnd_net_),
            .in3(N__31672),
            .lcout(n445),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10755_2_lut_3_lut_4_lut_LC_3_23_0 .C_ON=1'b0;
    defparam \c0.i10755_2_lut_3_lut_4_lut_LC_3_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10755_2_lut_3_lut_4_lut_LC_3_23_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10755_2_lut_3_lut_4_lut_LC_3_23_0  (
            .in0(N__23417),
            .in1(N__22996),
            .in2(N__28249),
            .in3(N__23236),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i15_LC_3_23_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i15_LC_3_23_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i15_LC_3_23_1 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i15_LC_3_23_1  (
            .in0(N__32913),
            .in1(N__33259),
            .in2(_gnd_net_),
            .in3(N__19036),
            .lcout(\c0.FRAME_MATCHER_i_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50415),
            .ce(),
            .sr(N__18337));
    defparam \c0.select_238_Select_15_i3_2_lut_3_lut_4_lut_LC_3_23_2 .C_ON=1'b0;
    defparam \c0.select_238_Select_15_i3_2_lut_3_lut_4_lut_LC_3_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_15_i3_2_lut_3_lut_4_lut_LC_3_23_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_15_i3_2_lut_3_lut_4_lut_LC_3_23_2  (
            .in0(N__29735),
            .in1(N__23008),
            .in2(N__28250),
            .in3(N__22704),
            .lcout(\c0.n3_adj_2242 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10756_2_lut_3_lut_4_lut_LC_3_23_3 .C_ON=1'b0;
    defparam \c0.i10756_2_lut_3_lut_4_lut_LC_3_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10756_2_lut_3_lut_4_lut_LC_3_23_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10756_2_lut_3_lut_4_lut_LC_3_23_3  (
            .in0(N__23237),
            .in1(N__28283),
            .in2(N__23046),
            .in3(N__23415),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_14_i3_2_lut_3_lut_4_lut_LC_3_23_4 .C_ON=1'b0;
    defparam \c0.select_238_Select_14_i3_2_lut_3_lut_4_lut_LC_3_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_14_i3_2_lut_3_lut_4_lut_LC_3_23_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_14_i3_2_lut_3_lut_4_lut_LC_3_23_4  (
            .in0(N__29734),
            .in1(N__23007),
            .in2(N__28290),
            .in3(N__22705),
            .lcout(\c0.n3_adj_2243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10757_2_lut_3_lut_4_lut_LC_3_23_5 .C_ON=1'b0;
    defparam \c0.i10757_2_lut_3_lut_4_lut_LC_3_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10757_2_lut_3_lut_4_lut_LC_3_23_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10757_2_lut_3_lut_4_lut_LC_3_23_5  (
            .in0(N__23238),
            .in1(N__24337),
            .in2(N__23047),
            .in3(N__23418),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_13_i3_2_lut_3_lut_4_lut_LC_3_23_6 .C_ON=1'b0;
    defparam \c0.select_238_Select_13_i3_2_lut_3_lut_4_lut_LC_3_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_13_i3_2_lut_3_lut_4_lut_LC_3_23_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_13_i3_2_lut_3_lut_4_lut_LC_3_23_6  (
            .in0(N__29733),
            .in1(N__23006),
            .in2(N__24347),
            .in3(N__22703),
            .lcout(\c0.n3_adj_2244 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10758_2_lut_3_lut_4_lut_LC_3_23_7 .C_ON=1'b0;
    defparam \c0.i10758_2_lut_3_lut_4_lut_LC_3_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10758_2_lut_3_lut_4_lut_LC_3_23_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10758_2_lut_3_lut_4_lut_LC_3_23_7  (
            .in0(N__23239),
            .in1(N__25470),
            .in2(N__23048),
            .in3(N__23416),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i25_LC_3_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i25_LC_3_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i25_LC_3_24_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i25_LC_3_24_0  (
            .in0(N__32914),
            .in1(N__33261),
            .in2(_gnd_net_),
            .in3(N__19150),
            .lcout(\c0.FRAME_MATCHER_i_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50425),
            .ce(),
            .sr(N__20290));
    defparam \c0.data_in_1__0__2273_LC_3_25_1 .C_ON=1'b0;
    defparam \c0.data_in_1__0__2273_LC_3_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__0__2273_LC_3_25_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_1__0__2273_LC_3_25_1  (
            .in0(N__27744),
            .in1(N__23572),
            .in2(_gnd_net_),
            .in3(N__20052),
            .lcout(data_in_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50433),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_54_i4_2_lut_LC_3_25_2 .C_ON=1'b0;
    defparam \c0.rx.equal_54_i4_2_lut_LC_3_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_54_i4_2_lut_LC_3_25_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.rx.equal_54_i4_2_lut_LC_3_25_2  (
            .in0(N__19918),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19971),
            .lcout(n4_adj_2460),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i7_LC_3_25_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i7_LC_3_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i7_LC_3_25_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i7_LC_3_25_3  (
            .in0(N__20718),
            .in1(N__33764),
            .in2(N__26490),
            .in3(N__20508),
            .lcout(rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50433),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__0__2265_LC_3_25_4 .C_ON=1'b0;
    defparam \c0.data_in_2__0__2265_LC_3_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__0__2265_LC_3_25_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_2__0__2265_LC_3_25_4  (
            .in0(N__23573),
            .in1(N__22110),
            .in2(_gnd_net_),
            .in3(N__27746),
            .lcout(data_in_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50433),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i5_LC_3_25_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i5_LC_3_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i5_LC_3_25_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i5_LC_3_25_5  (
            .in0(N__20539),
            .in1(N__33763),
            .in2(N__31202),
            .in3(N__20507),
            .lcout(rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50433),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__1__2272_LC_3_25_6 .C_ON=1'b0;
    defparam \c0.data_in_1__1__2272_LC_3_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__1__2272_LC_3_25_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_1__1__2272_LC_3_25_6  (
            .in0(N__19252),
            .in1(N__22408),
            .in2(_gnd_net_),
            .in3(N__27745),
            .lcout(data_in_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50433),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__5__2276_LC_3_25_7 .C_ON=1'b0;
    defparam \c0.data_in_0__5__2276_LC_3_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__5__2276_LC_3_25_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0__5__2276_LC_3_25_7  (
            .in0(N__27743),
            .in1(N__22077),
            .in2(_gnd_net_),
            .in3(N__18367),
            .lcout(data_in_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50433),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__3__2270_LC_3_26_0 .C_ON=1'b0;
    defparam \c0.data_in_1__3__2270_LC_3_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__3__2270_LC_3_26_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_1__3__2270_LC_3_26_0  (
            .in0(N__20595),
            .in1(N__27708),
            .in2(_gnd_net_),
            .in3(N__19542),
            .lcout(data_in_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50440),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14734_2_lut_LC_3_26_1 .C_ON=1'b0;
    defparam \c0.i14734_2_lut_LC_3_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14734_2_lut_LC_3_26_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i14734_2_lut_LC_3_26_1  (
            .in0(_gnd_net_),
            .in1(N__20048),
            .in2(_gnd_net_),
            .in3(N__20594),
            .lcout(),
            .ltout(\c0.n17172_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14824_4_lut_LC_3_26_2 .C_ON=1'b0;
    defparam \c0.i14824_4_lut_LC_3_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14824_4_lut_LC_3_26_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i14824_4_lut_LC_3_26_2  (
            .in0(N__18348),
            .in1(N__18365),
            .in2(N__18340),
            .in3(N__18378),
            .lcout(\c0.n17262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_567_LC_3_26_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_567_LC_3_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_567_LC_3_26_3 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.i2_3_lut_adj_567_LC_3_26_3  (
            .in0(N__25084),
            .in1(N__21653),
            .in2(_gnd_net_),
            .in3(N__32705),
            .lcout(\c0.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__7__2274_LC_3_26_4 .C_ON=1'b0;
    defparam \c0.data_in_0__7__2274_LC_3_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__7__2274_LC_3_26_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0__7__2274_LC_3_26_4  (
            .in0(N__18379),
            .in1(N__23539),
            .in2(_gnd_net_),
            .in3(N__27709),
            .lcout(data_in_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50440),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14826_3_lut_LC_3_26_5 .C_ON=1'b0;
    defparam \c0.i14826_3_lut_LC_3_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i14826_3_lut_LC_3_26_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i14826_3_lut_LC_3_26_5  (
            .in0(N__19541),
            .in1(N__19476),
            .in2(_gnd_net_),
            .in3(N__19599),
            .lcout(\c0.n17264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__5__2268_LC_3_26_6 .C_ON=1'b0;
    defparam \c0.data_in_1__5__2268_LC_3_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__5__2268_LC_3_26_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_1__5__2268_LC_3_26_6  (
            .in0(N__18366),
            .in1(N__25894),
            .in2(_gnd_net_),
            .in3(N__27710),
            .lcout(data_in_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50440),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__4__2277_LC_3_26_7 .C_ON=1'b0;
    defparam \c0.data_in_0__4__2277_LC_3_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__4__2277_LC_3_26_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0__4__2277_LC_3_26_7  (
            .in0(N__27707),
            .in1(N__19600),
            .in2(_gnd_net_),
            .in3(N__18349),
            .lcout(data_in_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50440),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i75_LC_3_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i75_LC_3_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i75_LC_3_27_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i75_LC_3_27_0  (
            .in0(N__26936),
            .in1(N__28803),
            .in2(N__22563),
            .in3(N__31135),
            .lcout(\c0.data_in_frame_9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50449),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__1__2256_LC_3_27_1 .C_ON=1'b0;
    defparam \c0.data_in_3__1__2256_LC_3_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__1__2256_LC_3_27_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_in_3__1__2256_LC_3_27_1  (
            .in0(N__27705),
            .in1(_gnd_net_),
            .in2(N__30665),
            .in3(N__19272),
            .lcout(data_in_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50449),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i4216_2_lut_LC_3_27_2 .C_ON=1'b0;
    defparam \c0.tx2.i4216_2_lut_LC_3_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i4216_2_lut_LC_3_27_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.tx2.i4216_2_lut_LC_3_27_2  (
            .in0(_gnd_net_),
            .in1(N__27248),
            .in2(_gnd_net_),
            .in3(N__29342),
            .lcout(\c0.tx2.n6480 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__6__2275_LC_3_27_3 .C_ON=1'b0;
    defparam \c0.data_in_0__6__2275_LC_3_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__6__2275_LC_3_27_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0__6__2275_LC_3_27_3  (
            .in0(N__27704),
            .in1(N__19477),
            .in2(_gnd_net_),
            .in3(N__27610),
            .lcout(data_in_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50449),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_LC_3_27_4 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_LC_3_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_LC_3_27_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.rx.i1_2_lut_LC_3_27_4  (
            .in0(_gnd_net_),
            .in1(N__20697),
            .in2(_gnd_net_),
            .in3(N__20658),
            .lcout(n9472),
            .ltout(n9472_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i1_LC_3_27_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i1_LC_3_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i1_LC_3_27_5 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.rx.r_Rx_Byte_i1_LC_3_27_5  (
            .in0(N__30649),
            .in1(N__20625),
            .in2(N__18427),
            .in3(N__33753),
            .lcout(rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50449),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i13_4_lut_4_lut_LC_3_27_6 .C_ON=1'b0;
    defparam \c0.rx.i13_4_lut_4_lut_LC_3_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i13_4_lut_4_lut_LC_3_27_6 .LUT_INIT=16'b0010010100000101;
    LogicCell40 \c0.rx.i13_4_lut_4_lut_LC_3_27_6  (
            .in0(N__30760),
            .in1(N__30875),
            .in2(N__33859),
            .in3(N__18420),
            .lcout(),
            .ltout(\c0.rx.n10086_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_52_LC_3_27_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_52_LC_3_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_DV_52_LC_3_27_7 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \c0.rx.r_Rx_DV_52_LC_3_27_7  (
            .in0(N__27706),
            .in1(N__30761),
            .in2(N__18424),
            .in3(N__30876),
            .lcout(rx_data_ready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50449),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i57_LC_3_28_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i57_LC_3_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i57_LC_3_28_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i57_LC_3_28_1  (
            .in0(N__25585),
            .in1(N__25770),
            .in2(_gnd_net_),
            .in3(N__20845),
            .lcout(data_in_frame_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50459),
            .ce(),
            .sr(_gnd_net_));
    defparam i14959_3_lut_LC_3_28_2.C_ON=1'b0;
    defparam i14959_3_lut_LC_3_28_2.SEQ_MODE=4'b0000;
    defparam i14959_3_lut_LC_3_28_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 i14959_3_lut_LC_3_28_2 (
            .in0(N__31343),
            .in1(N__35443),
            .in2(_gnd_net_),
            .in3(N__29368),
            .lcout(n17397),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i10646_2_lut_LC_3_28_4 .C_ON=1'b0;
    defparam \c0.tx2.i10646_2_lut_LC_3_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i10646_2_lut_LC_3_28_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx2.i10646_2_lut_LC_3_28_4  (
            .in0(_gnd_net_),
            .in1(N__29320),
            .in2(_gnd_net_),
            .in3(N__20001),
            .lcout(\c0.tx2.n1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_56_i4_2_lut_LC_3_28_5 .C_ON=1'b0;
    defparam \c0.rx.equal_56_i4_2_lut_LC_3_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_56_i4_2_lut_LC_3_28_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.equal_56_i4_2_lut_LC_3_28_5  (
            .in0(_gnd_net_),
            .in1(N__19961),
            .in2(_gnd_net_),
            .in3(N__19917),
            .lcout(n4_adj_2409),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_3_28_6 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_3_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_3_28_6 .LUT_INIT=16'b1101111100110011;
    LogicCell40 \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_3_28_6  (
            .in0(N__18574),
            .in1(N__33858),
            .in2(N__19970),
            .in3(N__18421),
            .lcout(n13440),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_4_lut_LC_3_29_0 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_4_lut_LC_3_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_4_lut_LC_3_29_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx.i1_2_lut_4_lut_LC_3_29_0  (
            .in0(N__19804),
            .in1(N__19825),
            .in2(N__19872),
            .in3(N__18470),
            .lcout(n14060),
            .ltout(n14060_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i14754_4_lut_LC_3_29_1 .C_ON=1'b0;
    defparam \c0.tx.i14754_4_lut_LC_3_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i14754_4_lut_LC_3_29_1 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \c0.tx.i14754_4_lut_LC_3_29_1  (
            .in0(N__24156),
            .in1(N__24043),
            .in2(N__18382),
            .in3(N__23892),
            .lcout(\c0.tx.n14082 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i0_LC_3_29_2 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i0_LC_3_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i0_LC_3_29_2 .LUT_INIT=16'b0000010000001110;
    LogicCell40 \c0.tx.r_SM_Main_i0_LC_3_29_2  (
            .in0(N__24169),
            .in1(N__19630),
            .in2(N__23933),
            .in3(N__24103),
            .lcout(r_SM_Main_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50471),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i5592_4_lut_LC_3_29_3 .C_ON=1'b0;
    defparam \c0.tx2.i5592_4_lut_LC_3_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i5592_4_lut_LC_3_29_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \c0.tx2.i5592_4_lut_LC_3_29_3  (
            .in0(N__31013),
            .in1(N__27249),
            .in2(N__29239),
            .in3(N__20002),
            .lcout(),
            .ltout(n7866_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i0_LC_3_29_4 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i0_LC_3_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i0_LC_3_29_4 .LUT_INIT=16'b0001000100110000;
    LogicCell40 \c0.tx2.r_SM_Main_i0_LC_3_29_4  (
            .in0(N__20003),
            .in1(N__31499),
            .in2(N__18505),
            .in3(N__29327),
            .lcout(r_SM_Main_0_adj_2445),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50471),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i14832_3_lut_4_lut_LC_3_29_5 .C_ON=1'b0;
    defparam \c0.rx.i14832_3_lut_4_lut_LC_3_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i14832_3_lut_4_lut_LC_3_29_5 .LUT_INIT=16'b1111111101001100;
    LogicCell40 \c0.rx.i14832_3_lut_4_lut_LC_3_29_5  (
            .in0(N__18572),
            .in1(N__30749),
            .in2(N__19969),
            .in3(N__18550),
            .lcout(n10425),
            .ltout(n10425_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i2_LC_3_29_6 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i2_LC_3_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i2_LC_3_29_6 .LUT_INIT=16'b1001000011000000;
    LogicCell40 \c0.rx.r_Bit_Index_i2_LC_3_29_6  (
            .in0(N__18551),
            .in1(N__19957),
            .in2(N__18502),
            .in3(N__18573),
            .lcout(r_Bit_Index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50471),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_4_lut_adj_402_LC_3_29_7 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_4_lut_adj_402_LC_3_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_4_lut_adj_402_LC_3_29_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx.i1_2_lut_4_lut_adj_402_LC_3_29_7  (
            .in0(N__19824),
            .in1(N__19865),
            .in2(N__24171),
            .in3(N__19803),
            .lcout(n12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i10933_2_lut_LC_3_30_0 .C_ON=1'b0;
    defparam \c0.tx.i10933_2_lut_LC_3_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i10933_2_lut_LC_3_30_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.i10933_2_lut_LC_3_30_0  (
            .in0(_gnd_net_),
            .in1(N__24039),
            .in2(_gnd_net_),
            .in3(N__23953),
            .lcout(n13276),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_LC_3_30_1.C_ON=1'b0;
    defparam i1_3_lut_4_lut_LC_3_30_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_LC_3_30_1.LUT_INIT=16'b0101000000010000;
    LogicCell40 i1_3_lut_4_lut_LC_3_30_1 (
            .in0(N__23954),
            .in1(N__19767),
            .in2(N__24064),
            .in3(N__18497),
            .lcout(),
            .ltout(n10_adj_2415_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_789_LC_3_30_2.C_ON=1'b0;
    defparam i1_4_lut_adj_789_LC_3_30_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_789_LC_3_30_2.LUT_INIT=16'b0000000011110010;
    LogicCell40 i1_4_lut_adj_789_LC_3_30_2 (
            .in0(N__18498),
            .in1(N__18481),
            .in2(N__18475),
            .in3(N__18472),
            .lcout(n16844),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i0_LC_3_30_3 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i0_LC_3_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i0_LC_3_30_3 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \c0.rx.r_Bit_Index_i0_LC_3_30_3  (
            .in0(N__20693),
            .in1(N__18552),
            .in2(_gnd_net_),
            .in3(N__18520),
            .lcout(r_Bit_Index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50484),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i1_LC_3_30_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i1_LC_3_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i1_LC_3_30_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i1_LC_3_30_4  (
            .in0(N__23958),
            .in1(N__18675),
            .in2(_gnd_net_),
            .in3(N__18685),
            .lcout(r_Clock_Count_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50484),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i1_LC_3_30_5 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i1_LC_3_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i1_LC_3_30_5 .LUT_INIT=16'b0000000101010001;
    LogicCell40 \c0.rx.r_SM_Main_i1_LC_3_30_5  (
            .in0(N__30874),
            .in1(N__18655),
            .in2(N__30768),
            .in3(N__18643),
            .lcout(r_SM_Main_1_adj_2440),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50484),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_2_lut_LC_3_30_6 .C_ON=1'b0;
    defparam \c0.rx.i2_2_lut_LC_3_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_2_lut_LC_3_30_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i2_2_lut_LC_3_30_6  (
            .in0(_gnd_net_),
            .in1(N__18626),
            .in2(_gnd_net_),
            .in3(N__18587),
            .lcout(\c0.rx.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i1_LC_3_30_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i1_LC_3_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i1_LC_3_30_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \c0.rx.r_Clock_Count__i1_LC_3_30_7  (
            .in0(N__18588),
            .in1(N__18604),
            .in2(_gnd_net_),
            .in3(N__20138),
            .lcout(r_Clock_Count_1_adj_2436),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50484),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_2_lut_3_lut_4_lut_LC_3_31_0 .C_ON=1'b0;
    defparam \c0.tx.i2_2_lut_3_lut_4_lut_LC_3_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_2_lut_3_lut_4_lut_LC_3_31_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.tx.i2_2_lut_3_lut_4_lut_LC_3_31_0  (
            .in0(N__31706),
            .in1(N__23956),
            .in2(N__24049),
            .in3(N__24172),
            .lcout(n8730),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14840_4_lut_LC_3_31_1 .C_ON=1'b0;
    defparam \c0.i14840_4_lut_LC_3_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14840_4_lut_LC_3_31_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14840_4_lut_LC_3_31_1  (
            .in0(N__21235),
            .in1(N__20929),
            .in2(N__20185),
            .in3(N__20026),
            .lcout(\c0.n17278 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_395_LC_3_31_2 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_395_LC_3_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_395_LC_3_31_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i1_2_lut_adj_395_LC_3_31_2  (
            .in0(_gnd_net_),
            .in1(N__19913),
            .in2(_gnd_net_),
            .in3(N__20685),
            .lcout(n4_adj_2411),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i1_LC_3_31_3 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i1_LC_3_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i1_LC_3_31_3 .LUT_INIT=16'b1101001000000000;
    LogicCell40 \c0.rx.r_Bit_Index_i1_LC_3_31_3  (
            .in0(N__20686),
            .in1(N__18553),
            .in2(N__19925),
            .in3(N__18519),
            .lcout(r_Bit_Index_1_adj_2438),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50494),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i5_LC_3_31_4 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i5_LC_3_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i5_LC_3_31_4 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i5_LC_3_31_4  (
            .in0(N__20141),
            .in1(N__18757),
            .in2(_gnd_net_),
            .in3(N__18778),
            .lcout(r_Clock_Count_5_adj_2432),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50494),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i3_LC_3_31_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i3_LC_3_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i3_LC_3_31_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \c0.rx.r_Clock_Count__i3_LC_3_31_5  (
            .in0(N__18718),
            .in1(N__18724),
            .in2(_gnd_net_),
            .in3(N__20140),
            .lcout(r_Clock_Count_3_adj_2434),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50494),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_3_lut_4_lut_LC_3_31_6 .C_ON=1'b0;
    defparam \c0.tx.i1_3_lut_4_lut_LC_3_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_3_lut_4_lut_LC_3_31_6 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.tx.i1_3_lut_4_lut_LC_3_31_6  (
            .in0(N__27532),
            .in1(N__24250),
            .in2(N__31721),
            .in3(N__31670),
            .lcout(n16886),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_401_LC_3_31_7 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_401_LC_3_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_401_LC_3_31_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.tx.i1_2_lut_adj_401_LC_3_31_7  (
            .in0(N__23955),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24023),
            .lcout(n9406),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_transmit_2156_LC_3_32_6 .C_ON=1'b0;
    defparam \c0.tx_transmit_2156_LC_3_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx_transmit_2156_LC_3_32_6 .LUT_INIT=16'b0000011100000010;
    LogicCell40 \c0.tx_transmit_2156_LC_3_32_6  (
            .in0(N__42607),
            .in1(N__27064),
            .in2(N__31612),
            .in3(N__27280),
            .lcout(\c0.r_SM_Main_2_N_2036_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50506),
            .ce(),
            .sr(N__45550));
    defparam \c0.FRAME_MATCHER_i_i24_LC_4_15_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i24_LC_4_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i24_LC_4_15_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i24_LC_4_15_0  (
            .in0(N__33185),
            .in1(N__33007),
            .in2(_gnd_net_),
            .in3(N__19162),
            .lcout(\c0.FRAME_MATCHER_i_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50396),
            .ce(),
            .sr(N__20317));
    defparam \c0.FRAME_MATCHER_i_i21_LC_4_16_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i21_LC_4_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i21_LC_4_16_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i21_LC_4_16_0  (
            .in0(N__33161),
            .in1(N__33006),
            .in2(_gnd_net_),
            .in3(N__19213),
            .lcout(\c0.FRAME_MATCHER_i_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50390),
            .ce(),
            .sr(N__20233));
    defparam \c0.FRAME_MATCHER_i_i28_LC_4_17_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i28_LC_4_17_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i28_LC_4_17_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i28_LC_4_17_0  (
            .in0(N__33098),
            .in1(N__32989),
            .in2(_gnd_net_),
            .in3(N__19111),
            .lcout(\c0.FRAME_MATCHER_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50382),
            .ce(),
            .sr(N__20227));
    defparam \c0.FRAME_MATCHER_i_i30_LC_4_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i30_LC_4_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i30_LC_4_18_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i30_LC_4_18_0  (
            .in0(N__33184),
            .in1(N__32947),
            .in2(_gnd_net_),
            .in3(N__19510),
            .lcout(\c0.FRAME_MATCHER_i_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50391),
            .ce(),
            .sr(N__18823));
    defparam \c0.FRAME_MATCHER_i_i29_LC_4_19_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i29_LC_4_19_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i29_LC_4_19_1 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i29_LC_4_19_1  (
            .in0(N__33186),
            .in1(N__32893),
            .in2(_gnd_net_),
            .in3(N__19522),
            .lcout(\c0.FRAME_MATCHER_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50397),
            .ce(),
            .sr(N__18832));
    defparam \c0.select_238_Select_29_i3_2_lut_3_lut_4_lut_LC_4_19_2 .C_ON=1'b0;
    defparam \c0.select_238_Select_29_i3_2_lut_3_lut_4_lut_LC_4_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_29_i3_2_lut_3_lut_4_lut_LC_4_19_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_29_i3_2_lut_3_lut_4_lut_LC_4_19_2  (
            .in0(N__23036),
            .in1(N__29679),
            .in2(N__22163),
            .in3(N__22674),
            .lcout(\c0.n3_adj_2217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_30_i3_2_lut_3_lut_4_lut_LC_4_19_4 .C_ON=1'b0;
    defparam \c0.select_238_Select_30_i3_2_lut_3_lut_4_lut_LC_4_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_30_i3_2_lut_3_lut_4_lut_LC_4_19_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_30_i3_2_lut_3_lut_4_lut_LC_4_19_4  (
            .in0(N__23037),
            .in1(N__29680),
            .in2(N__24908),
            .in3(N__22675),
            .lcout(\c0.n3_adj_2215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_31_i3_2_lut_3_lut_4_lut_LC_4_19_5 .C_ON=1'b0;
    defparam \c0.select_238_Select_31_i3_2_lut_3_lut_4_lut_LC_4_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_31_i3_2_lut_3_lut_4_lut_LC_4_19_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_31_i3_2_lut_3_lut_4_lut_LC_4_19_5  (
            .in0(N__22672),
            .in1(N__22494),
            .in2(N__29711),
            .in3(N__23038),
            .lcout(\c0.n3_adj_2210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_8_i3_2_lut_3_lut_4_lut_LC_4_19_6 .C_ON=1'b0;
    defparam \c0.select_238_Select_8_i3_2_lut_3_lut_4_lut_LC_4_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_8_i3_2_lut_3_lut_4_lut_LC_4_19_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_8_i3_2_lut_3_lut_4_lut_LC_4_19_6  (
            .in0(N__23039),
            .in1(N__29684),
            .in2(N__24868),
            .in3(N__22673),
            .lcout(\c0.n3_adj_2249 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_700_LC_4_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_700_LC_4_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_700_LC_4_19_7 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_700_LC_4_19_7  (
            .in0(N__22493),
            .in1(N__25179),
            .in2(_gnd_net_),
            .in3(N__23035),
            .lcout(\c0.n9393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i6_LC_4_20_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i6_LC_4_20_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i6_LC_4_20_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i6_LC_4_20_0  (
            .in0(N__33181),
            .in1(N__32946),
            .in2(_gnd_net_),
            .in3(N__18979),
            .lcout(\c0.FRAME_MATCHER_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50403),
            .ce(),
            .sr(N__20392));
    defparam \c0.i10768_2_lut_3_lut_4_lut_LC_4_21_0 .C_ON=1'b0;
    defparam \c0.i10768_2_lut_3_lut_4_lut_LC_4_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10768_2_lut_3_lut_4_lut_LC_4_21_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10768_2_lut_3_lut_4_lut_LC_4_21_0  (
            .in0(N__23430),
            .in1(N__23256),
            .in2(N__25080),
            .in3(N__23056),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_2 ),
            .ltout(\c0.FRAME_MATCHER_i_31_N_1312_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_2_i3_2_lut_LC_4_21_1 .C_ON=1'b0;
    defparam \c0.select_238_Select_2_i3_2_lut_LC_4_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_2_i3_2_lut_LC_4_21_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.select_238_Select_2_i3_2_lut_LC_4_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18781),
            .in3(N__29649),
            .lcout(\c0.n3_adj_2259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i2_LC_4_21_2 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i2_LC_4_21_2 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i2_LC_4_21_2 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i2_LC_4_21_2  (
            .in0(N__32848),
            .in1(N__33254),
            .in2(_gnd_net_),
            .in3(N__18856),
            .lcout(\c0.FRAME_MATCHER_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50409),
            .ce(),
            .sr(N__18931));
    defparam \c0.i1_2_lut_3_lut_adj_681_LC_4_21_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_681_LC_4_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_681_LC_4_21_3 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_681_LC_4_21_3  (
            .in0(N__25066),
            .in1(N__21641),
            .in2(_gnd_net_),
            .in3(N__18913),
            .lcout(n16896),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_627_LC_4_21_4 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_627_LC_4_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_627_LC_4_21_4 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \c0.i1_3_lut_adj_627_LC_4_21_4  (
            .in0(N__32690),
            .in1(N__18919),
            .in2(_gnd_net_),
            .in3(N__23714),
            .lcout(\c0.n16895 ),
            .ltout(\c0.n16895_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_651_LC_4_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_651_LC_4_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_651_LC_4_21_5 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_651_LC_4_21_5  (
            .in0(_gnd_net_),
            .in1(N__21640),
            .in2(N__18907),
            .in3(N__25062),
            .lcout(n16897),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10769_2_lut_3_lut_4_lut_LC_4_21_6 .C_ON=1'b0;
    defparam \c0.i10769_2_lut_3_lut_4_lut_LC_4_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10769_2_lut_3_lut_4_lut_LC_4_21_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10769_2_lut_3_lut_4_lut_LC_4_21_6  (
            .in0(N__23429),
            .in1(N__23257),
            .in2(N__21652),
            .in3(N__23057),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_1 ),
            .ltout(\c0.FRAME_MATCHER_i_31_N_1312_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_1_i3_2_lut_LC_4_21_7 .C_ON=1'b0;
    defparam \c0.select_238_Select_1_i3_2_lut_LC_4_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_1_i3_2_lut_LC_4_21_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.select_238_Select_1_i3_2_lut_LC_4_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18904),
            .in3(N__29648),
            .lcout(\c0.n3_adj_2260 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_2_lut_LC_4_22_0 .C_ON=1'b1;
    defparam \c0.add_997_2_lut_LC_4_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_2_lut_LC_4_22_0 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_997_2_lut_LC_4_22_0  (
            .in0(N__29574),
            .in1(N__19371),
            .in2(N__32709),
            .in3(N__18889),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_0 ),
            .ltout(),
            .carryin(bfn_4_22_0_),
            .carryout(\c0.n15622 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_3_lut_LC_4_22_1 .C_ON=1'b1;
    defparam \c0.add_997_3_lut_LC_4_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_3_lut_LC_4_22_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_3_lut_LC_4_22_1  (
            .in0(N__18886),
            .in1(N__21642),
            .in2(N__19439),
            .in3(N__18865),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_1 ),
            .ltout(),
            .carryin(\c0.n15622 ),
            .carryout(\c0.n15623 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_4_lut_LC_4_22_2 .C_ON=1'b1;
    defparam \c0.add_997_4_lut_LC_4_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_4_lut_LC_4_22_2 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_997_4_lut_LC_4_22_2  (
            .in0(N__18862),
            .in1(N__19375),
            .in2(N__25073),
            .in3(N__18850),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_2 ),
            .ltout(),
            .carryin(\c0.n15623 ),
            .carryout(\c0.n15624 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_5_lut_LC_4_22_3 .C_ON=1'b1;
    defparam \c0.add_997_5_lut_LC_4_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_5_lut_LC_4_22_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_5_lut_LC_4_22_3  (
            .in0(N__18847),
            .in1(N__25122),
            .in2(N__19440),
            .in3(N__19006),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_3 ),
            .ltout(),
            .carryin(\c0.n15624 ),
            .carryout(\c0.n15625 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_6_lut_LC_4_22_4 .C_ON=1'b1;
    defparam \c0.add_997_6_lut_LC_4_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_6_lut_LC_4_22_4 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_997_6_lut_LC_4_22_4  (
            .in0(N__19003),
            .in1(N__19379),
            .in2(N__24511),
            .in3(N__18997),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_4 ),
            .ltout(),
            .carryin(\c0.n15625 ),
            .carryout(\c0.n15626 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_7_lut_LC_4_22_5 .C_ON=1'b1;
    defparam \c0.add_997_7_lut_LC_4_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_7_lut_LC_4_22_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_7_lut_LC_4_22_5  (
            .in0(N__18994),
            .in1(N__24433),
            .in2(N__19441),
            .in3(N__18982),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_5 ),
            .ltout(),
            .carryin(\c0.n15626 ),
            .carryout(\c0.n15627 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_8_lut_LC_4_22_6 .C_ON=1'b1;
    defparam \c0.add_997_8_lut_LC_4_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_8_lut_LC_4_22_6 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_997_8_lut_LC_4_22_6  (
            .in0(N__20398),
            .in1(N__19383),
            .in2(N__21925),
            .in3(N__18970),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_6 ),
            .ltout(),
            .carryin(\c0.n15627 ),
            .carryout(\c0.n15628 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_9_lut_LC_4_22_7 .C_ON=1'b1;
    defparam \c0.add_997_9_lut_LC_4_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_9_lut_LC_4_22_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_9_lut_LC_4_22_7  (
            .in0(N__20257),
            .in1(N__21880),
            .in2(N__19442),
            .in3(N__18967),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_7 ),
            .ltout(),
            .carryin(\c0.n15628 ),
            .carryout(\c0.n15629 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_10_lut_LC_4_23_0 .C_ON=1'b1;
    defparam \c0.add_997_10_lut_LC_4_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_10_lut_LC_4_23_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_10_lut_LC_4_23_0  (
            .in0(N__20434),
            .in1(N__24847),
            .in2(N__19443),
            .in3(N__18955),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_8 ),
            .ltout(),
            .carryin(bfn_4_23_0_),
            .carryout(\c0.n15630 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_11_lut_LC_4_23_1 .C_ON=1'b1;
    defparam \c0.add_997_11_lut_LC_4_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_11_lut_LC_4_23_1 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_997_11_lut_LC_4_23_1  (
            .in0(N__20452),
            .in1(N__19390),
            .in2(N__21855),
            .in3(N__18940),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_9 ),
            .ltout(),
            .carryin(\c0.n15630 ),
            .carryout(\c0.n15631 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_12_lut_LC_4_23_2 .C_ON=1'b1;
    defparam \c0.add_997_12_lut_LC_4_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_12_lut_LC_4_23_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_12_lut_LC_4_23_2  (
            .in0(N__20338),
            .in1(N__28184),
            .in2(N__19444),
            .in3(N__18937),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_10 ),
            .ltout(),
            .carryin(\c0.n15631 ),
            .carryout(\c0.n15632 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_13_lut_LC_4_23_3 .C_ON=1'b1;
    defparam \c0.add_997_13_lut_LC_4_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_13_lut_LC_4_23_3 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_997_13_lut_LC_4_23_3  (
            .in0(N__20359),
            .in1(N__19394),
            .in2(N__28322),
            .in3(N__18934),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_11 ),
            .ltout(),
            .carryin(\c0.n15632 ),
            .carryout(\c0.n15633 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_14_lut_LC_4_23_4 .C_ON=1'b1;
    defparam \c0.add_997_14_lut_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_14_lut_LC_4_23_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_14_lut_LC_4_23_4  (
            .in0(N__19096),
            .in1(N__25469),
            .in2(N__19445),
            .in3(N__19087),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_12 ),
            .ltout(),
            .carryin(\c0.n15633 ),
            .carryout(\c0.n15634 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_15_lut_LC_4_23_5 .C_ON=1'b1;
    defparam \c0.add_997_15_lut_LC_4_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_15_lut_LC_4_23_5 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_997_15_lut_LC_4_23_5  (
            .in0(N__19084),
            .in1(N__19398),
            .in2(N__24349),
            .in3(N__19069),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_13 ),
            .ltout(),
            .carryin(\c0.n15634 ),
            .carryout(\c0.n15635 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_16_lut_LC_4_23_6 .C_ON=1'b1;
    defparam \c0.add_997_16_lut_LC_4_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_16_lut_LC_4_23_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_16_lut_LC_4_23_6  (
            .in0(N__19066),
            .in1(N__28282),
            .in2(N__19446),
            .in3(N__19048),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_14 ),
            .ltout(),
            .carryin(\c0.n15635 ),
            .carryout(\c0.n15636 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_17_lut_LC_4_23_7 .C_ON=1'b1;
    defparam \c0.add_997_17_lut_LC_4_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_17_lut_LC_4_23_7 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_997_17_lut_LC_4_23_7  (
            .in0(N__19045),
            .in1(N__19402),
            .in2(N__28254),
            .in3(N__19030),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_15 ),
            .ltout(),
            .carryin(\c0.n15636 ),
            .carryout(\c0.n15637 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_18_lut_LC_4_24_0 .C_ON=1'b1;
    defparam \c0.add_997_18_lut_LC_4_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_18_lut_LC_4_24_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_18_lut_LC_4_24_0  (
            .in0(N__23077),
            .in1(N__22752),
            .in2(N__19450),
            .in3(N__19027),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_16 ),
            .ltout(),
            .carryin(bfn_4_24_0_),
            .carryout(\c0.n15638 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_19_lut_LC_4_24_1 .C_ON=1'b1;
    defparam \c0.add_997_19_lut_LC_4_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_19_lut_LC_4_24_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_19_lut_LC_4_24_1  (
            .in0(N__23440),
            .in1(N__28081),
            .in2(N__19454),
            .in3(N__19024),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_17 ),
            .ltout(),
            .carryin(\c0.n15638 ),
            .carryout(\c0.n15639 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_20_lut_LC_4_24_2 .C_ON=1'b1;
    defparam \c0.add_997_20_lut_LC_4_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_20_lut_LC_4_24_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_20_lut_LC_4_24_2  (
            .in0(N__22258),
            .in1(N__23483),
            .in2(N__19451),
            .in3(N__19021),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_18 ),
            .ltout(),
            .carryin(\c0.n15639 ),
            .carryout(\c0.n15640 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_21_lut_LC_4_24_3 .C_ON=1'b1;
    defparam \c0.add_997_21_lut_LC_4_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_21_lut_LC_4_24_3 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_997_21_lut_LC_4_24_3  (
            .in0(N__20428),
            .in1(N__19420),
            .in2(N__21519),
            .in3(N__19009),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_19 ),
            .ltout(),
            .carryin(\c0.n15640 ),
            .carryout(\c0.n15641 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_22_lut_LC_4_24_4 .C_ON=1'b1;
    defparam \c0.add_997_22_lut_LC_4_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_22_lut_LC_4_24_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_22_lut_LC_4_24_4  (
            .in0(N__20422),
            .in1(N__24546),
            .in2(N__19452),
            .in3(N__19216),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_20 ),
            .ltout(),
            .carryin(\c0.n15641 ),
            .carryout(\c0.n15642 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_23_lut_LC_4_24_5 .C_ON=1'b1;
    defparam \c0.add_997_23_lut_LC_4_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_23_lut_LC_4_24_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_23_lut_LC_4_24_5  (
            .in0(N__20416),
            .in1(N__24403),
            .in2(N__19455),
            .in3(N__19198),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_21 ),
            .ltout(),
            .carryin(\c0.n15642 ),
            .carryout(\c0.n15643 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_24_lut_LC_4_24_6 .C_ON=1'b1;
    defparam \c0.add_997_24_lut_LC_4_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_24_lut_LC_4_24_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_24_lut_LC_4_24_6  (
            .in0(N__20458),
            .in1(N__24761),
            .in2(N__19453),
            .in3(N__19183),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_22 ),
            .ltout(),
            .carryin(\c0.n15643 ),
            .carryout(\c0.n15644 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_25_lut_LC_4_24_7 .C_ON=1'b1;
    defparam \c0.add_997_25_lut_LC_4_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_25_lut_LC_4_24_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_25_lut_LC_4_24_7  (
            .in0(N__20407),
            .in1(N__24722),
            .in2(N__19456),
            .in3(N__19165),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_23 ),
            .ltout(),
            .carryin(\c0.n15644 ),
            .carryout(\c0.n15645 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_26_lut_LC_4_25_0 .C_ON=1'b1;
    defparam \c0.add_997_26_lut_LC_4_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_26_lut_LC_4_25_0 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_997_26_lut_LC_4_25_0  (
            .in0(N__20470),
            .in1(N__19403),
            .in2(N__21472),
            .in3(N__19153),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_24 ),
            .ltout(),
            .carryin(bfn_4_25_0_),
            .carryout(\c0.n15646 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_27_lut_LC_4_25_1 .C_ON=1'b1;
    defparam \c0.add_997_27_lut_LC_4_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_27_lut_LC_4_25_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_27_lut_LC_4_25_1  (
            .in0(N__20482),
            .in1(N__24667),
            .in2(N__19447),
            .in3(N__19144),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_25 ),
            .ltout(),
            .carryin(\c0.n15646 ),
            .carryout(\c0.n15647 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_28_lut_LC_4_25_2 .C_ON=1'b1;
    defparam \c0.add_997_28_lut_LC_4_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_28_lut_LC_4_25_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_28_lut_LC_4_25_2  (
            .in0(N__20464),
            .in1(N__24818),
            .in2(N__19436),
            .in3(N__19129),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_26 ),
            .ltout(),
            .carryin(\c0.n15647 ),
            .carryout(\c0.n15648 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_29_lut_LC_4_25_3 .C_ON=1'b1;
    defparam \c0.add_997_29_lut_LC_4_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_29_lut_LC_4_25_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_29_lut_LC_4_25_3  (
            .in0(N__20518),
            .in1(N__24955),
            .in2(N__19448),
            .in3(N__19114),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_27 ),
            .ltout(),
            .carryin(\c0.n15648 ),
            .carryout(\c0.n15649 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_30_lut_LC_4_25_4 .C_ON=1'b1;
    defparam \c0.add_997_30_lut_LC_4_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_30_lut_LC_4_25_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_30_lut_LC_4_25_4  (
            .in0(N__20476),
            .in1(N__25017),
            .in2(N__19437),
            .in3(N__19099),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_28 ),
            .ltout(),
            .carryin(\c0.n15649 ),
            .carryout(\c0.n15650 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_31_lut_LC_4_25_5 .C_ON=1'b1;
    defparam \c0.add_997_31_lut_LC_4_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_31_lut_LC_4_25_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_31_lut_LC_4_25_5  (
            .in0(N__22123),
            .in1(N__22162),
            .in2(N__19449),
            .in3(N__19513),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_29 ),
            .ltout(),
            .carryin(\c0.n15650 ),
            .carryout(\c0.n15651 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_32_lut_LC_4_25_6 .C_ON=1'b1;
    defparam \c0.add_997_32_lut_LC_4_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_32_lut_LC_4_25_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_997_32_lut_LC_4_25_6  (
            .in0(N__20488),
            .in1(N__24907),
            .in2(N__19438),
            .in3(N__19498),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_30 ),
            .ltout(),
            .carryin(\c0.n15651 ),
            .carryout(\c0.n15652 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_997_33_lut_LC_4_25_7 .C_ON=1'b0;
    defparam \c0.add_997_33_lut_LC_4_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_997_33_lut_LC_4_25_7 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \c0.add_997_33_lut_LC_4_25_7  (
            .in0(N__19413),
            .in1(N__22500),
            .in2(N__20572),
            .in3(N__19495),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1280_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14836_4_lut_LC_4_26_0 .C_ON=1'b0;
    defparam \c0.i14836_4_lut_LC_4_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14836_4_lut_LC_4_26_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i14836_4_lut_LC_4_26_0  (
            .in0(N__22048),
            .in1(N__22099),
            .in2(N__26207),
            .in3(N__22073),
            .lcout(),
            .ltout(\c0.n17274_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_424_LC_4_26_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_424_LC_4_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_424_LC_4_26_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i3_4_lut_adj_424_LC_4_26_1  (
            .in0(N__19540),
            .in1(N__19475),
            .in2(N__19459),
            .in3(N__19597),
            .lcout(\c0.n9490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__1__2264_LC_4_26_2 .C_ON=1'b0;
    defparam \c0.data_in_2__1__2264_LC_4_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__1__2264_LC_4_26_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_in_2__1__2264_LC_4_26_2  (
            .in0(N__27672),
            .in1(_gnd_net_),
            .in2(N__19251),
            .in3(N__19271),
            .lcout(data_in_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50450),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15448_1_lut_LC_4_26_3 .C_ON=1'b0;
    defparam \c0.rx.i15448_1_lut_LC_4_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15448_1_lut_LC_4_26_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.rx.i15448_1_lut_LC_4_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27671),
            .lcout(\c0.n17889 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_433_LC_4_26_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_433_LC_4_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_433_LC_4_26_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i5_4_lut_adj_433_LC_4_26_4  (
            .in0(N__19273),
            .in1(N__20610),
            .in2(N__19250),
            .in3(N__19610),
            .lcout(\c0.n12_adj_2158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i80_LC_4_26_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i80_LC_4_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i80_LC_4_26_5 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i80_LC_4_26_5  (
            .in0(N__28764),
            .in1(N__23625),
            .in2(N__26539),
            .in3(N__31141),
            .lcout(\c0.data_in_frame_9_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50450),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__4__2261_LC_4_26_6 .C_ON=1'b0;
    defparam \c0.data_in_2__4__2261_LC_4_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__4__2261_LC_4_26_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_2__4__2261_LC_4_26_6  (
            .in0(N__22049),
            .in1(_gnd_net_),
            .in2(N__27713),
            .in3(N__19611),
            .lcout(data_in_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50450),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__4__2269_LC_4_26_7 .C_ON=1'b0;
    defparam \c0.data_in_1__4__2269_LC_4_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__4__2269_LC_4_26_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_1__4__2269_LC_4_26_7  (
            .in0(N__19612),
            .in1(N__27673),
            .in2(_gnd_net_),
            .in3(N__19598),
            .lcout(data_in_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50450),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i53_LC_4_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i53_LC_4_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i53_LC_4_27_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i53_LC_4_27_0  (
            .in0(N__31796),
            .in1(N__25992),
            .in2(_gnd_net_),
            .in3(N__25712),
            .lcout(data_in_frame_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50460),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i4_LC_4_27_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i4_LC_4_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i4_LC_4_27_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.tx2.r_Clock_Count__i4_LC_4_27_1  (
            .in0(N__19562),
            .in1(N__19582),
            .in2(_gnd_net_),
            .in3(N__31525),
            .lcout(r_Clock_Count_4_adj_2450),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50460),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i56_LC_4_27_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i56_LC_4_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i56_LC_4_27_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i56_LC_4_27_2  (
            .in0(N__26532),
            .in1(N__26049),
            .in2(_gnd_net_),
            .in3(N__25713),
            .lcout(data_in_frame_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50460),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__0__2257_LC_4_27_3 .C_ON=1'b0;
    defparam \c0.data_in_3__0__2257_LC_4_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__0__2257_LC_4_27_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_in_3__0__2257_LC_4_27_3  (
            .in0(N__27711),
            .in1(_gnd_net_),
            .in2(N__25589),
            .in3(N__22106),
            .lcout(data_in_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50460),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__3__2262_LC_4_27_4 .C_ON=1'b0;
    defparam \c0.data_in_2__3__2262_LC_4_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__3__2262_LC_4_27_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_2__3__2262_LC_4_27_4  (
            .in0(N__25801),
            .in1(N__19543),
            .in2(_gnd_net_),
            .in3(N__27712),
            .lcout(data_in_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50460),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i51_LC_4_27_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i51_LC_4_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i51_LC_4_27_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i51_LC_4_27_5  (
            .in0(N__26562),
            .in1(N__26911),
            .in2(_gnd_net_),
            .in3(N__25711),
            .lcout(data_in_frame_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50460),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i60_LC_4_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i60_LC_4_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i60_LC_4_27_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i60_LC_4_27_6  (
            .in0(N__30522),
            .in1(N__20850),
            .in2(_gnd_net_),
            .in3(N__28953),
            .lcout(data_in_frame_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50460),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_3_lut_4_lut_LC_4_27_7 .C_ON=1'b0;
    defparam \c0.tx2.i2_3_lut_4_lut_LC_4_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_3_lut_4_lut_LC_4_27_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx2.i2_3_lut_4_lut_LC_4_27_7  (
            .in0(N__31028),
            .in1(N__31524),
            .in2(N__27259),
            .in3(N__29341),
            .lcout(\c0.tx2.n8737 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i6_LC_4_28_0 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i6_LC_4_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i6_LC_4_28_0 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \c0.rx.r_Clock_Count__i6_LC_4_28_0  (
            .in0(N__19696),
            .in1(N__19659),
            .in2(_gnd_net_),
            .in3(N__20158),
            .lcout(r_Clock_Count_6_adj_2431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50472),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_678_LC_4_28_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_678_LC_4_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_678_LC_4_28_1 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_678_LC_4_28_1  (
            .in0(N__32710),
            .in1(N__25086),
            .in2(N__21658),
            .in3(N__31988),
            .lcout(n16893),
            .ltout(n16893_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i62_LC_4_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i62_LC_4_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i62_LC_4_28_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_frame_0__i62_LC_4_28_2  (
            .in0(N__31217),
            .in1(_gnd_net_),
            .in2(N__19633),
            .in3(N__28908),
            .lcout(data_in_frame_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50472),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i0_LC_4_28_3 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i0_LC_4_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i0_LC_4_28_3 .LUT_INIT=16'b1010101001000100;
    LogicCell40 \c0.tx.r_Bit_Index_i0_LC_4_28_3  (
            .in0(N__20811),
            .in1(N__24063),
            .in2(_gnd_net_),
            .in3(N__19753),
            .lcout(\c0.tx.r_Bit_Index_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50472),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i13_LC_4_28_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i13_LC_4_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i13_LC_4_28_5 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i13_LC_4_28_5  (
            .in0(N__28802),
            .in1(N__28568),
            .in2(N__31830),
            .in3(N__31989),
            .lcout(\c0.data_in_frame_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50472),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i54_LC_4_28_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i54_LC_4_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i54_LC_4_28_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i54_LC_4_28_6  (
            .in0(N__31216),
            .in1(N__28851),
            .in2(_gnd_net_),
            .in3(N__25715),
            .lcout(data_in_frame_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50472),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i52_LC_4_28_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i52_LC_4_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i52_LC_4_28_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i52_LC_4_28_7  (
            .in0(N__30523),
            .in1(N__26016),
            .in2(_gnd_net_),
            .in3(N__25714),
            .lcout(data_in_frame_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50472),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i9_3_lut_LC_4_29_0 .C_ON=1'b0;
    defparam \c0.tx.i9_3_lut_LC_4_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i9_3_lut_LC_4_29_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.i9_3_lut_LC_4_29_0  (
            .in0(N__24044),
            .in1(N__20818),
            .in2(_gnd_net_),
            .in3(N__31735),
            .lcout(n5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i6_LC_4_29_2 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i6_LC_4_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i6_LC_4_29_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i6_LC_4_29_2  (
            .in0(N__19827),
            .in1(N__23971),
            .in2(_gnd_net_),
            .in3(N__19624),
            .lcout(r_Clock_Count_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50485),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i14756_4_lut_LC_4_29_3 .C_ON=1'b0;
    defparam \c0.tx2.i14756_4_lut_LC_4_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i14756_4_lut_LC_4_29_3 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \c0.tx2.i14756_4_lut_LC_4_29_3  (
            .in0(N__31022),
            .in1(N__29321),
            .in2(N__31546),
            .in3(N__20005),
            .lcout(n17194),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_52_i4_2_lut_LC_4_29_4 .C_ON=1'b0;
    defparam \c0.rx.equal_52_i4_2_lut_LC_4_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_52_i4_2_lut_LC_4_29_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.rx.equal_52_i4_2_lut_LC_4_29_4  (
            .in0(N__19962),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19926),
            .lcout(n4_adj_2417),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_2_lut_4_lut_LC_4_29_5 .C_ON=1'b0;
    defparam \c0.tx.i2_2_lut_4_lut_LC_4_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_2_lut_4_lut_LC_4_29_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx.i2_2_lut_4_lut_LC_4_29_5  (
            .in0(N__19873),
            .in1(N__19826),
            .in2(N__24170),
            .in3(N__19802),
            .lcout(n9937),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i13245_2_lut_LC_4_29_6 .C_ON=1'b0;
    defparam \c0.tx.i13245_2_lut_LC_4_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i13245_2_lut_LC_4_29_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx.i13245_2_lut_LC_4_29_6  (
            .in0(_gnd_net_),
            .in1(N__20808),
            .in2(_gnd_net_),
            .in3(N__31383),
            .lcout(),
            .ltout(\c0.tx.n15683_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i2_LC_4_29_7 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i2_LC_4_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i2_LC_4_29_7 .LUT_INIT=16'b1010101001001000;
    LogicCell40 \c0.tx.r_Bit_Index_i2_LC_4_29_7  (
            .in0(N__20763),
            .in1(N__24045),
            .in2(N__19756),
            .in3(N__19748),
            .lcout(\c0.tx.r_Bit_Index_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50485),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_483_LC_4_30_0 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_483_LC_4_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_483_LC_4_30_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i8_4_lut_adj_483_LC_4_30_0  (
            .in0(N__26725),
            .in1(N__21220),
            .in2(N__20923),
            .in3(N__26668),
            .lcout(\c0.n20_adj_2267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i4_LC_4_30_1 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i4_LC_4_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i4_LC_4_30_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Clock_Count__i4_LC_4_30_1  (
            .in0(N__23962),
            .in1(N__19732),
            .in2(_gnd_net_),
            .in3(N__19721),
            .lcout(r_Clock_Count_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50495),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_461_LC_4_30_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_461_LC_4_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_461_LC_4_30_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_461_LC_4_30_2  (
            .in0(_gnd_net_),
            .in1(N__21359),
            .in2(_gnd_net_),
            .in3(N__21326),
            .lcout(\c0.n12993 ),
            .ltout(\c0.n12993_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14838_4_lut_LC_4_30_3 .C_ON=1'b0;
    defparam \c0.i14838_4_lut_LC_4_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14838_4_lut_LC_4_30_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14838_4_lut_LC_4_30_3  (
            .in0(N__21291),
            .in1(N__21129),
            .in2(N__19699),
            .in3(N__21066),
            .lcout(\c0.n17276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_462_LC_4_30_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_462_LC_4_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_462_LC_4_30_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_462_LC_4_30_4  (
            .in0(_gnd_net_),
            .in1(N__20876),
            .in2(_gnd_net_),
            .in3(N__21167),
            .lcout(\c0.n13298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i3_LC_4_30_5 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i3_LC_4_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i3_LC_4_30_5 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \c0.delay_counter_i0_i3_LC_4_30_5  (
            .in0(N__21168),
            .in1(N__27552),
            .in2(N__21154),
            .in3(N__20983),
            .lcout(\c0.delay_counter_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50495),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i4_LC_4_30_6 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i4_LC_4_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i4_LC_4_30_6 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \c0.delay_counter_i0_i4_LC_4_30_6  (
            .in0(N__20984),
            .in1(N__26669),
            .in2(N__21142),
            .in3(N__27559),
            .lcout(\c0.delay_counter_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50495),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i11_LC_4_30_7 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i11_LC_4_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i11_LC_4_30_7 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \c0.delay_counter_i0_i11_LC_4_30_7  (
            .in0(N__21327),
            .in1(N__27551),
            .in2(N__21313),
            .in3(N__20982),
            .lcout(\c0.delay_counter_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50495),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i1_LC_4_31_1 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i1_LC_4_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i1_LC_4_31_1 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \c0.delay_counter_i0_i1_LC_4_31_1  (
            .in0(N__27534),
            .in1(N__20860),
            .in2(N__20881),
            .in3(N__20985),
            .lcout(\c0.delay_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50507),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i5_LC_4_31_2 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i5_LC_4_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i5_LC_4_31_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.delay_counter_i0_i5_LC_4_31_2  (
            .in0(N__20987),
            .in1(N__21106),
            .in2(_gnd_net_),
            .in3(N__21130),
            .lcout(\c0.delay_counter_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50507),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_1_lut_LC_4_31_4.C_ON=1'b0;
    defparam i3_1_lut_LC_4_31_4.SEQ_MODE=4'b0000;
    defparam i3_1_lut_LC_4_31_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 i3_1_lut_LC_4_31_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27533),
            .lcout(n53),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_491_LC_4_31_5 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_491_LC_4_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_491_LC_4_31_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i9_4_lut_adj_491_LC_4_31_5  (
            .in0(N__21064),
            .in1(N__20032),
            .in2(N__21290),
            .in3(N__20025),
            .lcout(),
            .ltout(\c0.n21_adj_2271_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_adj_540_LC_4_31_6 .C_ON=1'b0;
    defparam \c0.i11_3_lut_adj_540_LC_4_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_adj_540_LC_4_31_6 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \c0.i11_3_lut_adj_540_LC_4_31_6  (
            .in0(_gnd_net_),
            .in1(N__20014),
            .in2(N__20008),
            .in3(N__20173),
            .lcout(n29),
            .ltout(n29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i9_LC_4_31_7 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i9_LC_4_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i9_LC_4_31_7 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \c0.delay_counter_i0_i9_LC_4_31_7  (
            .in0(N__21001),
            .in1(N__21019),
            .in2(N__20194),
            .in3(N__20986),
            .lcout(\c0.delay_counter_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50507),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_32_0 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_32_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_32_0  (
            .in0(N__20073),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(tx_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_464_LC_4_32_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_464_LC_4_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_464_LC_4_32_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i1_2_lut_adj_464_LC_4_32_1  (
            .in0(N__21097),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21017),
            .lcout(\c0.n12991 ),
            .ltout(\c0.n12991_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_489_LC_4_32_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_489_LC_4_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_489_LC_4_32_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_489_LC_4_32_2  (
            .in0(N__26649),
            .in1(N__21127),
            .in2(N__20176),
            .in3(N__26699),
            .lcout(\c0.n19_adj_2270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_LC_4_32_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_LC_4_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_LC_4_32_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \c0.i1_3_lut_4_lut_LC_4_32_3  (
            .in0(N__42592),
            .in1(N__46362),
            .in2(N__45952),
            .in3(N__27402),
            .lcout(n9361),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i1_LC_4_32_5 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i1_LC_4_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i1_LC_4_32_5 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \c0.tx.r_SM_Main_i1_LC_4_32_5  (
            .in0(N__24038),
            .in1(N__23964),
            .in2(N__24187),
            .in3(N__24115),
            .lcout(r_SM_Main_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50517),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i0_LC_4_32_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i0_LC_4_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i0_LC_4_32_6 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \c0.rx.r_Clock_Count__i0_LC_4_32_6  (
            .in0(N__20167),
            .in1(N__20096),
            .in2(_gnd_net_),
            .in3(N__20154),
            .lcout(r_Clock_Count_0_adj_2437),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50517),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_45_LC_4_32_7 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_45_LC_4_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.o_Tx_Serial_45_LC_4_32_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.tx.o_Tx_Serial_45_LC_4_32_7  (
            .in0(N__20734),
            .in1(N__23963),
            .in2(_gnd_net_),
            .in3(N__20072),
            .lcout(tx_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50517),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i3_LC_5_13_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i3_LC_5_13_3 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i3_LC_5_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i3_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(N__33397),
            .in2(_gnd_net_),
            .in3(N__34652),
            .lcout(\c0.FRAME_MATCHER_state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50416),
            .ce(),
            .sr(N__21187));
    defparam \c0.data_in_0__0__2281_LC_5_17_0 .C_ON=1'b0;
    defparam \c0.data_in_0__0__2281_LC_5_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__0__2281_LC_5_17_0 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_in_0__0__2281_LC_5_17_0  (
            .in0(N__27800),
            .in1(_gnd_net_),
            .in2(N__22205),
            .in3(N__20059),
            .lcout(data_in_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50386),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10680_2_lut_LC_5_17_1 .C_ON=1'b0;
    defparam \c0.i10680_2_lut_LC_5_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10680_2_lut_LC_5_17_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i10680_2_lut_LC_5_17_1  (
            .in0(_gnd_net_),
            .in1(N__22496),
            .in2(_gnd_net_),
            .in3(N__25180),
            .lcout(n3977),
            .ltout(n3977_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i2_LC_5_17_2 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i2_LC_5_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_state_i2_LC_5_17_2 .LUT_INIT=16'b1011101111111011;
    LogicCell40 \c0.FRAME_MATCHER_state_i2_LC_5_17_2  (
            .in0(N__21403),
            .in1(N__32447),
            .in2(N__20236),
            .in3(N__32996),
            .lcout(FRAME_MATCHER_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50386),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_LC_5_17_4 .C_ON=1'b0;
    defparam \c0.i3_3_lut_LC_5_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_LC_5_17_4 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \c0.i3_3_lut_LC_5_17_4  (
            .in0(N__32299),
            .in1(N__33476),
            .in2(_gnd_net_),
            .in3(N__29475),
            .lcout(\c0.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_21_i3_2_lut_3_lut_4_lut_LC_5_17_5 .C_ON=1'b0;
    defparam \c0.select_238_Select_21_i3_2_lut_3_lut_4_lut_LC_5_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_21_i3_2_lut_3_lut_4_lut_LC_5_17_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_21_i3_2_lut_3_lut_4_lut_LC_5_17_5  (
            .in0(N__22691),
            .in1(N__29712),
            .in2(N__24388),
            .in3(N__23044),
            .lcout(\c0.n3_adj_2233 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_28_i3_2_lut_3_lut_4_lut_LC_5_17_6 .C_ON=1'b0;
    defparam \c0.select_238_Select_28_i3_2_lut_3_lut_4_lut_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_28_i3_2_lut_3_lut_4_lut_LC_5_17_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_28_i3_2_lut_3_lut_4_lut_LC_5_17_6  (
            .in0(N__23045),
            .in1(N__24997),
            .in2(N__29732),
            .in3(N__22690),
            .lcout(\c0.n3_adj_2219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i6_LC_5_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i6_LC_5_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i6_LC_5_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i6_LC_5_18_0  (
            .in0(_gnd_net_),
            .in1(N__21774),
            .in2(_gnd_net_),
            .in3(N__34564),
            .lcout(\c0.FRAME_MATCHER_state_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50398),
            .ce(),
            .sr(N__20218));
    defparam \c0.FRAME_MATCHER_state_i4_LC_5_19_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i4_LC_5_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i4_LC_5_19_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i4_LC_5_19_0  (
            .in0(_gnd_net_),
            .in1(N__30018),
            .in2(_gnd_net_),
            .in3(N__34561),
            .lcout(\c0.FRAME_MATCHER_state_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50404),
            .ce(),
            .sr(N__29836));
    defparam \c0.select_238_Select_23_i3_2_lut_3_lut_4_lut_LC_5_20_0 .C_ON=1'b0;
    defparam \c0.select_238_Select_23_i3_2_lut_3_lut_4_lut_LC_5_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_23_i3_2_lut_3_lut_4_lut_LC_5_20_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_23_i3_2_lut_3_lut_4_lut_LC_5_20_0  (
            .in0(N__29657),
            .in1(N__22667),
            .in2(N__24726),
            .in3(N__23059),
            .lcout(\c0.n3_adj_2229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14770_3_lut_LC_5_20_1.C_ON=1'b0;
    defparam i14770_3_lut_LC_5_20_1.SEQ_MODE=4'b0000;
    defparam i14770_3_lut_LC_5_20_1.LUT_INIT=16'b1111111111011101;
    LogicCell40 i14770_3_lut_LC_5_20_1 (
            .in0(N__32306),
            .in1(N__37387),
            .in2(_gnd_net_),
            .in3(N__21811),
            .lcout(n17208),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_22_i3_2_lut_3_lut_4_lut_LC_5_20_2 .C_ON=1'b0;
    defparam \c0.select_238_Select_22_i3_2_lut_3_lut_4_lut_LC_5_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_22_i3_2_lut_3_lut_4_lut_LC_5_20_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_22_i3_2_lut_3_lut_4_lut_LC_5_20_2  (
            .in0(N__29656),
            .in1(N__22665),
            .in2(N__24772),
            .in3(N__23058),
            .lcout(\c0.n3_adj_2231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_24_i3_2_lut_3_lut_4_lut_LC_5_20_3 .C_ON=1'b0;
    defparam \c0.select_238_Select_24_i3_2_lut_3_lut_4_lut_LC_5_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_24_i3_2_lut_3_lut_4_lut_LC_5_20_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_24_i3_2_lut_3_lut_4_lut_LC_5_20_3  (
            .in0(N__23060),
            .in1(N__21466),
            .in2(N__22700),
            .in3(N__29658),
            .lcout(\c0.n3_adj_2227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_26_i3_2_lut_3_lut_4_lut_LC_5_20_4 .C_ON=1'b0;
    defparam \c0.select_238_Select_26_i3_2_lut_3_lut_4_lut_LC_5_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_26_i3_2_lut_3_lut_4_lut_LC_5_20_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_26_i3_2_lut_3_lut_4_lut_LC_5_20_4  (
            .in0(N__29660),
            .in1(N__22666),
            .in2(N__24822),
            .in3(N__23062),
            .lcout(\c0.n3_adj_2223 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_25_i3_2_lut_3_lut_4_lut_LC_5_20_5 .C_ON=1'b0;
    defparam \c0.select_238_Select_25_i3_2_lut_3_lut_4_lut_LC_5_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_25_i3_2_lut_3_lut_4_lut_LC_5_20_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_25_i3_2_lut_3_lut_4_lut_LC_5_20_5  (
            .in0(N__23061),
            .in1(N__24682),
            .in2(N__22701),
            .in3(N__29659),
            .lcout(\c0.n3_adj_2225 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11115_2_lut_3_lut_4_lut_LC_5_20_6 .C_ON=1'b0;
    defparam \c0.i11115_2_lut_3_lut_4_lut_LC_5_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11115_2_lut_3_lut_4_lut_LC_5_20_6 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \c0.i11115_2_lut_3_lut_4_lut_LC_5_20_6  (
            .in0(N__33530),
            .in1(N__22015),
            .in2(N__21799),
            .in3(N__32790),
            .lcout(\c0.n1439 ),
            .ltout(\c0.n1439_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_27_i3_2_lut_3_lut_4_lut_LC_5_20_7 .C_ON=1'b0;
    defparam \c0.select_238_Select_27_i3_2_lut_3_lut_4_lut_LC_5_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_27_i3_2_lut_3_lut_4_lut_LC_5_20_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_27_i3_2_lut_3_lut_4_lut_LC_5_20_7  (
            .in0(N__23063),
            .in1(N__22668),
            .in2(N__20275),
            .in3(N__24960),
            .lcout(\c0.n3_adj_2221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10763_2_lut_3_lut_4_lut_LC_5_21_0 .C_ON=1'b0;
    defparam \c0.i10763_2_lut_3_lut_4_lut_LC_5_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10763_2_lut_3_lut_4_lut_LC_5_21_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10763_2_lut_3_lut_4_lut_LC_5_21_0  (
            .in0(N__23422),
            .in1(N__23233),
            .in2(N__21886),
            .in3(N__22971),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i7_LC_5_21_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i7_LC_5_21_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i7_LC_5_21_1 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i7_LC_5_21_1  (
            .in0(N__33195),
            .in1(N__32803),
            .in2(_gnd_net_),
            .in3(N__20251),
            .lcout(\c0.FRAME_MATCHER_i_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50417),
            .ce(),
            .sr(N__20245));
    defparam \c0.select_238_Select_7_i3_2_lut_3_lut_4_lut_LC_5_21_2 .C_ON=1'b0;
    defparam \c0.select_238_Select_7_i3_2_lut_3_lut_4_lut_LC_5_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_7_i3_2_lut_3_lut_4_lut_LC_5_21_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_7_i3_2_lut_3_lut_4_lut_LC_5_21_2  (
            .in0(N__22695),
            .in1(N__21884),
            .in2(N__29707),
            .in3(N__22979),
            .lcout(\c0.n3_adj_2250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10764_2_lut_3_lut_4_lut_LC_5_21_3 .C_ON=1'b0;
    defparam \c0.i10764_2_lut_3_lut_4_lut_LC_5_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10764_2_lut_3_lut_4_lut_LC_5_21_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10764_2_lut_3_lut_4_lut_LC_5_21_3  (
            .in0(N__23234),
            .in1(N__21905),
            .in2(N__23042),
            .in3(N__23421),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_6_i3_2_lut_3_lut_4_lut_LC_5_21_4 .C_ON=1'b0;
    defparam \c0.select_238_Select_6_i3_2_lut_3_lut_4_lut_LC_5_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_6_i3_2_lut_3_lut_4_lut_LC_5_21_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_6_i3_2_lut_3_lut_4_lut_LC_5_21_4  (
            .in0(N__22696),
            .in1(N__21906),
            .in2(N__29706),
            .in3(N__22978),
            .lcout(\c0.n3_adj_2253 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_12_i3_2_lut_3_lut_4_lut_LC_5_21_5 .C_ON=1'b0;
    defparam \c0.select_238_Select_12_i3_2_lut_3_lut_4_lut_LC_5_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_12_i3_2_lut_3_lut_4_lut_LC_5_21_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_12_i3_2_lut_3_lut_4_lut_LC_5_21_5  (
            .in0(N__22975),
            .in1(N__29661),
            .in2(N__25477),
            .in3(N__22694),
            .lcout(\c0.n3_adj_2245 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_19_i3_2_lut_3_lut_4_lut_LC_5_21_6 .C_ON=1'b0;
    defparam \c0.select_238_Select_19_i3_2_lut_3_lut_4_lut_LC_5_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_19_i3_2_lut_3_lut_4_lut_LC_5_21_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_19_i3_2_lut_3_lut_4_lut_LC_5_21_6  (
            .in0(N__22693),
            .in1(N__21514),
            .in2(N__29705),
            .in3(N__22976),
            .lcout(\c0.n3_adj_2237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_20_i3_2_lut_3_lut_4_lut_LC_5_21_7 .C_ON=1'b0;
    defparam \c0.select_238_Select_20_i3_2_lut_3_lut_4_lut_LC_5_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_20_i3_2_lut_3_lut_4_lut_LC_5_21_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_20_i3_2_lut_3_lut_4_lut_LC_5_21_7  (
            .in0(N__22977),
            .in1(N__29665),
            .in2(N__24545),
            .in3(N__22692),
            .lcout(\c0.n3_adj_2235 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10759_2_lut_3_lut_4_lut_LC_5_22_0 .C_ON=1'b0;
    defparam \c0.i10759_2_lut_3_lut_4_lut_LC_5_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10759_2_lut_3_lut_4_lut_LC_5_22_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10759_2_lut_3_lut_4_lut_LC_5_22_0  (
            .in0(N__23367),
            .in1(N__23202),
            .in2(N__28323),
            .in3(N__22915),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i11_LC_5_22_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i11_LC_5_22_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i11_LC_5_22_1 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i11_LC_5_22_1  (
            .in0(N__32826),
            .in1(N__33182),
            .in2(_gnd_net_),
            .in3(N__20353),
            .lcout(\c0.FRAME_MATCHER_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50426),
            .ce(),
            .sr(N__20347));
    defparam \c0.select_238_Select_11_i3_2_lut_3_lut_4_lut_LC_5_22_2 .C_ON=1'b0;
    defparam \c0.select_238_Select_11_i3_2_lut_3_lut_4_lut_LC_5_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_11_i3_2_lut_3_lut_4_lut_LC_5_22_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_11_i3_2_lut_3_lut_4_lut_LC_5_22_2  (
            .in0(N__22699),
            .in1(N__29709),
            .in2(N__28324),
            .in3(N__22926),
            .lcout(\c0.n3_adj_2246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10760_2_lut_3_lut_4_lut_LC_5_22_3 .C_ON=1'b0;
    defparam \c0.i10760_2_lut_3_lut_4_lut_LC_5_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10760_2_lut_3_lut_4_lut_LC_5_22_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10760_2_lut_3_lut_4_lut_LC_5_22_3  (
            .in0(N__23203),
            .in1(N__28185),
            .in2(N__22993),
            .in3(N__23364),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_10_i3_2_lut_3_lut_4_lut_LC_5_22_4 .C_ON=1'b0;
    defparam \c0.select_238_Select_10_i3_2_lut_3_lut_4_lut_LC_5_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_10_i3_2_lut_3_lut_4_lut_LC_5_22_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_10_i3_2_lut_3_lut_4_lut_LC_5_22_4  (
            .in0(N__22697),
            .in1(N__29708),
            .in2(N__28189),
            .in3(N__22925),
            .lcout(\c0.n3_adj_2247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10761_2_lut_3_lut_4_lut_LC_5_22_5 .C_ON=1'b0;
    defparam \c0.i10761_2_lut_3_lut_4_lut_LC_5_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10761_2_lut_3_lut_4_lut_LC_5_22_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10761_2_lut_3_lut_4_lut_LC_5_22_5  (
            .in0(N__23204),
            .in1(N__21851),
            .in2(N__22994),
            .in3(N__23365),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_9_i3_2_lut_3_lut_4_lut_LC_5_22_6 .C_ON=1'b0;
    defparam \c0.select_238_Select_9_i3_2_lut_3_lut_4_lut_LC_5_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_9_i3_2_lut_3_lut_4_lut_LC_5_22_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_9_i3_2_lut_3_lut_4_lut_LC_5_22_6  (
            .in0(N__22698),
            .in1(N__29710),
            .in2(N__21856),
            .in3(N__22927),
            .lcout(\c0.n3_adj_2248 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10762_2_lut_3_lut_4_lut_LC_5_22_7 .C_ON=1'b0;
    defparam \c0.i10762_2_lut_3_lut_4_lut_LC_5_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10762_2_lut_3_lut_4_lut_LC_5_22_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10762_2_lut_3_lut_4_lut_LC_5_22_7  (
            .in0(N__23205),
            .in1(N__24860),
            .in2(N__22995),
            .in3(N__23366),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10751_2_lut_3_lut_4_lut_LC_5_23_0 .C_ON=1'b0;
    defparam \c0.i10751_2_lut_3_lut_4_lut_LC_5_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10751_2_lut_3_lut_4_lut_LC_5_23_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10751_2_lut_3_lut_4_lut_LC_5_23_0  (
            .in0(N__23188),
            .in1(N__21520),
            .in2(N__22989),
            .in3(N__23378),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10750_2_lut_3_lut_4_lut_LC_5_23_1 .C_ON=1'b0;
    defparam \c0.i10750_2_lut_3_lut_4_lut_LC_5_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10750_2_lut_3_lut_4_lut_LC_5_23_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10750_2_lut_3_lut_4_lut_LC_5_23_1  (
            .in0(N__23377),
            .in1(N__23187),
            .in2(N__24550),
            .in3(N__22891),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10749_2_lut_3_lut_4_lut_LC_5_23_2 .C_ON=1'b0;
    defparam \c0.i10749_2_lut_3_lut_4_lut_LC_5_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10749_2_lut_3_lut_4_lut_LC_5_23_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10749_2_lut_3_lut_4_lut_LC_5_23_2  (
            .in0(N__23186),
            .in1(N__24402),
            .in2(N__22988),
            .in3(N__23376),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10747_2_lut_3_lut_4_lut_LC_5_23_3 .C_ON=1'b0;
    defparam \c0.i10747_2_lut_3_lut_4_lut_LC_5_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10747_2_lut_3_lut_4_lut_LC_5_23_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10747_2_lut_3_lut_4_lut_LC_5_23_3  (
            .in0(N__23375),
            .in1(N__23185),
            .in2(N__24727),
            .in3(N__22887),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_454_LC_5_23_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_454_LC_5_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_454_LC_5_23_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_454_LC_5_23_5  (
            .in0(N__23581),
            .in1(N__22371),
            .in2(N__25294),
            .in3(N__22183),
            .lcout(),
            .ltout(\c0.n18_adj_2198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_456_LC_5_23_6 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_456_LC_5_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_456_LC_5_23_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i10_4_lut_adj_456_LC_5_23_6  (
            .in0(N__23494),
            .in1(N__20581),
            .in2(N__20401),
            .in3(N__22213),
            .lcout(\c0.n127_adj_2136 ),
            .ltout(\c0.n127_adj_2136_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10568_2_lut_3_lut_4_lut_LC_5_23_7 .C_ON=1'b0;
    defparam \c0.i10568_2_lut_3_lut_4_lut_LC_5_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10568_2_lut_3_lut_4_lut_LC_5_23_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10568_2_lut_3_lut_4_lut_LC_5_23_7  (
            .in0(N__32691),
            .in1(N__23184),
            .in2(N__20521),
            .in3(N__22886),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10743_2_lut_3_lut_4_lut_LC_5_24_0 .C_ON=1'b0;
    defparam \c0.i10743_2_lut_3_lut_4_lut_LC_5_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10743_2_lut_3_lut_4_lut_LC_5_24_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10743_2_lut_3_lut_4_lut_LC_5_24_0  (
            .in0(N__23370),
            .in1(N__23197),
            .in2(N__24961),
            .in3(N__22904),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i3_LC_5_24_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i3_LC_5_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i3_LC_5_24_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i3_LC_5_24_1  (
            .in0(N__20563),
            .in1(N__33758),
            .in2(N__30487),
            .in3(N__20512),
            .lcout(rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50441),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10736_2_lut_3_lut_4_lut_LC_5_24_2 .C_ON=1'b0;
    defparam \c0.i10736_2_lut_3_lut_4_lut_LC_5_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10736_2_lut_3_lut_4_lut_LC_5_24_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10736_2_lut_3_lut_4_lut_LC_5_24_2  (
            .in0(N__23368),
            .in1(N__23195),
            .in2(N__24913),
            .in3(N__22902),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10745_2_lut_3_lut_4_lut_LC_5_24_3 .C_ON=1'b0;
    defparam \c0.i10745_2_lut_3_lut_4_lut_LC_5_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10745_2_lut_3_lut_4_lut_LC_5_24_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10745_2_lut_3_lut_4_lut_LC_5_24_3  (
            .in0(N__23199),
            .in1(N__24680),
            .in2(N__22990),
            .in3(N__23374),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10742_2_lut_3_lut_4_lut_LC_5_24_4 .C_ON=1'b0;
    defparam \c0.i10742_2_lut_3_lut_4_lut_LC_5_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10742_2_lut_3_lut_4_lut_LC_5_24_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10742_2_lut_3_lut_4_lut_LC_5_24_4  (
            .in0(N__23369),
            .in1(N__23196),
            .in2(N__25018),
            .in3(N__22903),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10746_2_lut_3_lut_4_lut_LC_5_24_5 .C_ON=1'b0;
    defparam \c0.i10746_2_lut_3_lut_4_lut_LC_5_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10746_2_lut_3_lut_4_lut_LC_5_24_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10746_2_lut_3_lut_4_lut_LC_5_24_5  (
            .in0(N__23200),
            .in1(N__21471),
            .in2(N__22991),
            .in3(N__23373),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10744_2_lut_3_lut_4_lut_LC_5_24_6 .C_ON=1'b0;
    defparam \c0.i10744_2_lut_3_lut_4_lut_LC_5_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10744_2_lut_3_lut_4_lut_LC_5_24_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10744_2_lut_3_lut_4_lut_LC_5_24_6  (
            .in0(N__23371),
            .in1(N__23198),
            .in2(N__24823),
            .in3(N__22905),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10748_2_lut_3_lut_4_lut_LC_5_24_7 .C_ON=1'b0;
    defparam \c0.i10748_2_lut_3_lut_4_lut_LC_5_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10748_2_lut_3_lut_4_lut_LC_5_24_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10748_2_lut_3_lut_4_lut_LC_5_24_7  (
            .in0(N__23201),
            .in1(N__24768),
            .in2(N__22992),
            .in3(N__23372),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_425_LC_5_25_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_425_LC_5_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_425_LC_5_25_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_425_LC_5_25_0  (
            .in0(N__29085),
            .in1(N__28977),
            .in2(N__23734),
            .in3(N__25969),
            .lcout(\c0.n9743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_698_LC_5_25_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_698_LC_5_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_698_LC_5_25_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_698_LC_5_25_1  (
            .in0(N__23605),
            .in1(N__26152),
            .in2(N__22418),
            .in3(N__25860),
            .lcout(\c0.n12_adj_2200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_437_LC_5_25_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_437_LC_5_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_437_LC_5_25_2 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.i2_3_lut_adj_437_LC_5_25_2  (
            .in0(N__26151),
            .in1(N__22409),
            .in2(_gnd_net_),
            .in3(N__23604),
            .lcout(\c0.n9493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__7__2266_LC_5_25_3 .C_ON=1'b0;
    defparam \c0.data_in_1__7__2266_LC_5_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__7__2266_LC_5_25_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_1__7__2266_LC_5_25_3  (
            .in0(N__27761),
            .in1(N__25861),
            .in2(_gnd_net_),
            .in3(N__23535),
            .lcout(data_in_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50451),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__2__2255_LC_5_25_4 .C_ON=1'b0;
    defparam \c0.data_in_3__2__2255_LC_5_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__2__2255_LC_5_25_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__2__2255_LC_5_25_4  (
            .in0(N__26901),
            .in1(N__27762),
            .in2(_gnd_net_),
            .in3(N__26203),
            .lcout(data_in_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50451),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10733_2_lut_3_lut_4_lut_LC_5_25_5 .C_ON=1'b0;
    defparam \c0.i10733_2_lut_3_lut_4_lut_LC_5_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10733_2_lut_3_lut_4_lut_LC_5_25_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10733_2_lut_3_lut_4_lut_LC_5_25_5  (
            .in0(N__23240),
            .in1(N__23402),
            .in2(N__22501),
            .in3(N__23016),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__4__2253_LC_5_25_6 .C_ON=1'b0;
    defparam \c0.data_in_3__4__2253_LC_5_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__4__2253_LC_5_25_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__4__2253_LC_5_25_6  (
            .in0(N__31795),
            .in1(N__27763),
            .in2(_gnd_net_),
            .in3(N__22053),
            .lcout(data_in_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50451),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_40_i8_2_lut_3_lut_LC_5_25_7 .C_ON=1'b0;
    defparam \c0.equal_40_i8_2_lut_3_lut_LC_5_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.equal_40_i8_2_lut_3_lut_LC_5_25_7 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.equal_40_i8_2_lut_3_lut_LC_5_25_7  (
            .in0(N__21633),
            .in1(N__32704),
            .in2(_gnd_net_),
            .in3(N__25085),
            .lcout(\c0.n8_adj_2310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i2_LC_5_26_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i2_LC_5_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i2_LC_5_26_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i2_LC_5_26_0  (
            .in0(N__20562),
            .in1(N__33759),
            .in2(N__26918),
            .in3(N__20646),
            .lcout(rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50461),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i4_LC_5_26_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i4_LC_5_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i4_LC_5_26_1 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i4_LC_5_26_1  (
            .in0(N__20647),
            .in1(N__31794),
            .in2(N__33766),
            .in3(N__20535),
            .lcout(rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50461),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i16_LC_5_26_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i16_LC_5_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i16_LC_5_26_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i16_LC_5_26_2  (
            .in0(N__31995),
            .in1(N__28762),
            .in2(N__28611),
            .in3(N__26525),
            .lcout(\c0.data_in_frame_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50461),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__2__2279_LC_5_26_3 .C_ON=1'b0;
    defparam \c0.data_in_0__2__2279_LC_5_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__2__2279_LC_5_26_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0__2__2279_LC_5_26_3  (
            .in0(N__27768),
            .in1(N__26150),
            .in2(_gnd_net_),
            .in3(N__20611),
            .lcout(data_in_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50461),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__3__2278_LC_5_26_4 .C_ON=1'b0;
    defparam \c0.data_in_0__3__2278_LC_5_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__3__2278_LC_5_26_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0__3__2278_LC_5_26_4  (
            .in0(N__20599),
            .in1(N__23511),
            .in2(_gnd_net_),
            .in3(N__27769),
            .lcout(data_in_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50461),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i9_LC_5_26_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i9_LC_5_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i9_LC_5_26_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i9_LC_5_26_5  (
            .in0(N__28761),
            .in1(N__25594),
            .in2(N__26436),
            .in3(N__31997),
            .lcout(\c0.data_in_frame_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50461),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i22_LC_5_26_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i22_LC_5_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i22_LC_5_26_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i22_LC_5_26_6  (
            .in0(N__31996),
            .in1(N__31877),
            .in2(N__31229),
            .in3(N__26286),
            .lcout(\c0.data_in_frame_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50461),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i12_LC_5_26_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i12_LC_5_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i12_LC_5_26_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i12_LC_5_26_7  (
            .in0(N__28760),
            .in1(N__30505),
            .in2(N__28524),
            .in3(N__31994),
            .lcout(\c0.data_in_frame_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50461),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i24_LC_5_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i24_LC_5_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i24_LC_5_27_0 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i24_LC_5_27_0  (
            .in0(N__31918),
            .in1(N__23811),
            .in2(N__26537),
            .in3(N__31991),
            .lcout(\c0.data_in_frame_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50473),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_435_LC_5_27_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_435_LC_5_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_435_LC_5_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_435_LC_5_27_1  (
            .in0(N__23745),
            .in1(N__28393),
            .in2(_gnd_net_),
            .in3(N__28514),
            .lcout(\c0.n15939 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i17_LC_5_27_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i17_LC_5_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i17_LC_5_27_2 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i17_LC_5_27_2  (
            .in0(N__31917),
            .in1(N__30219),
            .in2(N__25593),
            .in3(N__31990),
            .lcout(\c0.data_in_frame_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50473),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_423_LC_5_27_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_423_LC_5_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_423_LC_5_27_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_423_LC_5_27_3  (
            .in0(_gnd_net_),
            .in1(N__28561),
            .in2(_gnd_net_),
            .in3(N__28513),
            .lcout(\c0.n17004 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i6_LC_5_27_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i6_LC_5_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i6_LC_5_27_4 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.rx.r_Rx_Byte_i6_LC_5_27_4  (
            .in0(N__25638),
            .in1(N__20725),
            .in2(N__33765),
            .in3(N__20640),
            .lcout(rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50473),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_585_LC_5_27_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_585_LC_5_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_585_LC_5_27_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_585_LC_5_27_6  (
            .in0(N__24453),
            .in1(N__24509),
            .in2(N__25140),
            .in3(N__23721),
            .lcout(\c0.n16891 ),
            .ltout(\c0.n16891_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i14_LC_5_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i14_LC_5_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i14_LC_5_27_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i14_LC_5_27_7  (
            .in0(N__28785),
            .in1(N__31212),
            .in2(N__20701),
            .in3(N__26249),
            .lcout(\c0.data_in_frame_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50473),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i63_LC_5_28_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i63_LC_5_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i63_LC_5_28_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i63_LC_5_28_0  (
            .in0(N__20848),
            .in1(N__25639),
            .in2(_gnd_net_),
            .in3(N__25749),
            .lcout(data_in_frame_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50486),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i59_LC_5_28_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i59_LC_5_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i59_LC_5_28_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i59_LC_5_28_1  (
            .in0(N__26577),
            .in1(N__26919),
            .in2(_gnd_net_),
            .in3(N__20847),
            .lcout(data_in_frame_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50486),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i11_LC_5_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i11_LC_5_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i11_LC_5_28_2 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i11_LC_5_28_2  (
            .in0(N__28801),
            .in1(N__28397),
            .in2(N__26932),
            .in3(N__31993),
            .lcout(\c0.data_in_frame_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50486),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_396_LC_5_28_4 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_396_LC_5_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_396_LC_5_28_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i1_2_lut_adj_396_LC_5_28_4  (
            .in0(_gnd_net_),
            .in1(N__20698),
            .in2(_gnd_net_),
            .in3(N__20662),
            .lcout(n9477),
            .ltout(n9477_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i0_LC_5_28_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i0_LC_5_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i0_LC_5_28_5 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.rx.r_Rx_Byte_i0_LC_5_28_5  (
            .in0(N__25562),
            .in1(N__20629),
            .in2(N__20614),
            .in3(N__33746),
            .lcout(rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50486),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i64_LC_5_28_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i64_LC_5_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i64_LC_5_28_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i64_LC_5_28_6  (
            .in0(N__20849),
            .in1(N__26521),
            .in2(_gnd_net_),
            .in3(N__26070),
            .lcout(data_in_frame_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50486),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i58_LC_5_28_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i58_LC_5_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i58_LC_5_28_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i58_LC_5_28_7  (
            .in0(N__30683),
            .in1(N__26322),
            .in2(_gnd_net_),
            .in3(N__20846),
            .lcout(data_in_frame_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50486),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i61_LC_5_29_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i61_LC_5_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i61_LC_5_29_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i61_LC_5_29_0  (
            .in0(N__31812),
            .in1(N__26304),
            .in2(_gnd_net_),
            .in3(N__20851),
            .lcout(data_in_frame_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50496),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i13_LC_5_29_1 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i13_LC_5_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i13_LC_5_29_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.delay_counter_i0_i13_LC_5_29_1  (
            .in0(N__21247),
            .in1(N__26732),
            .in2(_gnd_net_),
            .in3(N__20989),
            .lcout(\c0.delay_counter_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50496),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i15371_4_lut_LC_5_29_2 .C_ON=1'b0;
    defparam \c0.tx.i15371_4_lut_LC_5_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i15371_4_lut_LC_5_29_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx.i15371_4_lut_LC_5_29_2  (
            .in0(N__24104),
            .in1(N__20761),
            .in2(N__31384),
            .in3(N__20809),
            .lcout(\c0.tx.n17462 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i0_LC_5_29_3 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i0_LC_5_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i0_LC_5_29_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.delay_counter_i0_i0_LC_5_29_3  (
            .in0(N__20893),
            .in1(N__20928),
            .in2(_gnd_net_),
            .in3(N__20988),
            .lcout(\c0.delay_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50496),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_5_29_4 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_5_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_5_29_4 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_5_29_4  (
            .in0(N__20810),
            .in1(N__31315),
            .in2(N__20764),
            .in3(N__20776),
            .lcout(),
            .ltout(\c0.tx.n17975_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.n17975_bdd_4_lut_LC_5_29_5 .C_ON=1'b0;
    defparam \c0.tx.n17975_bdd_4_lut_LC_5_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.n17975_bdd_4_lut_LC_5_29_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.tx.n17975_bdd_4_lut_LC_5_29_5  (
            .in0(N__20762),
            .in1(N__29419),
            .in2(N__20740),
            .in3(N__23833),
            .lcout(),
            .ltout(\c0.tx.o_Tx_Serial_N_2064_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_5_29_6 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_5_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_5_29_6 .LUT_INIT=16'b1100110011110011;
    LogicCell40 \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_5_29_6  (
            .in0(_gnd_net_),
            .in1(N__24067),
            .in2(N__20737),
            .in3(N__24173),
            .lcout(n3_adj_2406),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i2_LC_5_30_0 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i2_LC_5_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i2_LC_5_30_0 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \c0.delay_counter_i0_i2_LC_5_30_0  (
            .in0(N__20977),
            .in1(N__21178),
            .in2(N__26650),
            .in3(N__27556),
            .lcout(\c0.delay_counter_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50508),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i10_LC_5_30_1 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i10_LC_5_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i10_LC_5_30_1 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \c0.delay_counter_i0_i10_LC_5_30_1  (
            .in0(N__21363),
            .in1(N__21343),
            .in2(N__27573),
            .in3(N__20976),
            .lcout(\c0.delay_counter_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50508),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i14_LC_5_30_2 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i14_LC_5_30_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i14_LC_5_30_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.delay_counter_i0_i14_LC_5_30_2  (
            .in0(N__20980),
            .in1(_gnd_net_),
            .in2(N__21199),
            .in3(N__21233),
            .lcout(\c0.delay_counter_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50508),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_616_LC_5_30_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_616_LC_5_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_616_LC_5_30_3 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \c0.i1_3_lut_adj_616_LC_5_30_3  (
            .in0(N__35761),
            .in1(N__45924),
            .in2(_gnd_net_),
            .in3(N__24196),
            .lcout(\c0.n1419 ),
            .ltout(\c0.n1419_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i6_LC_5_30_4 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i6_LC_5_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i6_LC_5_30_4 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \c0.delay_counter_i0_i6_LC_5_30_4  (
            .in0(N__21076),
            .in1(N__21096),
            .in2(N__20992),
            .in3(N__27557),
            .lcout(\c0.delay_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50508),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i12_LC_5_30_5 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i12_LC_5_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i12_LC_5_30_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.delay_counter_i0_i12_LC_5_30_5  (
            .in0(N__21259),
            .in1(N__21289),
            .in2(_gnd_net_),
            .in3(N__20979),
            .lcout(\c0.delay_counter_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50508),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i8_LC_5_30_6 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i8_LC_5_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i8_LC_5_30_6 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \c0.delay_counter_i0_i8_LC_5_30_6  (
            .in0(N__20978),
            .in1(N__26698),
            .in2(N__21034),
            .in3(N__27558),
            .lcout(\c0.delay_counter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50508),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i7_LC_5_30_7 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i7_LC_5_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i7_LC_5_30_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.delay_counter_i0_i7_LC_5_30_7  (
            .in0(N__21043),
            .in1(N__21067),
            .in2(_gnd_net_),
            .in3(N__20981),
            .lcout(\c0.delay_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50508),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_2_lut_LC_5_31_0 .C_ON=1'b1;
    defparam \c0.add_2495_2_lut_LC_5_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_2_lut_LC_5_31_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \c0.add_2495_2_lut_LC_5_31_0  (
            .in0(N__20935),
            .in1(N__20924),
            .in2(_gnd_net_),
            .in3(N__20884),
            .lcout(\c0.n17637 ),
            .ltout(),
            .carryin(bfn_5_31_0_),
            .carryout(\c0.n15514 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_3_lut_LC_5_31_1 .C_ON=1'b1;
    defparam \c0.add_2495_3_lut_LC_5_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_3_lut_LC_5_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2495_3_lut_LC_5_31_1  (
            .in0(_gnd_net_),
            .in1(N__20877),
            .in2(_gnd_net_),
            .in3(N__20854),
            .lcout(\c0.n6531 ),
            .ltout(),
            .carryin(\c0.n15514 ),
            .carryout(\c0.n15515 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_4_lut_LC_5_31_2 .C_ON=1'b1;
    defparam \c0.add_2495_4_lut_LC_5_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_4_lut_LC_5_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2495_4_lut_LC_5_31_2  (
            .in0(_gnd_net_),
            .in1(N__26635),
            .in2(_gnd_net_),
            .in3(N__21172),
            .lcout(\c0.n6530 ),
            .ltout(),
            .carryin(\c0.n15515 ),
            .carryout(\c0.n15516 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_5_lut_LC_5_31_3 .C_ON=1'b1;
    defparam \c0.add_2495_5_lut_LC_5_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_5_lut_LC_5_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2495_5_lut_LC_5_31_3  (
            .in0(_gnd_net_),
            .in1(N__21169),
            .in2(_gnd_net_),
            .in3(N__21145),
            .lcout(\c0.n6529 ),
            .ltout(),
            .carryin(\c0.n15516 ),
            .carryout(\c0.n15517 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_6_lut_LC_5_31_4 .C_ON=1'b1;
    defparam \c0.add_2495_6_lut_LC_5_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_6_lut_LC_5_31_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2495_6_lut_LC_5_31_4  (
            .in0(_gnd_net_),
            .in1(N__26670),
            .in2(_gnd_net_),
            .in3(N__21133),
            .lcout(\c0.n6528 ),
            .ltout(),
            .carryin(\c0.n15517 ),
            .carryout(\c0.n15518 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_7_lut_LC_5_31_5 .C_ON=1'b1;
    defparam \c0.add_2495_7_lut_LC_5_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_7_lut_LC_5_31_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2495_7_lut_LC_5_31_5  (
            .in0(N__27569),
            .in1(N__21128),
            .in2(_gnd_net_),
            .in3(N__21100),
            .lcout(\c0.n17574 ),
            .ltout(),
            .carryin(\c0.n15518 ),
            .carryout(\c0.n15519 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_8_lut_LC_5_31_6 .C_ON=1'b1;
    defparam \c0.add_2495_8_lut_LC_5_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_8_lut_LC_5_31_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2495_8_lut_LC_5_31_6  (
            .in0(_gnd_net_),
            .in1(N__21095),
            .in2(_gnd_net_),
            .in3(N__21070),
            .lcout(\c0.n6526 ),
            .ltout(),
            .carryin(\c0.n15519 ),
            .carryout(\c0.n15520 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_9_lut_LC_5_31_7 .C_ON=1'b1;
    defparam \c0.add_2495_9_lut_LC_5_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_9_lut_LC_5_31_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2495_9_lut_LC_5_31_7  (
            .in0(N__27568),
            .in1(N__21065),
            .in2(_gnd_net_),
            .in3(N__21037),
            .lcout(\c0.n17638 ),
            .ltout(),
            .carryin(\c0.n15520 ),
            .carryout(\c0.n15521 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_10_lut_LC_5_32_0 .C_ON=1'b1;
    defparam \c0.add_2495_10_lut_LC_5_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_10_lut_LC_5_32_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2495_10_lut_LC_5_32_0  (
            .in0(_gnd_net_),
            .in1(N__26703),
            .in2(_gnd_net_),
            .in3(N__21022),
            .lcout(\c0.n6524 ),
            .ltout(),
            .carryin(bfn_5_32_0_),
            .carryout(\c0.n15522 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_11_lut_LC_5_32_1 .C_ON=1'b1;
    defparam \c0.add_2495_11_lut_LC_5_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_11_lut_LC_5_32_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2495_11_lut_LC_5_32_1  (
            .in0(_gnd_net_),
            .in1(N__21018),
            .in2(_gnd_net_),
            .in3(N__20995),
            .lcout(\c0.n6523 ),
            .ltout(),
            .carryin(\c0.n15522 ),
            .carryout(\c0.n15523 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_12_lut_LC_5_32_2 .C_ON=1'b1;
    defparam \c0.add_2495_12_lut_LC_5_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_12_lut_LC_5_32_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2495_12_lut_LC_5_32_2  (
            .in0(_gnd_net_),
            .in1(N__21364),
            .in2(_gnd_net_),
            .in3(N__21334),
            .lcout(\c0.n6522 ),
            .ltout(),
            .carryin(\c0.n15523 ),
            .carryout(\c0.n15524 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_13_lut_LC_5_32_3 .C_ON=1'b1;
    defparam \c0.add_2495_13_lut_LC_5_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_13_lut_LC_5_32_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2495_13_lut_LC_5_32_3  (
            .in0(_gnd_net_),
            .in1(N__21331),
            .in2(_gnd_net_),
            .in3(N__21298),
            .lcout(\c0.n6521 ),
            .ltout(),
            .carryin(\c0.n15524 ),
            .carryout(\c0.n15525 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_14_lut_LC_5_32_4 .C_ON=1'b1;
    defparam \c0.add_2495_14_lut_LC_5_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_14_lut_LC_5_32_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2495_14_lut_LC_5_32_4  (
            .in0(N__27549),
            .in1(_gnd_net_),
            .in2(N__21295),
            .in3(N__21250),
            .lcout(\c0.n17575 ),
            .ltout(),
            .carryin(\c0.n15525 ),
            .carryout(\c0.n15526 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_15_lut_LC_5_32_5 .C_ON=1'b1;
    defparam \c0.add_2495_15_lut_LC_5_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_15_lut_LC_5_32_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2495_15_lut_LC_5_32_5  (
            .in0(N__27548),
            .in1(N__26734),
            .in2(_gnd_net_),
            .in3(N__21238),
            .lcout(\c0.n17639 ),
            .ltout(),
            .carryin(\c0.n15526 ),
            .carryout(\c0.n15527 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2495_16_lut_LC_5_32_6 .C_ON=1'b0;
    defparam \c0.add_2495_16_lut_LC_5_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_2495_16_lut_LC_5_32_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2495_16_lut_LC_5_32_6  (
            .in0(N__27550),
            .in1(N__21234),
            .in2(_gnd_net_),
            .in3(N__21202),
            .lcout(\c0.n17635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i29_LC_6_14_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i29_LC_6_14_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i29_LC_6_14_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.FRAME_MATCHER_state_i29_LC_6_14_0  (
            .in0(N__34653),
            .in1(N__21752),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_state_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50418),
            .ce(),
            .sr(N__21532));
    defparam \c0.i1_2_lut_adj_738_LC_6_15_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_738_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_738_LC_6_15_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.i1_2_lut_adj_738_LC_6_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29981),
            .in3(N__24601),
            .lcout(\c0.n16371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_703_LC_6_15_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_703_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_703_LC_6_15_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_703_LC_6_15_6  (
            .in0(_gnd_net_),
            .in1(N__33402),
            .in2(_gnd_net_),
            .in3(N__29968),
            .lcout(\c0.n16331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_719_LC_6_16_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_719_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_719_LC_6_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_719_LC_6_16_0  (
            .in0(_gnd_net_),
            .in1(N__25259),
            .in2(_gnd_net_),
            .in3(N__32590),
            .lcout(\c0.n16453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_4_lut_adj_565_LC_6_16_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_4_lut_adj_565_LC_6_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_4_lut_adj_565_LC_6_16_2 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \c0.i1_4_lut_4_lut_adj_565_LC_6_16_2  (
            .in0(N__33493),
            .in1(N__34281),
            .in2(N__32324),
            .in3(N__33401),
            .lcout(\c0.n8603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_760_LC_6_16_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_760_LC_6_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_760_LC_6_16_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_760_LC_6_16_5  (
            .in0(_gnd_net_),
            .in1(N__21754),
            .in2(_gnd_net_),
            .in3(N__29967),
            .lcout(\c0.n16381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_LC_6_17_0 .C_ON=1'b0;
    defparam \c0.i17_4_lut_LC_6_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_LC_6_17_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i17_4_lut_LC_6_17_0  (
            .in0(N__21518),
            .in1(N__23485),
            .in2(N__21470),
            .in3(N__22726),
            .lcout(\c0.n46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i16_LC_6_17_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i16_LC_6_17_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i16_LC_6_17_1 .LUT_INIT=16'b0101111100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i16_LC_6_17_1  (
            .in0(N__32895),
            .in1(_gnd_net_),
            .in2(N__33097),
            .in3(N__21421),
            .lcout(\c0.FRAME_MATCHER_i_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50392),
            .ce(),
            .sr(N__22576));
    defparam \c0.i1_2_lut_adj_528_LC_6_17_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_528_LC_6_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_528_LC_6_17_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i1_2_lut_adj_528_LC_6_17_2  (
            .in0(N__33478),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22020),
            .lcout(n9452),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10724_3_lut_LC_6_17_3 .C_ON=1'b0;
    defparam \c0.i10724_3_lut_LC_6_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10724_3_lut_LC_6_17_3 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \c0.i10724_3_lut_LC_6_17_3  (
            .in0(N__33517),
            .in1(N__23431),
            .in2(_gnd_net_),
            .in3(N__23225),
            .lcout(),
            .ltout(n1716_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_765_LC_6_17_4.C_ON=1'b0;
    defparam i1_4_lut_adj_765_LC_6_17_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_765_LC_6_17_4.LUT_INIT=16'b1011000000000000;
    LogicCell40 i1_4_lut_adj_765_LC_6_17_4 (
            .in0(N__21397),
            .in1(N__32894),
            .in2(N__21406),
            .in3(N__23043),
            .lcout(n14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_6_17_5.C_ON=1'b0;
    defparam i1_4_lut_LC_6_17_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_6_17_5.LUT_INIT=16'b1100110111111111;
    LogicCell40 i1_4_lut_LC_6_17_5 (
            .in0(N__33053),
            .in1(N__28029),
            .in2(N__21582),
            .in3(N__22353),
            .lcout(n16775),
            .ltout(n16775_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_802_LC_6_17_6.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_802_LC_6_17_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_802_LC_6_17_6.LUT_INIT=16'b1111000111110101;
    LogicCell40 i1_3_lut_4_lut_adj_802_LC_6_17_6 (
            .in0(N__21387),
            .in1(N__27906),
            .in2(N__21367),
            .in3(N__21672),
            .lcout(n16776),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_406_LC_6_17_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_406_LC_6_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_406_LC_6_17_7 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \c0.i1_2_lut_adj_406_LC_6_17_7  (
            .in0(N__22019),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33477),
            .lcout(n9453),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i14_LC_6_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i14_LC_6_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i14_LC_6_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i14_LC_6_18_0  (
            .in0(_gnd_net_),
            .in1(N__29816),
            .in2(_gnd_net_),
            .in3(N__34559),
            .lcout(\c0.FRAME_MATCHER_state_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50405),
            .ce(),
            .sr(N__25426));
    defparam \c0.i10695_4_lut_LC_6_19_0 .C_ON=1'b0;
    defparam \c0.i10695_4_lut_LC_6_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10695_4_lut_LC_6_19_0 .LUT_INIT=16'b0101010101000000;
    LogicCell40 \c0.i10695_4_lut_LC_6_19_0  (
            .in0(N__22492),
            .in1(N__32669),
            .in2(N__21657),
            .in3(N__25175),
            .lcout(n2275),
            .ltout(n2275_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15357_2_lut_3_lut_4_lut_LC_6_19_1 .C_ON=1'b0;
    defparam \c0.i15357_2_lut_3_lut_4_lut_LC_6_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15357_2_lut_3_lut_4_lut_LC_6_19_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.i15357_2_lut_3_lut_4_lut_LC_6_19_1  (
            .in0(N__23224),
            .in1(N__23420),
            .in2(N__21559),
            .in3(N__23040),
            .lcout(\c0.n17454 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4944_2_lut_LC_6_19_2 .C_ON=1'b0;
    defparam \c0.i4944_2_lut_LC_6_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4944_2_lut_LC_6_19_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i4944_2_lut_LC_6_19_2  (
            .in0(_gnd_net_),
            .in1(N__23419),
            .in2(_gnd_net_),
            .in3(N__23223),
            .lcout(\c0.n7212 ),
            .ltout(\c0.n7212_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15395_3_lut_4_lut_LC_6_19_3 .C_ON=1'b0;
    defparam \c0.i15395_3_lut_4_lut_LC_6_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15395_3_lut_4_lut_LC_6_19_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.i15395_3_lut_4_lut_LC_6_19_3  (
            .in0(N__27208),
            .in1(N__27943),
            .in2(N__21556),
            .in3(N__23041),
            .lcout(),
            .ltout(\c0.n17452_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_LC_6_19_4 .C_ON=1'b0;
    defparam \c0.i18_4_lut_LC_6_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_LC_6_19_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \c0.i18_4_lut_LC_6_19_4  (
            .in0(N__33531),
            .in1(N__22024),
            .in2(N__21553),
            .in3(N__21550),
            .lcout(\c0.n7 ),
            .ltout(\c0.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i5_LC_6_19_5 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i5_LC_6_19_5 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i5_LC_6_19_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i5_LC_6_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21544),
            .in3(N__21787),
            .lcout(\c0.FRAME_MATCHER_state_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50410),
            .ce(),
            .sr(N__21541));
    defparam \c0.i1_2_lut_adj_707_LC_6_19_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_707_LC_6_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_707_LC_6_19_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_707_LC_6_19_6  (
            .in0(N__21786),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29920),
            .lcout(\c0.n16335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_467_LC_6_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_467_LC_6_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_467_LC_6_19_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_467_LC_6_19_7  (
            .in0(_gnd_net_),
            .in1(N__21785),
            .in2(_gnd_net_),
            .in3(N__21770),
            .lcout(\c0.n6_adj_2213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_458_LC_6_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_458_LC_6_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_458_LC_6_20_0 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \c0.i1_2_lut_adj_458_LC_6_20_0  (
            .in0(N__25329),
            .in1(N__21753),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n59 ),
            .ltout(\c0.n59_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_476_LC_6_20_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_476_LC_6_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_476_LC_6_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_4_lut_adj_476_LC_6_20_1  (
            .in0(N__29775),
            .in1(N__33412),
            .in2(N__21733),
            .in3(N__24615),
            .lcout(),
            .ltout(\c0.n5_adj_2262_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_479_LC_6_20_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_479_LC_6_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_479_LC_6_20_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_479_LC_6_20_2  (
            .in0(N__28140),
            .in1(N__25366),
            .in2(N__21730),
            .in3(N__24580),
            .lcout(\c0.n16876 ),
            .ltout(\c0.n16876_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_415_LC_6_20_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_415_LC_6_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_415_LC_6_20_3 .LUT_INIT=16'b1111110011111100;
    LogicCell40 \c0.i1_2_lut_adj_415_LC_6_20_3  (
            .in0(_gnd_net_),
            .in1(N__29509),
            .in2(N__21727),
            .in3(_gnd_net_),
            .lcout(\c0.n60 ),
            .ltout(\c0.n60_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14820_4_lut_LC_6_20_4 .C_ON=1'b0;
    defparam \c0.i14820_4_lut_LC_6_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14820_4_lut_LC_6_20_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14820_4_lut_LC_6_20_4  (
            .in0(N__24313),
            .in1(N__21952),
            .in2(N__21724),
            .in3(N__32368),
            .lcout(\c0.n17258 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i23_LC_6_20_5 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i23_LC_6_20_5 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i23_LC_6_20_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i23_LC_6_20_5  (
            .in0(N__34558),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21688),
            .lcout(\c0.FRAME_MATCHER_state_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50419),
            .ce(),
            .sr(N__21721));
    defparam \c0.i1_2_lut_adj_747_LC_6_20_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_747_LC_6_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_747_LC_6_20_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_747_LC_6_20_6  (
            .in0(N__21687),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29919),
            .lcout(\c0.n16363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_635_LC_6_20_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_635_LC_6_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_635_LC_6_20_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i1_2_lut_adj_635_LC_6_20_7  (
            .in0(N__21711),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21686),
            .lcout(\c0.n16898 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_LC_6_21_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_LC_6_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_LC_6_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i4_4_lut_LC_6_21_0  (
            .in0(N__30084),
            .in1(N__30025),
            .in2(N__32341),
            .in3(N__21958),
            .lcout(\c0.n9451 ),
            .ltout(\c0.n9451_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10592_2_lut_3_lut_LC_6_21_1 .C_ON=1'b0;
    defparam \c0.i10592_2_lut_3_lut_LC_6_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10592_2_lut_3_lut_LC_6_21_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.i10592_2_lut_3_lut_LC_6_21_1  (
            .in0(N__27937),
            .in1(_gnd_net_),
            .in2(N__22030),
            .in3(N__33522),
            .lcout(n12933),
            .ltout(n12933_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10929_2_lut_3_lut_4_lut_LC_6_21_2 .C_ON=1'b0;
    defparam \c0.i10929_2_lut_3_lut_4_lut_LC_6_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10929_2_lut_3_lut_4_lut_LC_6_21_2 .LUT_INIT=16'b0000110001001100;
    LogicCell40 \c0.i10929_2_lut_3_lut_4_lut_LC_6_21_2  (
            .in0(N__22009),
            .in1(N__27770),
            .in2(N__22027),
            .in3(N__33534),
            .lcout(\c0.n13272 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i33_3_lut_LC_6_21_3 .C_ON=1'b0;
    defparam \c0.i33_3_lut_LC_6_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i33_3_lut_LC_6_21_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.i33_3_lut_LC_6_21_3  (
            .in0(N__27938),
            .in1(N__33523),
            .in2(_gnd_net_),
            .in3(N__22008),
            .lcout(),
            .ltout(\c0.n28_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_404_LC_6_21_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_404_LC_6_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_404_LC_6_21_4 .LUT_INIT=16'b0010111111111111;
    LogicCell40 \c0.i1_4_lut_adj_404_LC_6_21_4  (
            .in0(N__21985),
            .in1(N__21973),
            .in2(N__21967),
            .in3(N__32783),
            .lcout(n16795),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_LC_6_21_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_LC_6_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_LC_6_21_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_LC_6_21_5  (
            .in0(N__29474),
            .in1(N__24312),
            .in2(_gnd_net_),
            .in3(N__21964),
            .lcout(\c0.n16879 ),
            .ltout(\c0.n16879_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_419_LC_6_21_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_419_LC_6_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_419_LC_6_21_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_419_LC_6_21_6  (
            .in0(N__33521),
            .in1(N__21948),
            .in2(N__21928),
            .in3(N__32367),
            .lcout(n9445),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_LC_6_21_7 .C_ON=1'b0;
    defparam \c0.i21_4_lut_LC_6_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_LC_6_21_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i21_4_lut_LC_6_21_7  (
            .in0(N__21918),
            .in1(N__21885),
            .in2(N__21847),
            .in3(N__22164),
            .lcout(\c0.n50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_422_LC_6_22_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_422_LC_6_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_422_LC_6_22_0 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \c0.i1_2_lut_adj_422_LC_6_22_0  (
            .in0(N__21810),
            .in1(N__32292),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n9488 ),
            .ltout(\c0.n9488_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_436_LC_6_22_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_436_LC_6_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_436_LC_6_22_1 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i1_4_lut_adj_436_LC_6_22_1  (
            .in0(N__25837),
            .in1(N__22240),
            .in2(N__22228),
            .in3(N__22225),
            .lcout(\c0.n9485 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_740_LC_6_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_740_LC_6_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_740_LC_6_22_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_740_LC_6_22_2  (
            .in0(_gnd_net_),
            .in1(N__27990),
            .in2(_gnd_net_),
            .in3(N__29893),
            .lcout(\c0.n16369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14802_2_lut_LC_6_22_3 .C_ON=1'b0;
    defparam \c0.i14802_2_lut_LC_6_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14802_2_lut_LC_6_22_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i14802_2_lut_LC_6_22_3  (
            .in0(N__26144),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23611),
            .lcout(\c0.n17240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__1__2280_LC_6_22_4 .C_ON=1'b0;
    defparam \c0.data_in_0__1__2280_LC_6_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__1__2280_LC_6_22_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0__1__2280_LC_6_22_4  (
            .in0(N__22426),
            .in1(N__27782),
            .in2(_gnd_net_),
            .in3(N__25292),
            .lcout(data_in_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50434),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14818_4_lut_LC_6_22_5 .C_ON=1'b0;
    defparam \c0.i14818_4_lut_LC_6_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i14818_4_lut_LC_6_22_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i14818_4_lut_LC_6_22_5  (
            .in0(N__22207),
            .in1(N__25925),
            .in2(N__25828),
            .in3(N__27609),
            .lcout(\c0.n17256 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_410_LC_6_22_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_410_LC_6_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_410_LC_6_22_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i4_4_lut_adj_410_LC_6_22_6  (
            .in0(N__27608),
            .in1(N__22206),
            .in2(N__25929),
            .in3(N__22182),
            .lcout(),
            .ltout(\c0.n10_adj_2149_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_LC_6_22_7 .C_ON=1'b0;
    defparam \c0.i5_4_lut_LC_6_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_LC_6_22_7 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \c0.i5_4_lut_LC_6_22_7  (
            .in0(N__25824),
            .in1(N__25270),
            .in2(N__22171),
            .in3(N__23548),
            .lcout(\c0.n9482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10741_2_lut_3_lut_4_lut_LC_6_23_0 .C_ON=1'b0;
    defparam \c0.i10741_2_lut_3_lut_4_lut_LC_6_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10741_2_lut_3_lut_4_lut_LC_6_23_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10741_2_lut_3_lut_4_lut_LC_6_23_0  (
            .in0(N__23354),
            .in1(N__22168),
            .in2(N__22954),
            .in3(N__23182),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_411_LC_6_23_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_411_LC_6_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_411_LC_6_23_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i5_4_lut_adj_411_LC_6_23_1  (
            .in0(N__22111),
            .in1(N__22081),
            .in2(N__22057),
            .in3(N__22383),
            .lcout(),
            .ltout(\c0.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_LC_6_23_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_LC_6_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_LC_6_23_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i6_4_lut_LC_6_23_2  (
            .in0(N__22531),
            .in1(N__22519),
            .in2(N__22504),
            .in3(N__26208),
            .lcout(n127_adj_2418),
            .ltout(n127_adj_2418_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_691_LC_6_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_691_LC_6_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_691_LC_6_23_3 .LUT_INIT=16'b1011000000000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_691_LC_6_23_3  (
            .in0(N__22495),
            .in1(N__25168),
            .in2(N__22435),
            .in3(N__23352),
            .lcout(n9435),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_LC_6_23_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_LC_6_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_LC_6_23_4 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i3_4_lut_LC_6_23_4  (
            .in0(N__22432),
            .in1(N__22425),
            .in2(N__22387),
            .in3(N__22375),
            .lcout(n127),
            .ltout(n127_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_751_LC_6_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_751_LC_6_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_751_LC_6_23_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_751_LC_6_23_5  (
            .in0(N__22349),
            .in1(N__23351),
            .in2(N__22327),
            .in3(N__22856),
            .lcout(\c0.n2 ),
            .ltout(\c0.n2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_LC_6_23_6 .C_ON=1'b0;
    defparam \c0.i1_4_lut_LC_6_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_LC_6_23_6 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \c0.i1_4_lut_LC_6_23_6  (
            .in0(N__32834),
            .in1(N__23183),
            .in2(N__22312),
            .in3(N__22299),
            .lcout(\c0.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4924_2_lut_LC_6_23_7 .C_ON=1'b0;
    defparam \c0.i4924_2_lut_LC_6_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4924_2_lut_LC_6_23_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i4924_2_lut_LC_6_23_7  (
            .in0(_gnd_net_),
            .in1(N__23353),
            .in2(_gnd_net_),
            .in3(N__22855),
            .lcout(n7198),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10752_2_lut_3_lut_4_lut_LC_6_24_0 .C_ON=1'b0;
    defparam \c0.i10752_2_lut_3_lut_4_lut_LC_6_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10752_2_lut_3_lut_4_lut_LC_6_24_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10752_2_lut_3_lut_4_lut_LC_6_24_0  (
            .in0(N__23357),
            .in1(N__23189),
            .in2(N__23484),
            .in3(N__22895),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i18_LC_6_24_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i18_LC_6_24_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i18_LC_6_24_1 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i18_LC_6_24_1  (
            .in0(N__33183),
            .in1(N__32835),
            .in2(_gnd_net_),
            .in3(N__22249),
            .lcout(\c0.FRAME_MATCHER_i_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50452),
            .ce(),
            .sr(N__23449));
    defparam \c0.select_238_Select_18_i3_2_lut_3_lut_4_lut_LC_6_24_2 .C_ON=1'b0;
    defparam \c0.select_238_Select_18_i3_2_lut_3_lut_4_lut_LC_6_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_18_i3_2_lut_3_lut_4_lut_LC_6_24_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_18_i3_2_lut_3_lut_4_lut_LC_6_24_2  (
            .in0(N__22708),
            .in1(N__23479),
            .in2(N__29749),
            .in3(N__22901),
            .lcout(\c0.n3_adj_2239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_764_LC_6_24_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_764_LC_6_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_764_LC_6_24_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_764_LC_6_24_3  (
            .in0(N__22898),
            .in1(_gnd_net_),
            .in2(N__23235),
            .in3(N__23358),
            .lcout(n8828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10753_2_lut_3_lut_4_lut_LC_6_24_4 .C_ON=1'b0;
    defparam \c0.i10753_2_lut_3_lut_4_lut_LC_6_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10753_2_lut_3_lut_4_lut_LC_6_24_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10753_2_lut_3_lut_4_lut_LC_6_24_4  (
            .in0(N__23356),
            .in1(N__23190),
            .in2(N__28082),
            .in3(N__22896),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_17_i3_2_lut_3_lut_4_lut_LC_6_24_5 .C_ON=1'b0;
    defparam \c0.select_238_Select_17_i3_2_lut_3_lut_4_lut_LC_6_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_17_i3_2_lut_3_lut_4_lut_LC_6_24_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_17_i3_2_lut_3_lut_4_lut_LC_6_24_5  (
            .in0(N__22900),
            .in1(N__29745),
            .in2(N__28083),
            .in3(N__22707),
            .lcout(\c0.n3_adj_2240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10754_2_lut_3_lut_4_lut_LC_6_24_6 .C_ON=1'b0;
    defparam \c0.i10754_2_lut_3_lut_4_lut_LC_6_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10754_2_lut_3_lut_4_lut_LC_6_24_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10754_2_lut_3_lut_4_lut_LC_6_24_6  (
            .in0(N__23355),
            .in1(N__23191),
            .in2(N__22753),
            .in3(N__22897),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1312_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_16_i3_2_lut_3_lut_4_lut_LC_6_24_7 .C_ON=1'b0;
    defparam \c0.select_238_Select_16_i3_2_lut_3_lut_4_lut_LC_6_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_16_i3_2_lut_3_lut_4_lut_LC_6_24_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.select_238_Select_16_i3_2_lut_3_lut_4_lut_LC_6_24_7  (
            .in0(N__22899),
            .in1(N__29744),
            .in2(N__22751),
            .in3(N__22706),
            .lcout(\c0.n3_adj_2241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_438_LC_6_25_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_438_LC_6_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_438_LC_6_25_0 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \c0.i5_4_lut_adj_438_LC_6_25_0  (
            .in0(N__29133),
            .in1(N__22564),
            .in2(N__22543),
            .in3(N__26428),
            .lcout(\c0.n21_adj_2171 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i5_LC_6_25_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i5_LC_6_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i5_LC_6_25_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i5_LC_6_25_1  (
            .in0(N__30422),
            .in1(N__31797),
            .in2(_gnd_net_),
            .in3(N__30339),
            .lcout(data_in_frame_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50462),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_420_LC_6_25_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_420_LC_6_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_420_LC_6_25_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_420_LC_6_25_2  (
            .in0(_gnd_net_),
            .in1(N__28603),
            .in2(_gnd_net_),
            .in3(N__26858),
            .lcout(\c0.n17013 ),
            .ltout(\c0.n17013_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_440_LC_6_25_3 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_440_LC_6_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_440_LC_6_25_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_440_LC_6_25_3  (
            .in0(N__23668),
            .in1(N__23781),
            .in2(N__23644),
            .in3(N__26253),
            .lcout(\c0.n17015 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__6__2259_LC_6_25_4 .C_ON=1'b0;
    defparam \c0.data_in_2__6__2259_LC_6_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__6__2259_LC_6_25_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_2__6__2259_LC_6_25_4  (
            .in0(N__23607),
            .in1(_gnd_net_),
            .in2(N__27783),
            .in3(N__27828),
            .lcout(data_in_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50462),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_430_LC_6_25_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_430_LC_6_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_430_LC_6_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_430_LC_6_25_5  (
            .in0(N__23641),
            .in1(N__23782),
            .in2(N__23632),
            .in3(N__26831),
            .lcout(\c0.n17014 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i3_LC_6_25_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i3_LC_6_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i3_LC_6_25_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i3_LC_6_25_6  (
            .in0(N__26910),
            .in1(N__25951),
            .in2(_gnd_net_),
            .in3(N__30421),
            .lcout(data_in_frame_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50462),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__6__2251_LC_6_25_7 .C_ON=1'b0;
    defparam \c0.data_in_3__6__2251_LC_6_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__6__2251_LC_6_25_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__6__2251_LC_6_25_7  (
            .in0(N__25672),
            .in1(N__27764),
            .in2(_gnd_net_),
            .in3(N__23606),
            .lcout(data_in_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50462),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14830_3_lut_LC_6_26_0 .C_ON=1'b0;
    defparam \c0.i14830_3_lut_LC_6_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14830_3_lut_LC_6_26_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i14830_3_lut_LC_6_26_0  (
            .in0(N__23580),
            .in1(N__23507),
            .in2(_gnd_net_),
            .in3(N__23530),
            .lcout(\c0.n17268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i82_LC_6_26_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i82_LC_6_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i82_LC_6_26_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i82_LC_6_26_1  (
            .in0(N__31111),
            .in1(N__30697),
            .in2(N__23797),
            .in3(N__31878),
            .lcout(\c0.data_in_frame_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50474),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i87_LC_6_26_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i87_LC_6_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i87_LC_6_26_2 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i87_LC_6_26_2  (
            .in0(N__31879),
            .in1(N__23764),
            .in2(N__25675),
            .in3(N__31112),
            .lcout(\c0.data_in_frame_10_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50474),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_LC_6_26_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_LC_6_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_LC_6_26_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i8_4_lut_LC_6_26_3  (
            .in0(N__23531),
            .in1(N__25887),
            .in2(N__23512),
            .in3(N__26173),
            .lcout(\c0.n19_adj_2199 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i79_LC_6_26_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i79_LC_6_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i79_LC_6_26_4 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i79_LC_6_26_4  (
            .in0(N__28763),
            .in1(N__23680),
            .in2(N__25674),
            .in3(N__31110),
            .lcout(\c0.data_in_frame_9_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50474),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_427_LC_6_26_5 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_427_LC_6_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_427_LC_6_26_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_427_LC_6_26_5  (
            .in0(N__26241),
            .in1(N__26832),
            .in2(N__23796),
            .in3(N__23780),
            .lcout(),
            .ltout(\c0.n16954_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_439_LC_6_26_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_439_LC_6_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_439_LC_6_26_6 .LUT_INIT=16'b1111001111111100;
    LogicCell40 \c0.i2_3_lut_adj_439_LC_6_26_6  (
            .in0(_gnd_net_),
            .in1(N__30575),
            .in2(N__23767),
            .in3(N__23691),
            .lcout(),
            .ltout(\c0.n18_adj_2174_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_455_LC_6_26_7 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_455_LC_6_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_455_LC_6_26_7 .LUT_INIT=16'b1111011011111111;
    LogicCell40 \c0.i9_4_lut_adj_455_LC_6_26_7  (
            .in0(N__23763),
            .in1(N__30271),
            .in2(N__23755),
            .in3(N__23752),
            .lcout(\c0.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i77_LC_6_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i77_LC_6_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i77_LC_6_27_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i77_LC_6_27_0  (
            .in0(N__31109),
            .in1(N__28799),
            .in2(N__31826),
            .in3(N__23746),
            .lcout(\c0.data_in_frame_9_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50487),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_421_LC_6_27_1 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_421_LC_6_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_421_LC_6_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_3_lut_adj_421_LC_6_27_1  (
            .in0(N__28392),
            .in1(N__29114),
            .in2(_gnd_net_),
            .in3(N__29049),
            .lcout(\c0.n6_adj_2152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_666_LC_6_27_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_666_LC_6_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_666_LC_6_27_2 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_666_LC_6_27_2  (
            .in0(N__24454),
            .in1(N__24510),
            .in2(N__25144),
            .in3(N__23722),
            .lcout(\c0.n16882 ),
            .ltout(\c0.n16882_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i85_LC_6_27_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i85_LC_6_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i85_LC_6_27_3 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i85_LC_6_27_3  (
            .in0(N__31919),
            .in1(N__31819),
            .in2(N__23695),
            .in3(N__23692),
            .lcout(\c0.data_in_frame_10_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50487),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_429_LC_6_27_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_429_LC_6_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_429_LC_6_27_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_429_LC_6_27_4  (
            .in0(N__23679),
            .in1(N__26242),
            .in2(_gnd_net_),
            .in3(N__28575),
            .lcout(\c0.n15938 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i73_LC_6_27_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i73_LC_6_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i73_LC_6_27_5 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i73_LC_6_27_5  (
            .in0(N__28796),
            .in1(N__28992),
            .in2(N__25595),
            .in3(N__31107),
            .lcout(\c0.data_in_frame_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50487),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i10_LC_6_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i10_LC_6_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i10_LC_6_27_6 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0__i10_LC_6_27_6  (
            .in0(N__29115),
            .in1(N__28798),
            .in2(N__30693),
            .in3(N__31992),
            .lcout(\c0.data_in_frame_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50487),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i76_LC_6_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i76_LC_6_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i76_LC_6_27_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i76_LC_6_27_7  (
            .in0(N__28797),
            .in1(N__28356),
            .in2(N__30531),
            .in3(N__31108),
            .lcout(\c0.data_in_frame_9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50487),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i15_LC_6_28_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i15_LC_6_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i15_LC_6_28_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i15_LC_6_28_0  (
            .in0(N__28800),
            .in1(N__25649),
            .in2(N__26833),
            .in3(N__31998),
            .lcout(\c0.data_in_frame_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50497),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_4_lut_adj_566_LC_6_28_1 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_adj_566_LC_6_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_adj_566_LC_6_28_1 .LUT_INIT=16'b1101011101111101;
    LogicCell40 \c0.i6_3_lut_4_lut_adj_566_LC_6_28_1  (
            .in0(N__26820),
            .in1(N__29036),
            .in2(N__23812),
            .in3(N__30300),
            .lcout(\c0.n22_adj_2301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i88_LC_6_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i88_LC_6_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i88_LC_6_28_2 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i88_LC_6_28_2  (
            .in0(N__31923),
            .in1(N__28467),
            .in2(N__26538),
            .in3(N__31114),
            .lcout(\c0.data_in_frame_10_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50497),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i20_LC_6_28_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i20_LC_6_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i20_LC_6_28_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i20_LC_6_28_3  (
            .in0(N__32000),
            .in1(N__31921),
            .in2(N__30532),
            .in3(N__26271),
            .lcout(\c0.data_in_frame_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50497),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i49_LC_6_28_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i49_LC_6_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i49_LC_6_28_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i49_LC_6_28_4  (
            .in0(N__28872),
            .in1(N__25563),
            .in2(_gnd_net_),
            .in3(N__25735),
            .lcout(data_in_frame_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50497),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i23_LC_6_28_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i23_LC_6_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i23_LC_6_28_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i23_LC_6_28_5  (
            .in0(N__32001),
            .in1(N__31922),
            .in2(N__25665),
            .in3(N__30237),
            .lcout(\c0.data_in_frame_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50497),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i19_LC_6_28_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i19_LC_6_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i19_LC_6_28_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i19_LC_6_28_7  (
            .in0(N__31999),
            .in1(N__31920),
            .in2(N__26940),
            .in3(N__26349),
            .lcout(\c0.data_in_frame_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50497),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i7_LC_6_29_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i7_LC_6_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i7_LC_6_29_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i7_LC_6_29_0  (
            .in0(N__25664),
            .in1(N__29045),
            .in2(_gnd_net_),
            .in3(N__30441),
            .lcout(data_in_frame_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50509),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_LC_6_29_1 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_LC_6_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_LC_6_29_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.tx.i1_2_lut_LC_6_29_1  (
            .in0(_gnd_net_),
            .in1(N__23824),
            .in2(_gnd_net_),
            .in3(N__31642),
            .lcout(\c0.n65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i43_4_lut_LC_6_29_2 .C_ON=1'b0;
    defparam \c0.i43_4_lut_LC_6_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i43_4_lut_LC_6_29_2 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \c0.i43_4_lut_LC_6_29_2  (
            .in0(N__46395),
            .in1(N__26755),
            .in2(N__42749),
            .in3(N__24301),
            .lcout(\c0.n25_adj_2324 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i15400_3_lut_4_lut_4_lut_LC_6_29_3 .C_ON=1'b0;
    defparam \c0.tx.i15400_3_lut_4_lut_4_lut_LC_6_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i15400_3_lut_4_lut_4_lut_LC_6_29_3 .LUT_INIT=16'b1000010110000000;
    LogicCell40 \c0.tx.i15400_3_lut_4_lut_4_lut_LC_6_29_3  (
            .in0(N__24182),
            .in1(N__24113),
            .in2(N__24075),
            .in3(N__31736),
            .lcout(),
            .ltout(n4_adj_2458_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_47_LC_6_29_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_47_LC_6_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Active_47_LC_6_29_4 .LUT_INIT=16'b1010101000111010;
    LogicCell40 \c0.tx.r_Tx_Active_47_LC_6_29_4  (
            .in0(N__31643),
            .in1(N__24074),
            .in2(N__24190),
            .in3(N__23878),
            .lcout(tx_active),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50509),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i2_LC_6_29_5 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i2_LC_6_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i2_LC_6_29_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.tx.r_SM_Main_i2_LC_6_29_5  (
            .in0(N__24183),
            .in1(N__24114),
            .in2(N__24076),
            .in3(N__23877),
            .lcout(r_SM_Main_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50509),
            .ce(),
            .sr(_gnd_net_));
    defparam i14957_3_lut_LC_6_29_6.C_ON=1'b0;
    defparam i14957_3_lut_LC_6_29_6.SEQ_MODE=4'b0000;
    defparam i14957_3_lut_LC_6_29_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 i14957_3_lut_LC_6_29_6 (
            .in0(N__26745),
            .in1(N__32083),
            .in2(_gnd_net_),
            .in3(N__31378),
            .lcout(n17395),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_active_prev_2155_LC_6_29_7 .C_ON=1'b0;
    defparam \c0.tx_active_prev_2155_LC_6_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx_active_prev_2155_LC_6_29_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.tx_active_prev_2155_LC_6_29_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31644),
            .lcout(\c0.tx_active_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50509),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2494_2_lut_LC_6_30_0 .C_ON=1'b1;
    defparam \c0.add_2494_2_lut_LC_6_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_2494_2_lut_LC_6_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2494_2_lut_LC_6_30_0  (
            .in0(_gnd_net_),
            .in1(N__23818),
            .in2(N__51887),
            .in3(_gnd_net_),
            .lcout(\c0.tx_transmit_N_1949_0 ),
            .ltout(),
            .carryin(bfn_6_30_0_),
            .carryout(\c0.n15653 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2494_3_lut_LC_6_30_1 .C_ON=1'b1;
    defparam \c0.add_2494_3_lut_LC_6_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_2494_3_lut_LC_6_30_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2494_3_lut_LC_6_30_1  (
            .in0(_gnd_net_),
            .in1(N__52175),
            .in2(_gnd_net_),
            .in3(N__24217),
            .lcout(\c0.tx_transmit_N_1949_1 ),
            .ltout(),
            .carryin(\c0.n15653 ),
            .carryout(\c0.n15654 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2494_4_lut_LC_6_30_2 .C_ON=1'b1;
    defparam \c0.add_2494_4_lut_LC_6_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_2494_4_lut_LC_6_30_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2494_4_lut_LC_6_30_2  (
            .in0(_gnd_net_),
            .in1(N__52351),
            .in2(_gnd_net_),
            .in3(N__24214),
            .lcout(\c0.tx_transmit_N_1949_2 ),
            .ltout(),
            .carryin(\c0.n15654 ),
            .carryout(\c0.n15655 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2494_5_lut_LC_6_30_3 .C_ON=1'b1;
    defparam \c0.add_2494_5_lut_LC_6_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_2494_5_lut_LC_6_30_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2494_5_lut_LC_6_30_3  (
            .in0(_gnd_net_),
            .in1(N__43078),
            .in2(_gnd_net_),
            .in3(N__24211),
            .lcout(\c0.tx_transmit_N_1949_3 ),
            .ltout(),
            .carryin(\c0.n15655 ),
            .carryout(\c0.n15656 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2494_6_lut_LC_6_30_4 .C_ON=1'b1;
    defparam \c0.add_2494_6_lut_LC_6_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_2494_6_lut_LC_6_30_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2494_6_lut_LC_6_30_4  (
            .in0(_gnd_net_),
            .in1(N__35471),
            .in2(_gnd_net_),
            .in3(N__24208),
            .lcout(\c0.tx_transmit_N_1949_4 ),
            .ltout(),
            .carryin(\c0.n15656 ),
            .carryout(\c0.n15657 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2494_7_lut_LC_6_30_5 .C_ON=1'b1;
    defparam \c0.add_2494_7_lut_LC_6_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_2494_7_lut_LC_6_30_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2494_7_lut_LC_6_30_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26596),
            .in3(N__24205),
            .lcout(\c0.tx_transmit_N_1949_5 ),
            .ltout(),
            .carryin(\c0.n15657 ),
            .carryout(\c0.n15658 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2494_8_lut_LC_6_30_6 .C_ON=1'b1;
    defparam \c0.add_2494_8_lut_LC_6_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_2494_8_lut_LC_6_30_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2494_8_lut_LC_6_30_6  (
            .in0(_gnd_net_),
            .in1(N__27012),
            .in2(_gnd_net_),
            .in3(N__24202),
            .lcout(\c0.tx_transmit_N_1949_6 ),
            .ltout(),
            .carryin(\c0.n15658 ),
            .carryout(\c0.n15659 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2494_9_lut_LC_6_30_7 .C_ON=1'b0;
    defparam \c0.add_2494_9_lut_LC_6_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_2494_9_lut_LC_6_30_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2494_9_lut_LC_6_30_7  (
            .in0(_gnd_net_),
            .in1(N__27105),
            .in2(_gnd_net_),
            .in3(N__24199),
            .lcout(\c0.tx_transmit_N_1949_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i1_LC_6_31_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i1_LC_6_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i1_LC_6_31_1 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.byte_transmit_counter__i1_LC_6_31_1  (
            .in0(N__24238),
            .in1(N__35745),
            .in2(N__52236),
            .in3(N__27145),
            .lcout(\c0.byte_transmit_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50526),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i152_2_lut_4_lut_LC_6_31_2 .C_ON=1'b0;
    defparam \c0.i152_2_lut_4_lut_LC_6_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.i152_2_lut_4_lut_LC_6_31_2 .LUT_INIT=16'b1111111111110001;
    LogicCell40 \c0.i152_2_lut_4_lut_LC_6_31_2  (
            .in0(N__27171),
            .in1(N__27189),
            .in2(N__31737),
            .in3(N__31660),
            .lcout(\c0.n456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_LC_6_31_3 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_LC_6_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_LC_6_31_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i3_2_lut_3_lut_LC_6_31_3  (
            .in0(N__26957),
            .in1(N__27026),
            .in2(_gnd_net_),
            .in3(N__27039),
            .lcout(\c0.n8938 ),
            .ltout(\c0.n8938_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_677_LC_6_31_4 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_677_LC_6_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_677_LC_6_31_4 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_677_LC_6_31_4  (
            .in0(N__27170),
            .in1(N__27338),
            .in2(N__24253),
            .in3(N__27308),
            .lcout(\c0.n22_adj_2164 ),
            .ltout(\c0.n22_adj_2164_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_4_lut_LC_6_31_5 .C_ON=1'b0;
    defparam \c0.i1_4_lut_4_lut_LC_6_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_4_lut_LC_6_31_5 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \c0.i1_4_lut_4_lut_LC_6_31_5  (
            .in0(N__42574),
            .in1(N__46415),
            .in2(N__24241),
            .in3(N__27385),
            .lcout(\c0.n42_adj_2165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_604_LC_6_31_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_604_LC_6_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_604_LC_6_31_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.i1_2_lut_adj_604_LC_6_31_6  (
            .in0(N__26973),
            .in1(N__24237),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n4_adj_2311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15441_2_lut_3_lut_LC_6_31_7 .C_ON=1'b0;
    defparam \c0.i15441_2_lut_3_lut_LC_6_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15441_2_lut_3_lut_LC_6_31_7 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \c0.i15441_2_lut_3_lut_LC_6_31_7  (
            .in0(N__42575),
            .in1(_gnd_net_),
            .in2(N__45848),
            .in3(N__46416),
            .lcout(data_out_10__7__N_110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6219_4_lut_LC_6_32_0 .C_ON=1'b0;
    defparam \c0.i6219_4_lut_LC_6_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6219_4_lut_LC_6_32_0 .LUT_INIT=16'b1010111110101100;
    LogicCell40 \c0.i6219_4_lut_LC_6_32_0  (
            .in0(N__24283),
            .in1(N__24300),
            .in2(N__42645),
            .in3(N__45761),
            .lcout(\c0.n8631 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_697_LC_6_32_1 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_697_LC_6_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_697_LC_6_32_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \c0.i2_4_lut_adj_697_LC_6_32_1  (
            .in0(N__46302),
            .in1(N__34309),
            .in2(N__45549),
            .in3(N__27427),
            .lcout(),
            .ltout(\c0.n15868_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_701_LC_6_32_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_701_LC_6_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_701_LC_6_32_2 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \c0.i1_4_lut_adj_701_LC_6_32_2  (
            .in0(N__27576),
            .in1(N__46303),
            .in2(N__24229),
            .in3(N__24226),
            .lcout(),
            .ltout(n10141_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.UART_TRANSMITTER_state_i0_i1_LC_6_32_3 .C_ON=1'b0;
    defparam \c0.UART_TRANSMITTER_state_i0_i1_LC_6_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.UART_TRANSMITTER_state_i0_i1_LC_6_32_3 .LUT_INIT=16'b0101101000001010;
    LogicCell40 \c0.UART_TRANSMITTER_state_i0_i1_LC_6_32_3  (
            .in0(N__46304),
            .in1(_gnd_net_),
            .in2(N__24220),
            .in3(N__45907),
            .lcout(UART_TRANSMITTER_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50537),
            .ce(),
            .sr(_gnd_net_));
    defparam i14724_2_lut_LC_6_32_4.C_ON=1'b0;
    defparam i14724_2_lut_LC_6_32_4.SEQ_MODE=4'b0000;
    defparam i14724_2_lut_LC_6_32_4.LUT_INIT=16'b1111111110101010;
    LogicCell40 i14724_2_lut_LC_6_32_4 (
            .in0(N__34310),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46301),
            .lcout(n17162),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__6__2214_LC_6_32_5 .C_ON=1'b0;
    defparam \c0.data_out_3__6__2214_LC_6_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__6__2214_LC_6_32_5 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \c0.data_out_3__6__2214_LC_6_32_5  (
            .in0(N__46305),
            .in1(N__34053),
            .in2(N__46150),
            .in3(N__42580),
            .lcout(\c0.data_out_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50537),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i142_2_lut_4_lut_LC_6_32_6 .C_ON=1'b0;
    defparam \c0.i142_2_lut_4_lut_LC_6_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.i142_2_lut_4_lut_LC_6_32_6 .LUT_INIT=16'b1111000011110111;
    LogicCell40 \c0.i142_2_lut_4_lut_LC_6_32_6  (
            .in0(N__27357),
            .in1(N__27310),
            .in2(N__27464),
            .in3(N__27375),
            .lcout(\c0.n446 ),
            .ltout(\c0.n446_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15401_4_lut_LC_6_32_7 .C_ON=1'b0;
    defparam \c0.i15401_4_lut_LC_6_32_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15401_4_lut_LC_6_32_7 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \c0.i15401_4_lut_LC_6_32_7  (
            .in0(N__45760),
            .in1(N__42576),
            .in2(N__24286),
            .in3(N__24282),
            .lcout(n10031),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i19_LC_7_15_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i19_LC_7_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i19_LC_7_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i19_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__24602),
            .in2(_gnd_net_),
            .in3(N__34654),
            .lcout(\c0.FRAME_MATCHER_state_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50420),
            .ce(),
            .sr(N__24274));
    defparam \c0.FRAME_MATCHER_state_i10_LC_7_17_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i10_LC_7_17_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i10_LC_7_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i10_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__25260),
            .in2(_gnd_net_),
            .in3(N__34644),
            .lcout(\c0.FRAME_MATCHER_state_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50399),
            .ce(),
            .sr(N__24262));
    defparam \c0.FRAME_MATCHER_state_i21_LC_7_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i21_LC_7_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i21_LC_7_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i21_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(N__25412),
            .in2(_gnd_net_),
            .in3(N__34562),
            .lcout(\c0.FRAME_MATCHER_state_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50411),
            .ce(),
            .sr(N__25387));
    defparam \c0.FRAME_MATCHER_state_i22_LC_7_19_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i22_LC_7_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i22_LC_7_19_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i22_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__25515),
            .in2(_gnd_net_),
            .in3(N__34560),
            .lcout(\c0.FRAME_MATCHER_state_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50421),
            .ce(),
            .sr(N__25498));
    defparam \c0.i4_4_lut_adj_649_LC_7_19_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_649_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_649_LC_7_19_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i4_4_lut_adj_649_LC_7_19_1  (
            .in0(N__28141),
            .in1(N__25374),
            .in2(N__29536),
            .in3(N__24604),
            .lcout(\c0.n10_adj_2336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_466_LC_7_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_466_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_466_LC_7_19_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i1_2_lut_adj_466_LC_7_19_2  (
            .in0(N__25408),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25514),
            .lcout(),
            .ltout(\c0.n61_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_443_LC_7_19_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_443_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_443_LC_7_19_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_443_LC_7_19_3  (
            .in0(N__24637),
            .in1(N__27991),
            .in2(N__24628),
            .in3(N__27880),
            .lcout(),
            .ltout(\c0.n16133_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_650_LC_7_19_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_650_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_650_LC_7_19_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_4_lut_adj_650_LC_7_19_4  (
            .in0(N__24625),
            .in1(N__32403),
            .in2(N__24619),
            .in3(N__24616),
            .lcout(\c0.n62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_695_LC_7_19_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_695_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_695_LC_7_19_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_695_LC_7_19_6  (
            .in0(N__24603),
            .in1(N__25513),
            .in2(N__25413),
            .in3(N__29809),
            .lcout(\c0.n52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_732_LC_7_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_732_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_732_LC_7_19_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_732_LC_7_19_7  (
            .in0(N__32404),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29945),
            .lcout(\c0.n16347 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i26_LC_7_20_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i26_LC_7_20_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i26_LC_7_20_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i26_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__25373),
            .in2(_gnd_net_),
            .in3(N__34563),
            .lcout(\c0.FRAME_MATCHER_state_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50427),
            .ce(),
            .sr(N__25345));
    defparam \c0.FRAME_MATCHER_i_i4_LC_7_21_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i4_LC_7_21_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i4_LC_7_21_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i4_LC_7_21_0  (
            .in0(N__33247),
            .in1(N__32802),
            .in2(_gnd_net_),
            .in3(N__24574),
            .lcout(\c0.FRAME_MATCHER_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50435),
            .ce(),
            .sr(N__24562));
    defparam \c0.i1_2_lut_adj_408_LC_7_21_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_408_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_408_LC_7_21_1 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \c0.i1_2_lut_adj_408_LC_7_21_1  (
            .in0(N__24535),
            .in1(N__24475),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_LC_7_21_2 .C_ON=1'b0;
    defparam \c0.i22_4_lut_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_LC_7_21_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i22_4_lut_LC_7_21_2  (
            .in0(N__24446),
            .in1(N__24398),
            .in2(N__24352),
            .in3(N__24348),
            .lcout(\c0.n51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_441_LC_7_21_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_441_LC_7_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_441_LC_7_21_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_441_LC_7_21_3  (
            .in0(N__27983),
            .in1(N__27879),
            .in2(N__30064),
            .in3(N__25231),
            .lcout(\c0.n56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_468_LC_7_21_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_468_LC_7_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_468_LC_7_21_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i4_4_lut_adj_468_LC_7_21_4  (
            .in0(N__25261),
            .in1(N__32614),
            .in2(N__34441),
            .in3(N__25240),
            .lcout(\c0.n16869 ),
            .ltout(\c0.n16869_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_471_LC_7_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_471_LC_7_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_471_LC_7_21_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \c0.i1_2_lut_adj_471_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25225),
            .in3(N__30028),
            .lcout(\c0.n16871 ),
            .ltout(\c0.n16871_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_496_LC_7_21_6 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_496_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_496_LC_7_21_6 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i5_4_lut_adj_496_LC_7_21_6  (
            .in0(N__29532),
            .in1(N__32310),
            .in2(N__25222),
            .in3(N__25219),
            .lcout(\c0.n12_adj_2189 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i27_4_lut_LC_7_22_0 .C_ON=1'b0;
    defparam \c0.i27_4_lut_LC_7_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i27_4_lut_LC_7_22_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i27_4_lut_LC_7_22_0  (
            .in0(N__28213),
            .in1(N__24643),
            .in2(N__25213),
            .in3(N__24778),
            .lcout(),
            .ltout(\c0.n56_adj_2146_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i28_4_lut_LC_7_22_1 .C_ON=1'b0;
    defparam \c0.i28_4_lut_LC_7_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i28_4_lut_LC_7_22_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i28_4_lut_LC_7_22_1  (
            .in0(N__24967),
            .in1(N__25204),
            .in2(N__25189),
            .in3(N__25186),
            .lcout(\c0.n9346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_LC_7_22_2 .C_ON=1'b0;
    defparam \c0.i16_4_lut_LC_7_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_LC_7_22_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i16_4_lut_LC_7_22_2  (
            .in0(N__25121),
            .in1(N__25087),
            .in2(N__25016),
            .in3(N__25451),
            .lcout(\c0.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_407_LC_7_22_3 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_407_LC_7_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_407_LC_7_22_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i18_4_lut_adj_407_LC_7_22_3  (
            .in0(N__24956),
            .in1(N__24909),
            .in2(N__24864),
            .in3(N__24808),
            .lcout(\c0.n47_adj_2144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_LC_7_22_4 .C_ON=1'b0;
    defparam \c0.i20_4_lut_LC_7_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_LC_7_22_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i20_4_lut_LC_7_22_4  (
            .in0(N__24751),
            .in1(N__24712),
            .in2(N__28084),
            .in3(N__24681),
            .lcout(\c0.n49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_744_LC_7_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_744_LC_7_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_744_LC_7_22_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_744_LC_7_22_5  (
            .in0(_gnd_net_),
            .in1(N__25519),
            .in2(_gnd_net_),
            .in3(N__29894),
            .lcout(\c0.n16365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i12_LC_7_23_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i12_LC_7_23_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i12_LC_7_23_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i12_LC_7_23_0  (
            .in0(N__33209),
            .in1(N__32847),
            .in2(_gnd_net_),
            .in3(N__25486),
            .lcout(\c0.FRAME_MATCHER_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50453),
            .ce(),
            .sr(N__25438));
    defparam \c0.i1_2_lut_adj_728_LC_7_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_728_LC_7_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_728_LC_7_23_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_728_LC_7_23_1  (
            .in0(_gnd_net_),
            .in1(N__29824),
            .in2(_gnd_net_),
            .in3(N__29884),
            .lcout(\c0.n16351 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_742_LC_7_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_742_LC_7_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_742_LC_7_23_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_742_LC_7_23_3  (
            .in0(_gnd_net_),
            .in1(N__25414),
            .in2(_gnd_net_),
            .in3(N__29885),
            .lcout(\c0.n16367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_752_LC_7_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_752_LC_7_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_752_LC_7_23_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.i1_2_lut_adj_752_LC_7_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29917),
            .in3(N__28139),
            .lcout(\c0.n16359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_754_LC_7_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_754_LC_7_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_754_LC_7_23_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_754_LC_7_23_5  (
            .in0(_gnd_net_),
            .in1(N__25375),
            .in2(_gnd_net_),
            .in3(N__29889),
            .lcout(\c0.n16357 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_756_LC_7_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_756_LC_7_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_756_LC_7_23_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.i1_2_lut_adj_756_LC_7_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29918),
            .in3(N__25333),
            .lcout(\c0.n16355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14828_4_lut_LC_7_24_1 .C_ON=1'b0;
    defparam \c0.i14828_4_lut_LC_7_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14828_4_lut_LC_7_24_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i14828_4_lut_LC_7_24_1  (
            .in0(N__25293),
            .in1(N__26176),
            .in2(N__25886),
            .in3(N__25850),
            .lcout(\c0.n17266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i50_LC_7_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i50_LC_7_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i50_LC_7_24_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i50_LC_7_24_2  (
            .in0(N__30696),
            .in1(N__26035),
            .in2(_gnd_net_),
            .in3(N__25724),
            .lcout(data_in_frame_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50463),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__5__2260_LC_7_24_3 .C_ON=1'b0;
    defparam \c0.data_in_2__5__2260_LC_7_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__5__2260_LC_7_24_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_2__5__2260_LC_7_24_3  (
            .in0(N__25879),
            .in1(N__27803),
            .in2(_gnd_net_),
            .in3(N__25930),
            .lcout(data_in_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50463),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__7__2258_LC_7_24_4 .C_ON=1'b0;
    defparam \c0.data_in_2__7__2258_LC_7_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__7__2258_LC_7_24_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_2__7__2258_LC_7_24_4  (
            .in0(N__25851),
            .in1(_gnd_net_),
            .in2(N__27808),
            .in3(N__25818),
            .lcout(data_in_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50463),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_432_LC_7_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_432_LC_7_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_432_LC_7_24_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_432_LC_7_24_5  (
            .in0(_gnd_net_),
            .in1(N__25790),
            .in2(_gnd_net_),
            .in3(N__27824),
            .lcout(\c0.n8_adj_2157 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__7__2250_LC_7_24_6 .C_ON=1'b0;
    defparam \c0.data_in_3__7__2250_LC_7_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__7__2250_LC_7_24_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_3__7__2250_LC_7_24_6  (
            .in0(N__27802),
            .in1(N__26520),
            .in2(_gnd_net_),
            .in3(N__25817),
            .lcout(data_in_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50463),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__3__2254_LC_7_24_7 .C_ON=1'b0;
    defparam \c0.data_in_3__3__2254_LC_7_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__3__2254_LC_7_24_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_3__3__2254_LC_7_24_7  (
            .in0(N__25794),
            .in1(N__27804),
            .in2(_gnd_net_),
            .in3(N__30488),
            .lcout(data_in_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50463),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_412_LC_7_25_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_412_LC_7_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_412_LC_7_25_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \c0.i1_4_lut_adj_412_LC_7_25_0  (
            .in0(N__30267),
            .in1(N__25774),
            .in2(N__25756),
            .in3(N__30191),
            .lcout(\c0.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1028_2_lut_LC_7_25_1 .C_ON=1'b0;
    defparam \c0.i1028_2_lut_LC_7_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1028_2_lut_LC_7_25_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1028_2_lut_LC_7_25_1  (
            .in0(N__30377),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25950),
            .lcout(\c0.n2334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i55_LC_7_25_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i55_LC_7_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i55_LC_7_25_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i55_LC_7_25_2  (
            .in0(N__25731),
            .in1(N__25673),
            .in2(_gnd_net_),
            .in3(N__26091),
            .lcout(data_in_frame_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50475),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i1_LC_7_25_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i1_LC_7_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i1_LC_7_25_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i1_LC_7_25_3  (
            .in0(N__26852),
            .in1(N__25603),
            .in2(_gnd_net_),
            .in3(N__30436),
            .lcout(data_in_frame_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50475),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i2_LC_7_25_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i2_LC_7_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i2_LC_7_25_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i2_LC_7_25_4  (
            .in0(N__30437),
            .in1(N__30695),
            .in2(_gnd_net_),
            .in3(N__26780),
            .lcout(data_in_frame_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50475),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_746_LC_7_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_746_LC_7_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_746_LC_7_25_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_746_LC_7_25_5  (
            .in0(N__29055),
            .in1(N__28649),
            .in2(_gnd_net_),
            .in3(N__25962),
            .lcout(\c0.n2351 ),
            .ltout(\c0.n2351_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1046_2_lut_LC_7_25_6 .C_ON=1'b0;
    defparam \c0.i1046_2_lut_LC_7_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1046_2_lut_LC_7_25_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1046_2_lut_LC_7_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26056),
            .in3(N__26851),
            .lcout(\c0.n2352 ),
            .ltout(\c0.n2352_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_LC_7_25_7 .C_ON=1'b0;
    defparam \c0.i7_4_lut_LC_7_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_LC_7_25_7 .LUT_INIT=16'b1011011111101101;
    LogicCell40 \c0.i7_4_lut_LC_7_25_7  (
            .in0(N__26053),
            .in1(N__26034),
            .in2(N__26023),
            .in3(N__28650),
            .lcout(\c0.n23_adj_2145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_LC_7_26_0 .C_ON=1'b0;
    defparam \c0.i14_4_lut_LC_7_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_LC_7_26_0 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \c0.i14_4_lut_LC_7_26_0  (
            .in0(N__26020),
            .in1(N__26545),
            .in2(N__26002),
            .in3(N__25978),
            .lcout(\c0.n30_adj_2148 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i137_LC_7_26_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i137_LC_7_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i137_LC_7_26_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i137_LC_7_26_1  (
            .in0(N__48769),
            .in1(N__34785),
            .in2(_gnd_net_),
            .in3(N__51249),
            .lcout(data_out_frame2_17_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50488),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_416_LC_7_26_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_416_LC_7_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_416_LC_7_26_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_416_LC_7_26_2  (
            .in0(_gnd_net_),
            .in1(N__25948),
            .in2(_gnd_net_),
            .in3(N__26773),
            .lcout(\c0.n9541 ),
            .ltout(\c0.n9541_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_414_LC_7_26_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_414_LC_7_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_414_LC_7_26_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_414_LC_7_26_3  (
            .in0(N__30334),
            .in1(N__30378),
            .in2(N__25972),
            .in3(N__30299),
            .lcout(\c0.n16943 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_715_LC_7_26_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_715_LC_7_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_715_LC_7_26_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_715_LC_7_26_4  (
            .in0(N__28610),
            .in1(N__25949),
            .in2(N__26109),
            .in3(N__26774),
            .lcout(\c0.n15929 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1030_2_lut_LC_7_26_5 .C_ON=1'b0;
    defparam \c0.i1030_2_lut_LC_7_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1030_2_lut_LC_7_26_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1030_2_lut_LC_7_26_5  (
            .in0(N__30335),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30379),
            .lcout(\c0.n2336 ),
            .ltout(\c0.n2336_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_655_LC_7_26_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_655_LC_7_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_655_LC_7_26_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \c0.i4_4_lut_adj_655_LC_7_26_6  (
            .in0(N__26287),
            .in1(N__26272),
            .in2(N__26257),
            .in3(N__28887),
            .lcout(),
            .ltout(\c0.n20_adj_2340_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_659_LC_7_26_7 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_659_LC_7_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_659_LC_7_26_7 .LUT_INIT=16'b1111110111110111;
    LogicCell40 \c0.i10_4_lut_adj_659_LC_7_26_7  (
            .in0(N__26254),
            .in1(N__28827),
            .in2(N__26215),
            .in3(N__26435),
            .lcout(\c0.n26_adj_2344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15345_2_lut_LC_7_27_0 .C_ON=1'b0;
    defparam \c0.i15345_2_lut_LC_7_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15345_2_lut_LC_7_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15345_2_lut_LC_7_27_0  (
            .in0(_gnd_net_),
            .in1(N__40243),
            .in2(_gnd_net_),
            .in3(N__51938),
            .lcout(\c0.n17548 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1036_2_lut_LC_7_27_1 .C_ON=1'b0;
    defparam \c0.i1036_2_lut_LC_7_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1036_2_lut_LC_7_27_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1036_2_lut_LC_7_27_1  (
            .in0(_gnd_net_),
            .in1(N__28645),
            .in2(_gnd_net_),
            .in3(N__29050),
            .lcout(\c0.n2342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__2__2263_LC_7_27_2 .C_ON=1'b0;
    defparam \c0.data_in_2__2__2263_LC_7_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__2__2263_LC_7_27_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_2__2__2263_LC_7_27_2  (
            .in0(N__26174),
            .in1(N__27742),
            .in2(_gnd_net_),
            .in3(N__26212),
            .lcout(data_in_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50498),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__2__2271_LC_7_27_3 .C_ON=1'b0;
    defparam \c0.data_in_1__2__2271_LC_7_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__2__2271_LC_7_27_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_1__2__2271_LC_7_27_3  (
            .in0(N__27741),
            .in1(N__26131),
            .in2(_gnd_net_),
            .in3(N__26175),
            .lcout(data_in_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50498),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i84_LC_7_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i84_LC_7_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i84_LC_7_27_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i84_LC_7_27_4  (
            .in0(N__31925),
            .in1(N__30512),
            .in2(N__26110),
            .in3(N__31113),
            .lcout(\c0.data_in_frame_10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50498),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_4_lut_adj_716_LC_7_27_5 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_adj_716_LC_7_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_adj_716_LC_7_27_5 .LUT_INIT=16'b1101011101111101;
    LogicCell40 \c0.i6_3_lut_4_lut_adj_716_LC_7_27_5  (
            .in0(N__26092),
            .in1(N__29051),
            .in2(N__26077),
            .in3(N__30304),
            .lcout(),
            .ltout(\c0.n22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_LC_7_27_6 .C_ON=1'b0;
    defparam \c0.i11_4_lut_LC_7_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_LC_7_27_6 .LUT_INIT=16'b1111011111111011;
    LogicCell40 \c0.i11_4_lut_LC_7_27_6  (
            .in0(N__26581),
            .in1(N__26563),
            .in2(N__26548),
            .in3(N__26356),
            .lcout(\c0.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i6_LC_7_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i6_LC_7_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i6_LC_7_27_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i6_LC_7_27_7  (
            .in0(N__31221),
            .in1(N__30305),
            .in2(_gnd_net_),
            .in3(N__30434),
            .lcout(data_in_frame_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50498),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i8_LC_7_28_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i8_LC_7_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i8_LC_7_28_0 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.data_in_frame_0__i8_LC_7_28_0  (
            .in0(N__28644),
            .in1(_gnd_net_),
            .in2(N__26536),
            .in3(N__30435),
            .lcout(data_in_frame_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50510),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_413_LC_7_28_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_413_LC_7_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_413_LC_7_28_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_413_LC_7_28_1  (
            .in0(_gnd_net_),
            .in1(N__26437),
            .in2(_gnd_net_),
            .in3(N__28643),
            .lcout(\c0.n17001 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i6_LC_7_28_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i6_LC_7_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i6_LC_7_28_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i6_LC_7_28_2  (
            .in0(N__26378),
            .in1(N__31550),
            .in2(_gnd_net_),
            .in3(N__26401),
            .lcout(r_Clock_Count_6_adj_2448),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50510),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_417_LC_7_28_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_417_LC_7_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_417_LC_7_28_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_417_LC_7_28_3  (
            .in0(N__26859),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26781),
            .lcout(\c0.n9585 ),
            .ltout(\c0.n9585_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_657_LC_7_28_4 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_657_LC_7_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_657_LC_7_28_4 .LUT_INIT=16'b1101111011111111;
    LogicCell40 \c0.i11_4_lut_adj_657_LC_7_28_4  (
            .in0(N__26350),
            .in1(N__26335),
            .in2(N__26329),
            .in3(N__28398),
            .lcout(\c0.n27_adj_2342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_LC_7_28_5 .C_ON=1'b0;
    defparam \c0.i2_4_lut_LC_7_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_LC_7_28_5 .LUT_INIT=16'b1011111001111101;
    LogicCell40 \c0.i2_4_lut_LC_7_28_5  (
            .in0(N__26326),
            .in1(N__30580),
            .in2(N__26308),
            .in3(N__30556),
            .lcout(\c0.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i83_LC_7_28_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i83_LC_7_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i83_LC_7_28_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i83_LC_7_28_6  (
            .in0(N__31115),
            .in1(N__31933),
            .in2(N__26941),
            .in3(N__26793),
            .lcout(\c0.data_in_frame_10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50510),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_702_LC_7_28_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_702_LC_7_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_702_LC_7_28_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_702_LC_7_28_7  (
            .in0(N__26860),
            .in1(N__26824),
            .in2(N__26794),
            .in3(N__26782),
            .lcout(\c0.n15930 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15216_3_lut_LC_7_29_0 .C_ON=1'b0;
    defparam \c0.i15216_3_lut_LC_7_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15216_3_lut_LC_7_29_0 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \c0.i15216_3_lut_LC_7_29_0  (
            .in0(N__27471),
            .in1(N__27073),
            .in2(_gnd_net_),
            .in3(N__27193),
            .lcout(\c0.n17460 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i3_LC_7_29_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i3_LC_7_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i3_LC_7_29_2 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \c0.tx.r_Tx_Data_i3_LC_7_29_2  (
            .in0(N__26749),
            .in1(N__43039),
            .in2(N__35617),
            .in3(N__35511),
            .lcout(r_Tx_Data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50518),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14798_2_lut_LC_7_29_3 .C_ON=1'b0;
    defparam \c0.i14798_2_lut_LC_7_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14798_2_lut_LC_7_29_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i14798_2_lut_LC_7_29_3  (
            .in0(N__26733),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26704),
            .lcout(\c0.n17236 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_2_lut_LC_7_29_4 .C_ON=1'b0;
    defparam \c0.i21_2_lut_LC_7_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i21_2_lut_LC_7_29_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i21_2_lut_LC_7_29_4  (
            .in0(_gnd_net_),
            .in1(N__38106),
            .in2(_gnd_net_),
            .in3(N__42403),
            .lcout(\c0.n9530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i150_LC_7_29_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i150_LC_7_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i150_LC_7_29_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i150_LC_7_29_5  (
            .in0(N__41470),
            .in1(N__30897),
            .in2(_gnd_net_),
            .in3(N__51271),
            .lcout(data_out_frame2_18_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50518),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_581_LC_7_30_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_581_LC_7_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_581_LC_7_30_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \c0.i10_4_lut_adj_581_LC_7_30_0  (
            .in0(N__26674),
            .in1(N__26645),
            .in2(N__26614),
            .in3(N__26602),
            .lcout(\c0.n23_adj_2309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i5_LC_7_30_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i5_LC_7_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i5_LC_7_30_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \c0.byte_transmit_counter__i5_LC_7_30_1  (
            .in0(N__27147),
            .in1(N__35763),
            .in2(N__27052),
            .in3(N__26595),
            .lcout(\c0.byte_transmit_counter_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50527),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14816_3_lut_4_lut_LC_7_30_2 .C_ON=1'b0;
    defparam \c0.i14816_3_lut_4_lut_LC_7_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14816_3_lut_4_lut_LC_7_30_2 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.i14816_3_lut_4_lut_LC_7_30_2  (
            .in0(N__27309),
            .in1(N__27347),
            .in2(N__46399),
            .in3(N__27172),
            .lcout(\c0.n17254 ),
            .ltout(\c0.n17254_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14852_3_lut_4_lut_LC_7_30_3 .C_ON=1'b0;
    defparam \c0.i14852_3_lut_4_lut_LC_7_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14852_3_lut_4_lut_LC_7_30_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14852_3_lut_4_lut_LC_7_30_3  (
            .in0(N__26958),
            .in1(N__27027),
            .in2(N__27067),
            .in3(N__27040),
            .lcout(\c0.n17290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i2_LC_7_30_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i2_LC_7_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i2_LC_7_30_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter__i2_LC_7_30_4  (
            .in0(N__35762),
            .in1(N__27348),
            .in2(N__52437),
            .in3(N__27146),
            .lcout(byte_transmit_counter_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50527),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_610_LC_7_30_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_610_LC_7_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_610_LC_7_30_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i1_2_lut_adj_610_LC_7_30_5  (
            .in0(N__27048),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27117),
            .lcout(\c0.n5_adj_2319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i6_LC_7_30_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i6_LC_7_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i6_LC_7_30_6 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \c0.byte_transmit_counter__i6_LC_7_30_6  (
            .in0(N__27028),
            .in1(N__27013),
            .in2(N__35772),
            .in3(N__27148),
            .lcout(\c0.byte_transmit_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50527),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__6__2238_LC_7_30_7 .C_ON=1'b0;
    defparam \c0.data_out_0__6__2238_LC_7_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__6__2238_LC_7_30_7 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \c0.data_out_0__6__2238_LC_7_30_7  (
            .in0(N__32055),
            .in1(N__42644),
            .in2(N__46149),
            .in3(N__46321),
            .lcout(\c0.data_out_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50527),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_582_LC_7_31_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_582_LC_7_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_582_LC_7_31_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.i1_4_lut_adj_582_LC_7_31_0  (
            .in0(N__27001),
            .in1(N__26995),
            .in2(N__31608),
            .in3(N__26986),
            .lcout(\c0.n16839 ),
            .ltout(\c0.n16839_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i0_LC_7_31_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i0_LC_7_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i0_LC_7_31_1 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \c0.byte_transmit_counter__i0_LC_7_31_1  (
            .in0(N__35767),
            .in1(N__26974),
            .in2(N__26962),
            .in3(N__51972),
            .lcout(\c0.byte_transmit_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50538),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i4_LC_7_31_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i4_LC_7_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i4_LC_7_31_2 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \c0.byte_transmit_counter__i4_LC_7_31_2  (
            .in0(N__35490),
            .in1(N__26959),
            .in2(N__35760),
            .in3(N__27143),
            .lcout(byte_transmit_counter_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50538),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11084_2_lut_LC_7_31_3 .C_ON=1'b0;
    defparam \c0.i11084_2_lut_LC_7_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11084_2_lut_LC_7_31_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i11084_2_lut_LC_7_31_3  (
            .in0(_gnd_net_),
            .in1(N__27168),
            .in2(_gnd_net_),
            .in3(N__27188),
            .lcout(n9357),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i3_LC_7_31_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i3_LC_7_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i3_LC_7_31_4 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.byte_transmit_counter__i3_LC_7_31_4  (
            .in0(N__27169),
            .in1(N__35768),
            .in2(N__43139),
            .in3(N__27142),
            .lcout(byte_transmit_counter_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50538),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i7_LC_7_31_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i7_LC_7_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i7_LC_7_31_5 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \c0.byte_transmit_counter__i7_LC_7_31_5  (
            .in0(N__27144),
            .in1(N__27106),
            .in2(N__35773),
            .in3(N__27118),
            .lcout(\c0.byte_transmit_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50538),
            .ce(),
            .sr(_gnd_net_));
    defparam i15393_3_lut_4_lut_LC_7_31_6.C_ON=1'b0;
    defparam i15393_3_lut_4_lut_LC_7_31_6.SEQ_MODE=4'b0000;
    defparam i15393_3_lut_4_lut_LC_7_31_6.LUT_INIT=16'b1010101010000000;
    LogicCell40 i15393_3_lut_4_lut_LC_7_31_6 (
            .in0(N__42646),
            .in1(N__46306),
            .in2(N__45928),
            .in3(N__27577),
            .lcout(),
            .ltout(n17834_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.UART_TRANSMITTER_state_i0_i0_LC_7_31_7 .C_ON=1'b0;
    defparam \c0.UART_TRANSMITTER_state_i0_i0_LC_7_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.UART_TRANSMITTER_state_i0_i0_LC_7_31_7 .LUT_INIT=16'b1000100010001101;
    LogicCell40 \c0.UART_TRANSMITTER_state_i0_i0_LC_7_31_7  (
            .in0(N__45844),
            .in1(N__45548),
            .in2(N__27094),
            .in3(N__27091),
            .lcout(UART_TRANSMITTER_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50538),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.UART_TRANSMITTER_state_i0_i2_LC_7_32_0 .C_ON=1'b0;
    defparam \c0.UART_TRANSMITTER_state_i0_i2_LC_7_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.UART_TRANSMITTER_state_i0_i2_LC_7_32_0 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \c0.UART_TRANSMITTER_state_i0_i2_LC_7_32_0  (
            .in0(N__34291),
            .in1(N__27079),
            .in2(N__42623),
            .in3(N__27391),
            .lcout(UART_TRANSMITTER_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50547),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_692_LC_7_32_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_692_LC_7_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_692_LC_7_32_1 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_692_LC_7_32_1  (
            .in0(N__27377),
            .in1(N__27353),
            .in2(_gnd_net_),
            .in3(N__27312),
            .lcout(),
            .ltout(n9358_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_792_LC_7_32_2.C_ON=1'b0;
    defparam i1_4_lut_adj_792_LC_7_32_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_792_LC_7_32_2.LUT_INIT=16'b1111111100100000;
    LogicCell40 i1_4_lut_adj_792_LC_7_32_2 (
            .in0(N__27574),
            .in1(N__31601),
            .in2(N__27085),
            .in3(N__27426),
            .lcout(),
            .ltout(n41_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_4_lut_LC_7_32_3.C_ON=1'b0;
    defparam i2_4_lut_4_lut_LC_7_32_3.SEQ_MODE=4'b0000;
    defparam i2_4_lut_4_lut_LC_7_32_3.LUT_INIT=16'b1111111111110111;
    LogicCell40 i2_4_lut_4_lut_LC_7_32_3 (
            .in0(N__45905),
            .in1(N__46299),
            .in2(N__27082),
            .in3(N__34317),
            .lcout(n35),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15262_4_lut_LC_7_32_4.C_ON=1'b0;
    defparam i15262_4_lut_LC_7_32_4.SEQ_MODE=4'b0000;
    defparam i15262_4_lut_LC_7_32_4.LUT_INIT=16'b0000000011110111;
    LogicCell40 i15262_4_lut_LC_7_32_4 (
            .in0(N__27575),
            .in1(N__27378),
            .in2(N__27475),
            .in3(N__27425),
            .lcout(),
            .ltout(n17479_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i57_4_lut_LC_7_32_5.C_ON=1'b0;
    defparam i57_4_lut_LC_7_32_5.SEQ_MODE=4'b0000;
    defparam i57_4_lut_LC_7_32_5.LUT_INIT=16'b1101000111000000;
    LogicCell40 i57_4_lut_LC_7_32_5 (
            .in0(N__45906),
            .in1(N__46300),
            .in2(N__27412),
            .in3(N__27409),
            .lcout(n38),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_690_LC_7_32_6 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_690_LC_7_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_690_LC_7_32_6 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_690_LC_7_32_6  (
            .in0(N__27352),
            .in1(N__27311),
            .in2(N__42622),
            .in3(N__27376),
            .lcout(\c0.n44_adj_2163 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15277_3_lut_4_lut_LC_7_32_7 .C_ON=1'b0;
    defparam \c0.i15277_3_lut_4_lut_LC_7_32_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15277_3_lut_4_lut_LC_7_32_7 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \c0.i15277_3_lut_4_lut_LC_7_32_7  (
            .in0(N__27379),
            .in1(N__46298),
            .in2(N__27358),
            .in3(N__27313),
            .lcout(\c0.n17475 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i15437_2_lut_3_lut_LC_9_17_1 .C_ON=1'b0;
    defparam \c0.tx2.i15437_2_lut_3_lut_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i15437_2_lut_3_lut_LC_9_17_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \c0.tx2.i15437_2_lut_3_lut_LC_9_17_1  (
            .in0(N__27268),
            .in1(N__30604),
            .in2(_gnd_net_),
            .in3(N__27230),
            .lcout(\c0.tx2_transmit_N_1997 ),
            .ltout(\c0.tx2_transmit_N_1997_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_transmit_2249_LC_9_17_2 .C_ON=1'b0;
    defparam \c0.tx2_transmit_2249_LC_9_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2_transmit_2249_LC_9_17_2 .LUT_INIT=16'b1000000011101110;
    LogicCell40 \c0.tx2_transmit_2249_LC_9_17_2  (
            .in0(N__32317),
            .in1(N__33516),
            .in2(N__27271),
            .in3(N__34275),
            .lcout(\c0.r_SM_Main_2_N_2036_0_adj_2261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50412),
            .ce(),
            .sr(N__33580));
    defparam \c0.tx2.i3_4_lut_LC_9_17_4 .C_ON=1'b0;
    defparam \c0.tx2.i3_4_lut_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i3_4_lut_LC_9_17_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx2.i3_4_lut_LC_9_17_4  (
            .in0(N__32203),
            .in1(N__34756),
            .in2(N__34735),
            .in3(N__34708),
            .lcout(\c0.tx2.n113 ),
            .ltout(\c0.tx2.n113_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_2_lut_3_lut_LC_9_17_5 .C_ON=1'b0;
    defparam \c0.tx2.i1_2_lut_3_lut_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_2_lut_3_lut_LC_9_17_5 .LUT_INIT=16'b1111111111001111;
    LogicCell40 \c0.tx2.i1_2_lut_3_lut_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(N__30603),
            .in2(N__27262),
            .in3(N__27229),
            .lcout(n491),
            .ltout(n491_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_9_17_6.C_ON=1'b0;
    defparam i1_3_lut_LC_9_17_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_9_17_6.LUT_INIT=16'b0000000011000000;
    LogicCell40 i1_3_lut_LC_9_17_6 (
            .in0(_gnd_net_),
            .in1(N__33515),
            .in2(N__27196),
            .in3(N__27939),
            .lcout(n17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i20_LC_9_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i20_LC_9_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i20_LC_9_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i20_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__27981),
            .in2(_gnd_net_),
            .in3(N__34648),
            .lcout(\c0.FRAME_MATCHER_state_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50428),
            .ce(),
            .sr(N__28012));
    defparam \c0.FRAME_MATCHER_state_i24_LC_9_19_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i24_LC_9_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i24_LC_9_19_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i24_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__29473),
            .in2(_gnd_net_),
            .in3(N__34613),
            .lcout(\c0.FRAME_MATCHER_state_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50436),
            .ce(),
            .sr(N__29434));
    defparam \c0.FRAME_MATCHER_state_i18_LC_9_20_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i18_LC_9_20_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i18_LC_9_20_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i18_LC_9_20_0  (
            .in0(N__34645),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27878),
            .lcout(\c0.FRAME_MATCHER_state_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50442),
            .ce(),
            .sr(N__27841));
    defparam \c0.i6_3_lut_4_lut_LC_9_21_0 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_LC_9_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_3_lut_4_lut_LC_9_21_0  (
            .in0(N__28000),
            .in1(N__27982),
            .in2(N__30088),
            .in3(N__27864),
            .lcout(n9460),
            .ltout(n9460_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_519_LC_9_21_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_519_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_519_LC_9_21_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \c0.i1_2_lut_adj_519_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27910),
            .in3(N__33535),
            .lcout(n9462),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i64_LC_9_21_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i64_LC_9_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i64_LC_9_21_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i64_LC_9_21_4  (
            .in0(N__51224),
            .in1(N__44944),
            .in2(_gnd_net_),
            .in3(N__41318),
            .lcout(data_out_frame2_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50454),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_736_LC_9_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_736_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_736_LC_9_21_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_736_LC_9_21_5  (
            .in0(N__27865),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29954),
            .lcout(\c0.n16343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__6__2267_LC_9_21_6 .C_ON=1'b0;
    defparam \c0.data_in_1__6__2267_LC_9_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__6__2267_LC_9_21_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_1__6__2267_LC_9_21_6  (
            .in0(N__27835),
            .in1(N__27596),
            .in2(_gnd_net_),
            .in3(N__27790),
            .lcout(data_in_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50454),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3112_3_lut_4_lut_LC_9_21_7 .C_ON=1'b0;
    defparam \c0.i3112_3_lut_4_lut_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3112_3_lut_4_lut_LC_9_21_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \c0.i3112_3_lut_4_lut_LC_9_21_7  (
            .in0(N__33320),
            .in1(N__33352),
            .in2(N__28342),
            .in3(N__32318),
            .lcout(\c0.n5543 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_LC_9_22_0 .C_ON=1'b0;
    defparam \c0.i19_4_lut_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_LC_9_22_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i19_4_lut_LC_9_22_0  (
            .in0(N__28321),
            .in1(N__28291),
            .in2(N__28258),
            .in3(N__28169),
            .lcout(\c0.n48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i10_LC_9_22_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i10_LC_9_22_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i10_LC_9_22_1 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i10_LC_9_22_1  (
            .in0(N__33276),
            .in1(N__32918),
            .in2(_gnd_net_),
            .in3(N__28204),
            .lcout(\c0.FRAME_MATCHER_i_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50464),
            .ce(),
            .sr(N__28156));
    defparam \c0.i1_2_lut_4_lut_adj_665_LC_9_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_665_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_665_LC_9_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_665_LC_9_22_2  (
            .in0(N__40905),
            .in1(N__35232),
            .in2(N__43909),
            .in3(N__48882),
            .lcout(\c0.n6_adj_2293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_520_LC_9_22_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_520_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_520_LC_9_22_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_3_lut_adj_520_LC_9_22_3  (
            .in0(N__48883),
            .in1(_gnd_net_),
            .in2(N__35239),
            .in3(N__43906),
            .lcout(),
            .ltout(\c0.n9819_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_449_LC_9_22_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_449_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_449_LC_9_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_449_LC_9_22_4  (
            .in0(N__37021),
            .in1(N__49633),
            .in2(N__28144),
            .in3(N__43585),
            .lcout(\c0.n17_adj_2193 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15294_2_lut_LC_9_22_5 .C_ON=1'b0;
    defparam \c0.i15294_2_lut_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15294_2_lut_LC_9_22_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i15294_2_lut_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(N__40904),
            .in2(_gnd_net_),
            .in3(N__48211),
            .lcout(\c0.n17560 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i25_LC_9_23_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i25_LC_9_23_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i25_LC_9_23_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i25_LC_9_23_0  (
            .in0(N__34646),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28132),
            .lcout(\c0.FRAME_MATCHER_state_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50476),
            .ce(),
            .sr(N__28102));
    defparam \c0.FRAME_MATCHER_i_i17_LC_9_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i17_LC_9_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i17_LC_9_24_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i17_LC_9_24_0  (
            .in0(N__33277),
            .in1(N__32988),
            .in2(_gnd_net_),
            .in3(N__28093),
            .lcout(\c0.FRAME_MATCHER_i_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50489),
            .ce(),
            .sr(N__28666));
    defparam \c0.i7_4_lut_adj_656_LC_9_25_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_656_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_656_LC_9_25_1 .LUT_INIT=16'b1111011001101111;
    LogicCell40 \c0.i7_4_lut_adj_656_LC_9_25_1  (
            .in0(N__29132),
            .in1(N__28654),
            .in2(N__28615),
            .in3(N__30192),
            .lcout(),
            .ltout(\c0.n23_adj_2341_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_660_LC_9_25_2 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_660_LC_9_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_660_LC_9_25_2 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \c0.i14_4_lut_adj_660_LC_9_25_2  (
            .in0(N__28579),
            .in1(N__28540),
            .in2(N__28528),
            .in3(N__28525),
            .lcout(\c0.n30_adj_2345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_452_LC_9_25_4 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_452_LC_9_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_452_LC_9_25_4 .LUT_INIT=16'b1011111111101111;
    LogicCell40 \c0.i11_4_lut_adj_452_LC_9_25_4  (
            .in0(N__28495),
            .in1(N__29005),
            .in2(N__28486),
            .in3(N__28471),
            .lcout(\c0.n27_adj_2196 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14914_3_lut_LC_9_25_6 .C_ON=1'b0;
    defparam \c0.i14914_3_lut_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i14914_3_lut_LC_9_25_6 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \c0.i14914_3_lut_LC_9_25_6  (
            .in0(N__40900),
            .in1(N__37478),
            .in2(_gnd_net_),
            .in3(N__35018),
            .lcout(),
            .ltout(\c0.n17352_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i1_LC_9_25_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i1_LC_9_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i1_LC_9_25_7 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.data_out_frame2_0___i1_LC_9_25_7  (
            .in0(N__37479),
            .in1(N__34956),
            .in2(N__28453),
            .in3(N__37548),
            .lcout(\c0.data_out_frame2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50499),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_460_LC_9_26_0 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_460_LC_9_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_460_LC_9_26_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15_4_lut_adj_460_LC_9_26_0  (
            .in0(N__28420),
            .in1(N__29062),
            .in2(N__28450),
            .in3(N__28441),
            .lcout(\c0.n15846 ),
            .ltout(\c0.n15846_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14903_3_lut_LC_9_26_1 .C_ON=1'b0;
    defparam \c0.i14903_3_lut_LC_9_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14903_3_lut_LC_9_26_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.i14903_3_lut_LC_9_26_1  (
            .in0(_gnd_net_),
            .in1(N__37472),
            .in2(N__28432),
            .in3(N__37382),
            .lcout(\c0.n17769 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_442_LC_9_26_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_442_LC_9_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_442_LC_9_26_2 .LUT_INIT=16'b1111111101111011;
    LogicCell40 \c0.i10_4_lut_adj_442_LC_9_26_2  (
            .in0(N__28938),
            .in1(N__28429),
            .in2(N__31057),
            .in3(N__28960),
            .lcout(\c0.n26_adj_2184 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_431_LC_9_26_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_431_LC_9_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_431_LC_9_26_4 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \c0.i7_4_lut_adj_431_LC_9_26_4  (
            .in0(N__28414),
            .in1(N__28402),
            .in2(N__28363),
            .in3(N__29137),
            .lcout(),
            .ltout(\c0.n23_adj_2156_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_LC_9_26_5 .C_ON=1'b0;
    defparam \c0.i12_4_lut_LC_9_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_LC_9_26_5 .LUT_INIT=16'b1111011111111011;
    LogicCell40 \c0.i12_4_lut_LC_9_26_5  (
            .in0(N__28815),
            .in1(N__29101),
            .in2(N__29089),
            .in3(N__29086),
            .lcout(\c0.n28_adj_2183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1034_2_lut_LC_9_26_7 .C_ON=1'b0;
    defparam \c0.i1034_2_lut_LC_9_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1034_2_lut_LC_9_26_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1034_2_lut_LC_9_26_7  (
            .in0(_gnd_net_),
            .in1(N__29056),
            .in2(_gnd_net_),
            .in3(N__30316),
            .lcout(\c0.n2340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_434_LC_9_27_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_434_LC_9_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_434_LC_9_27_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \c0.i3_4_lut_adj_434_LC_9_27_0  (
            .in0(N__28704),
            .in1(N__28833),
            .in2(N__28996),
            .in3(N__28978),
            .lcout(\c0.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_409_LC_9_27_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_409_LC_9_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_409_LC_9_27_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \c0.i4_4_lut_adj_409_LC_9_27_1  (
            .in0(N__28954),
            .in1(N__28939),
            .in2(N__28918),
            .in3(N__28894),
            .lcout(),
            .ltout(\c0.n20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_LC_9_27_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_LC_9_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_LC_9_27_2 .LUT_INIT=16'b1111101111110111;
    LogicCell40 \c0.i10_4_lut_LC_9_27_2  (
            .in0(N__28876),
            .in1(N__28858),
            .in2(N__28837),
            .in3(N__28834),
            .lcout(\c0.n26_adj_2147 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i74_LC_9_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i74_LC_9_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i74_LC_9_27_4 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i74_LC_9_27_4  (
            .in0(N__30679),
            .in1(N__28816),
            .in2(N__28804),
            .in3(N__31133),
            .lcout(\c0.data_in_frame_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50519),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i78_LC_9_27_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i78_LC_9_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i78_LC_9_27_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i78_LC_9_27_5  (
            .in0(N__31134),
            .in1(N__28795),
            .in2(N__31231),
            .in3(N__28705),
            .lcout(\c0.data_in_frame_9_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50519),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_45_LC_9_27_6 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_45_LC_9_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.o_Tx_Serial_45_LC_9_27_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx2.o_Tx_Serial_45_LC_9_27_6  (
            .in0(N__28677),
            .in1(N__31545),
            .in2(_gnd_net_),
            .in3(N__29275),
            .lcout(tx2_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50519),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14905_3_lut_LC_9_27_7 .C_ON=1'b0;
    defparam \c0.i14905_3_lut_LC_9_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i14905_3_lut_LC_9_27_7 .LUT_INIT=16'b0000101011111010;
    LogicCell40 \c0.i14905_3_lut_LC_9_27_7  (
            .in0(N__35853),
            .in1(_gnd_net_),
            .in2(N__37483),
            .in3(N__35004),
            .lcout(\c0.n17343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i1_LC_9_28_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i1_LC_9_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i1_LC_9_28_2 .LUT_INIT=16'b1101001000000000;
    LogicCell40 \c0.tx2.r_Bit_Index_i1_LC_9_28_2  (
            .in0(N__35343),
            .in1(N__29184),
            .in2(N__35391),
            .in3(N__29193),
            .lcout(r_Bit_Index_1_adj_2456),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50528),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i2_LC_9_28_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i2_LC_9_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i2_LC_9_28_4 .LUT_INIT=16'b1001101000000000;
    LogicCell40 \c0.tx2.r_Bit_Index_i2_LC_9_28_4  (
            .in0(N__29256),
            .in1(N__29185),
            .in2(N__29266),
            .in3(N__29194),
            .lcout(r_Bit_Index_2_adj_2455),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50528),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.n17903_bdd_4_lut_LC_9_28_5 .C_ON=1'b0;
    defparam \c0.tx2.n17903_bdd_4_lut_LC_9_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.n17903_bdd_4_lut_LC_9_28_5 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.tx2.n17903_bdd_4_lut_LC_9_28_5  (
            .in0(N__35101),
            .in1(N__35381),
            .in2(N__51484),
            .in3(N__35314),
            .lcout(\c0.tx2.n17906 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_9_28_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_9_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_9_28_6 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_9_28_6  (
            .in0(N__36793),
            .in1(N__35342),
            .in2(N__35390),
            .in3(N__32509),
            .lcout(),
            .ltout(\c0.tx2.n18113_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.n18113_bdd_4_lut_LC_9_28_7 .C_ON=1'b0;
    defparam \c0.tx2.n18113_bdd_4_lut_LC_9_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.n18113_bdd_4_lut_LC_9_28_7 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.tx2.n18113_bdd_4_lut_LC_9_28_7  (
            .in0(N__34822),
            .in1(N__33949),
            .in2(N__29197),
            .in3(N__35380),
            .lcout(\c0.tx2.n18116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i14834_3_lut_LC_9_29_0 .C_ON=1'b0;
    defparam \c0.tx2.i14834_3_lut_LC_9_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i14834_3_lut_LC_9_29_0 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \c0.tx2.i14834_3_lut_LC_9_29_0  (
            .in0(N__29232),
            .in1(N__31027),
            .in2(_gnd_net_),
            .in3(N__29182),
            .lcout(n10398),
            .ltout(n10398_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i0_LC_9_29_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i0_LC_9_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i0_LC_9_29_1 .LUT_INIT=16'b1010000001010000;
    LogicCell40 \c0.tx2.r_Bit_Index_i0_LC_9_29_1  (
            .in0(N__29183),
            .in1(_gnd_net_),
            .in2(N__29155),
            .in3(N__35349),
            .lcout(r_Bit_Index_0_adj_2457),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50539),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i11207211_i1_3_lut_LC_9_29_2 .C_ON=1'b0;
    defparam \c0.tx2.i11207211_i1_3_lut_LC_9_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i11207211_i1_3_lut_LC_9_29_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.tx2.i11207211_i1_3_lut_LC_9_29_2  (
            .in0(N__29152),
            .in1(N__29146),
            .in2(_gnd_net_),
            .in3(N__29255),
            .lcout(),
            .ltout(\c0.tx2.o_Tx_Serial_N_2064_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_29_3 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_29_3 .LUT_INIT=16'b1100110011110011;
    LogicCell40 \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_29_3  (
            .in0(_gnd_net_),
            .in1(N__31026),
            .in2(N__29347),
            .in3(N__29340),
            .lcout(n3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2595_2_lut_LC_9_29_4 .C_ON=1'b0;
    defparam \c0.tx2.i2595_2_lut_LC_9_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2595_2_lut_LC_9_29_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.tx2.i2595_2_lut_LC_9_29_4  (
            .in0(N__35348),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35386),
            .lcout(n5029),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_2_lut_3_lut_LC_9_29_5 .C_ON=1'b0;
    defparam \c0.tx2.i2_2_lut_3_lut_LC_9_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_2_lut_3_lut_LC_9_29_5 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \c0.tx2.i2_2_lut_3_lut_LC_9_29_5  (
            .in0(N__35385),
            .in1(_gnd_net_),
            .in2(N__29257),
            .in3(N__35347),
            .lcout(\c0.tx2.n13281 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_9_29_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_9_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_9_29_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_9_29_7  (
            .in0(N__42968),
            .in1(N__47138),
            .in2(_gnd_net_),
            .in3(N__52043),
            .lcout(\c0.n8_adj_2160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_9_30_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_9_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_9_30_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_9_30_1  (
            .in0(N__52044),
            .in1(N__34075),
            .in2(_gnd_net_),
            .in3(N__33976),
            .lcout(),
            .ltout(\c0.n2_adj_2266_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18095_bdd_4_lut_LC_9_30_2 .C_ON=1'b0;
    defparam \c0.n18095_bdd_4_lut_LC_9_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18095_bdd_4_lut_LC_9_30_2 .LUT_INIT=16'b1100110011100010;
    LogicCell40 \c0.n18095_bdd_4_lut_LC_9_30_2  (
            .in0(N__41911),
            .in1(N__52150),
            .in2(N__29221),
            .in3(N__52408),
            .lcout(),
            .ltout(\c0.n18098_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_LC_9_30_3 .C_ON=1'b0;
    defparam \c0.i24_4_lut_LC_9_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_LC_9_30_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.i24_4_lut_LC_9_30_3  (
            .in0(N__52409),
            .in1(N__31564),
            .in2(N__29218),
            .in3(N__43150),
            .lcout(),
            .ltout(\c0.n10_adj_2139_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i0_LC_9_30_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i0_LC_9_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i0_LC_9_30_4 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \c0.tx.r_Tx_Data_i0_LC_9_30_4  (
            .in0(N__29428),
            .in1(N__35604),
            .in2(N__29215),
            .in3(N__35518),
            .lcout(r_Tx_Data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50548),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_50_LC_9_30_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_50_LC_9_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_50_LC_9_30_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.rx.r_Rx_Data_50_LC_9_30_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29212),
            .lcout(r_Rx_Data),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50548),
            .ce(),
            .sr(_gnd_net_));
    defparam i14956_3_lut_LC_9_30_7.C_ON=1'b0;
    defparam i14956_3_lut_LC_9_30_7.SEQ_MODE=4'b0000;
    defparam i14956_3_lut_LC_9_30_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 i14956_3_lut_LC_9_30_7 (
            .in0(N__29391),
            .in1(N__29427),
            .in2(_gnd_net_),
            .in3(N__31379),
            .lcout(n17394),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__7__2213_LC_9_31_1 .C_ON=1'b0;
    defparam \c0.data_out_3__7__2213_LC_9_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__7__2213_LC_9_31_1 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \c0.data_out_3__7__2213_LC_9_31_1  (
            .in0(N__45515),
            .in1(N__32098),
            .in2(N__45929),
            .in3(N__46422),
            .lcout(data_out_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50557),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_9_31_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_9_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_9_31_4 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_9_31_4  (
            .in0(N__29407),
            .in1(N__52232),
            .in2(N__47101),
            .in3(N__51970),
            .lcout(n10_adj_2426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30_4_lut_LC_9_31_5 .C_ON=1'b0;
    defparam \c0.i30_4_lut_LC_9_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i30_4_lut_LC_9_31_5 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \c0.i30_4_lut_LC_9_31_5  (
            .in0(N__51971),
            .in1(N__35653),
            .in2(N__52264),
            .in3(N__46756),
            .lcout(),
            .ltout(\c0.n15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i31_4_lut_LC_9_31_6 .C_ON=1'b0;
    defparam \c0.i31_4_lut_LC_9_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i31_4_lut_LC_9_31_6 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \c0.i31_4_lut_LC_9_31_6  (
            .in0(N__32158),
            .in1(N__43120),
            .in2(N__29398),
            .in3(N__52460),
            .lcout(),
            .ltout(\c0.n12_adj_2150_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i2_LC_9_31_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i2_LC_9_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i2_LC_9_31_7 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.tx.r_Tx_Data_i2_LC_9_31_7  (
            .in0(N__35521),
            .in1(N__29392),
            .in2(N__29395),
            .in3(N__35564),
            .lcout(r_Tx_Data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50557),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_LC_9_32_0.C_ON=1'b0;
    defparam i24_4_lut_LC_9_32_0.SEQ_MODE=4'b0000;
    defparam i24_4_lut_LC_9_32_0.LUT_INIT=16'b0101000011001100;
    LogicCell40 i24_4_lut_LC_9_32_0 (
            .in0(N__52459),
            .in1(N__29557),
            .in2(N__29380),
            .in3(N__43151),
            .lcout(),
            .ltout(n10_adj_2407_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i4_LC_9_32_1 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i4_LC_9_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i4_LC_9_32_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \c0.tx.r_Tx_Data_i4_LC_9_32_1  (
            .in0(N__35522),
            .in1(N__35603),
            .in2(N__29371),
            .in3(N__29361),
            .lcout(r_Tx_Data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50567),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15288_2_lut_LC_9_32_4 .C_ON=1'b0;
    defparam \c0.i15288_2_lut_LC_9_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15288_2_lut_LC_9_32_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.i15288_2_lut_LC_9_32_4  (
            .in0(N__51997),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32478),
            .lcout(),
            .ltout(\c0.n17590_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18023_bdd_4_lut_LC_9_32_5 .C_ON=1'b0;
    defparam \c0.n18023_bdd_4_lut_LC_9_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18023_bdd_4_lut_LC_9_32_5 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n18023_bdd_4_lut_LC_9_32_5  (
            .in0(N__42898),
            .in1(N__32017),
            .in2(N__29560),
            .in3(N__52458),
            .lcout(n18026),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15348_2_lut_LC_9_32_7 .C_ON=1'b0;
    defparam \c0.i15348_2_lut_LC_9_32_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15348_2_lut_LC_9_32_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15348_2_lut_LC_9_32_7  (
            .in0(_gnd_net_),
            .in1(N__42383),
            .in2(_gnd_net_),
            .in3(N__51996),
            .lcout(\c0.n17547 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i16_LC_10_17_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i16_LC_10_17_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i16_LC_10_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i16_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__32396),
            .in2(_gnd_net_),
            .in3(N__34650),
            .lcout(\c0.FRAME_MATCHER_state_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50422),
            .ce(),
            .sr(N__29551));
    defparam \c0.FRAME_MATCHER_state_i17_LC_10_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i17_LC_10_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i17_LC_10_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i17_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__30057),
            .in2(_gnd_net_),
            .in3(N__34649),
            .lcout(\c0.FRAME_MATCHER_state_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50430),
            .ce(),
            .sr(N__30034));
    defparam \c0.i3_4_lut_adj_495_LC_10_19_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_495_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_495_LC_10_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_495_LC_10_19_0  (
            .in0(N__32192),
            .in1(N__30055),
            .in2(N__29476),
            .in3(N__29503),
            .lcout(\c0.n16761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i28_LC_10_19_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i28_LC_10_19_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i28_LC_10_19_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i28_LC_10_19_1  (
            .in0(N__29505),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34641),
            .lcout(\c0.FRAME_MATCHER_state_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50437),
            .ce(),
            .sr(N__29485));
    defparam \c0.i1_2_lut_adj_758_LC_10_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_758_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_758_LC_10_19_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.i1_2_lut_adj_758_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29983),
            .in3(N__29504),
            .lcout(\c0.n16353 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_LC_10_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_LC_10_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__32193),
            .in2(_gnd_net_),
            .in3(N__29972),
            .lcout(\c0.n16377 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_749_LC_10_19_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_749_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_749_LC_10_19_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \c0.i1_2_lut_adj_749_LC_10_19_4  (
            .in0(N__29472),
            .in1(_gnd_net_),
            .in2(N__29982),
            .in3(_gnd_net_),
            .lcout(\c0.n16361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_734_LC_10_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_734_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_734_LC_10_19_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_734_LC_10_19_5  (
            .in0(N__30056),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29974),
            .lcout(\c0.n16345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_705_LC_10_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_705_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_705_LC_10_19_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_705_LC_10_19_7  (
            .in0(N__30026),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29973),
            .lcout(\c0.n16339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i12_LC_10_20_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i12_LC_10_20_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i12_LC_10_20_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i12_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__32610),
            .in2(_gnd_net_),
            .in3(N__34647),
            .lcout(\c0.FRAME_MATCHER_state_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50443),
            .ce(),
            .sr(N__32542));
    defparam \c0.data_out_frame2_0___i147_LC_10_21_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i147_LC_10_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i147_LC_10_21_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i147_LC_10_21_0  (
            .in0(N__36442),
            .in1(N__32529),
            .in2(_gnd_net_),
            .in3(N__51250),
            .lcout(data_out_frame2_18_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50455),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_640_LC_10_21_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_640_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_640_LC_10_21_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_640_LC_10_21_1  (
            .in0(N__30133),
            .in1(N__29823),
            .in2(N__29788),
            .in3(N__29776),
            .lcout(\c0.n13464 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_10_21_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_10_21_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_10_21_4  (
            .in0(N__48194),
            .in1(N__33556),
            .in2(_gnd_net_),
            .in3(N__34913),
            .lcout(\c0.n5_adj_2322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14911_3_lut_LC_10_21_5 .C_ON=1'b0;
    defparam \c0.i14911_3_lut_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i14911_3_lut_LC_10_21_5 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \c0.i14911_3_lut_LC_10_21_5  (
            .in0(N__37109),
            .in1(N__37434),
            .in2(_gnd_net_),
            .in3(N__35037),
            .lcout(),
            .ltout(\c0.n17349_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i2_LC_10_21_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i2_LC_10_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i2_LC_10_21_6 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.data_out_frame2_0___i2_LC_10_21_6  (
            .in0(N__37435),
            .in1(N__37538),
            .in2(N__29752),
            .in3(N__34978),
            .lcout(\c0.data_out_frame2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50455),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_238_Select_0_i3_2_lut_LC_10_21_7 .C_ON=1'b0;
    defparam \c0.select_238_Select_0_i3_2_lut_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_238_Select_0_i3_2_lut_LC_10_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_238_Select_0_i3_2_lut_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(N__29743),
            .in2(_gnd_net_),
            .in3(N__29581),
            .lcout(\c0.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_10_22_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_10_22_0 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_10_22_0  (
            .in0(N__48209),
            .in1(N__30148),
            .in2(N__35071),
            .in3(N__48541),
            .lcout(\c0.n6_adj_2187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_10_22_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_10_22_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_10_22_1  (
            .in0(N__38607),
            .in1(N__48208),
            .in2(_gnd_net_),
            .in3(N__41521),
            .lcout(),
            .ltout(\c0.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_10_22_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_10_22_2 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_10_22_2  (
            .in0(N__48210),
            .in1(N__48542),
            .in2(N__30139),
            .in3(N__39021),
            .lcout(\c0.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14890_3_lut_LC_10_22_3 .C_ON=1'b0;
    defparam \c0.i14890_3_lut_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14890_3_lut_LC_10_22_3 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \c0.i14890_3_lut_LC_10_22_3  (
            .in0(N__37431),
            .in1(N__49525),
            .in2(_gnd_net_),
            .in3(N__35036),
            .lcout(),
            .ltout(\c0.n17328_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i8_LC_10_22_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i8_LC_10_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i8_LC_10_22_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.data_out_frame2_0___i8_LC_10_22_4  (
            .in0(N__37539),
            .in1(N__37432),
            .in2(N__30136),
            .in3(N__34977),
            .lcout(\c0.data_out_frame2_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50465),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_596_LC_10_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_596_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_596_LC_10_22_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_596_LC_10_22_5  (
            .in0(_gnd_net_),
            .in1(N__34912),
            .in2(_gnd_net_),
            .in3(N__38524),
            .lcout(\c0.n9758 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_LC_10_22_7 .C_ON=1'b0;
    defparam \c0.i1_3_lut_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_LC_10_22_7 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.i1_3_lut_LC_10_22_7  (
            .in0(N__30129),
            .in1(N__34276),
            .in2(_gnd_net_),
            .in3(N__32397),
            .lcout(\c0.n16905 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_699_LC_10_23_0 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_699_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_699_LC_10_23_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_699_LC_10_23_0  (
            .in0(N__41703),
            .in1(_gnd_net_),
            .in2(N__33568),
            .in3(N__36073),
            .lcout(\c0.n16_adj_2197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i124_LC_10_23_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i124_LC_10_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i124_LC_10_23_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i124_LC_10_23_1  (
            .in0(N__36074),
            .in1(N__48839),
            .in2(_gnd_net_),
            .in3(N__51273),
            .lcout(data_out_frame2_15_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50477),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14899_3_lut_LC_10_23_3 .C_ON=1'b0;
    defparam \c0.i14899_3_lut_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14899_3_lut_LC_10_23_3 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \c0.i14899_3_lut_LC_10_23_3  (
            .in0(N__35809),
            .in1(N__37433),
            .in2(_gnd_net_),
            .in3(N__35035),
            .lcout(),
            .ltout(\c0.n17337_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i5_LC_10_23_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i5_LC_10_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i5_LC_10_23_4 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \c0.data_out_frame2_0___i5_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(N__37541),
            .in2(N__30349),
            .in3(N__31294),
            .lcout(\c0.data_out_frame2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50477),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i91_LC_10_23_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i91_LC_10_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i91_LC_10_23_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i91_LC_10_23_5  (
            .in0(N__36622),
            .in1(N__40861),
            .in2(_gnd_net_),
            .in3(N__51274),
            .lcout(data_out_frame2_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50477),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i4_LC_10_23_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i4_LC_10_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i4_LC_10_23_6 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \c0.data_out_frame2_0___i4_LC_10_23_6  (
            .in0(N__32494),
            .in1(N__37540),
            .in2(_gnd_net_),
            .in3(N__31293),
            .lcout(\c0.data_out_frame2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50477),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1032_2_lut_LC_10_24_1 .C_ON=1'b0;
    defparam \c0.i1032_2_lut_LC_10_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1032_2_lut_LC_10_24_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1032_2_lut_LC_10_24_1  (
            .in0(_gnd_net_),
            .in1(N__30346),
            .in2(_gnd_net_),
            .in3(N__30315),
            .lcout(\c0.n2338 ),
            .ltout(\c0.n2338_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_661_LC_10_24_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_661_LC_10_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_661_LC_10_24_2 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \c0.i1_4_lut_adj_661_LC_10_24_2  (
            .in0(N__30244),
            .in1(N__30223),
            .in2(N__30199),
            .in3(N__30196),
            .lcout(),
            .ltout(\c0.n17_adj_2346_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_662_LC_10_24_3 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_662_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_662_LC_10_24_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15_4_lut_adj_662_LC_10_24_3  (
            .in0(N__30172),
            .in1(N__30538),
            .in2(N__30160),
            .in3(N__30157),
            .lcout(n31),
            .ltout(n31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_653_LC_10_24_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_653_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_653_LC_10_24_4 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \c0.i1_4_lut_adj_653_LC_10_24_4  (
            .in0(N__33356),
            .in1(N__33322),
            .in2(N__30151),
            .in3(N__34282),
            .lcout(\c0.n5_adj_2339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i127_LC_10_24_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i127_LC_10_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i127_LC_10_24_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i127_LC_10_24_6  (
            .in0(N__51279),
            .in1(N__49102),
            .in2(_gnd_net_),
            .in3(N__44378),
            .lcout(data_out_frame2_15_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50490),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i84_LC_10_24_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i84_LC_10_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i84_LC_10_24_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i84_LC_10_24_7  (
            .in0(N__36731),
            .in1(N__41815),
            .in2(_gnd_net_),
            .in3(N__51280),
            .lcout(data_out_frame2_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50490),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15387_3_lut_LC_10_25_0 .C_ON=1'b0;
    defparam \c0.i15387_3_lut_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15387_3_lut_LC_10_25_0 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \c0.i15387_3_lut_LC_10_25_0  (
            .in0(N__48227),
            .in1(N__38707),
            .in2(_gnd_net_),
            .in3(N__48667),
            .lcout(\c0.n17571 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Active_47_LC_10_25_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Active_47_LC_10_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Active_47_LC_10_25_2 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \c0.tx2.r_Tx_Active_47_LC_10_25_2  (
            .in0(N__31039),
            .in1(N__30597),
            .in2(_gnd_net_),
            .in3(N__30910),
            .lcout(\c0.tx2.tx2_active ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50500),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14896_3_lut_LC_10_25_3 .C_ON=1'b0;
    defparam \c0.i14896_3_lut_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14896_3_lut_LC_10_25_3 .LUT_INIT=16'b0111010001110100;
    LogicCell40 \c0.i14896_3_lut_LC_10_25_3  (
            .in0(N__35017),
            .in1(N__37476),
            .in2(N__38717),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n17334_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i6_LC_10_25_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i6_LC_10_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i6_LC_10_25_4 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.data_out_frame2_0___i6_LC_10_25_4  (
            .in0(N__37477),
            .in1(N__37553),
            .in2(N__30583),
            .in3(N__34957),
            .lcout(\c0.data_out_frame2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50500),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_10_25_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_10_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_10_25_5 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_10_25_5  (
            .in0(N__43963),
            .in1(N__48665),
            .in2(N__41287),
            .in3(N__48226),
            .lcout(\c0.n6_adj_2278 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_658_LC_10_25_6 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_658_LC_10_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_658_LC_10_25_6 .LUT_INIT=16'b1101111001111011;
    LogicCell40 \c0.i2_4_lut_adj_658_LC_10_25_6  (
            .in0(N__30579),
            .in1(N__30619),
            .in2(N__31759),
            .in3(N__30555),
            .lcout(\c0.n18_adj_2343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i4_LC_10_25_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i4_LC_10_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i4_LC_10_25_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i4_LC_10_25_7  (
            .in0(N__30524),
            .in1(N__30371),
            .in2(_gnd_net_),
            .in3(N__30442),
            .lcout(data_in_frame_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50500),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i77_LC_10_26_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i77_LC_10_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i77_LC_10_26_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i77_LC_10_26_0  (
            .in0(N__39210),
            .in1(N__35215),
            .in2(_gnd_net_),
            .in3(N__51180),
            .lcout(data_out_frame2_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50511),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17915_bdd_4_lut_LC_10_26_2 .C_ON=1'b0;
    defparam \c0.n17915_bdd_4_lut_LC_10_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.n17915_bdd_4_lut_LC_10_26_2 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \c0.n17915_bdd_4_lut_LC_10_26_2  (
            .in0(N__41594),
            .in1(N__48666),
            .in2(N__49603),
            .in3(N__33655),
            .lcout(),
            .ltout(\c0.n17918_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15636_LC_10_26_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15636_LC_10_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15636_LC_10_26_3 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15636_LC_10_26_3  (
            .in0(N__41662),
            .in1(N__51644),
            .in2(N__31303),
            .in3(N__47711),
            .lcout(\c0.n18107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i3_LC_10_26_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i3_LC_10_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i3_LC_10_26_5 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \c0.data_out_frame2_0___i3_LC_10_26_5  (
            .in0(N__37554),
            .in1(N__31300),
            .in2(_gnd_net_),
            .in3(N__31284),
            .lcout(\c0.data_out_frame2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50511),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_LC_10_26_7 .C_ON=1'b0;
    defparam \c0.i15_4_lut_LC_10_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_LC_10_26_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15_4_lut_LC_10_26_7  (
            .in0(N__31273),
            .in1(N__31261),
            .in2(N__31249),
            .in3(N__31240),
            .lcout(\c0.n16148 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i86_LC_10_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i86_LC_10_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i86_LC_10_27_0 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i86_LC_10_27_0  (
            .in0(N__31936),
            .in1(N__31053),
            .in2(N__31230),
            .in3(N__31136),
            .lcout(\c0.data_in_frame_10_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50520),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_4_lut_LC_10_27_1 .C_ON=1'b0;
    defparam \c0.tx2.i1_4_lut_LC_10_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_4_lut_LC_10_27_1 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \c0.tx2.i1_4_lut_LC_10_27_1  (
            .in0(N__31552),
            .in1(N__31038),
            .in2(N__30943),
            .in3(N__30925),
            .lcout(\c0.tx2.n10101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15533_LC_10_27_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15533_LC_10_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15533_LC_10_27_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15533_LC_10_27_2  (
            .in0(N__30901),
            .in1(N__48641),
            .in2(N__35986),
            .in3(N__48186),
            .lcout(\c0.n17981 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i0_LC_10_27_3 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i0_LC_10_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i0_LC_10_27_3 .LUT_INIT=16'b0001010100010000;
    LogicCell40 \c0.rx.r_SM_Main_i0_LC_10_27_3  (
            .in0(N__30883),
            .in1(N__30802),
            .in2(N__30787),
            .in3(N__33661),
            .lcout(r_SM_Main_0_adj_2441),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50520),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i18_LC_10_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i18_LC_10_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i18_LC_10_27_6 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i18_LC_10_27_6  (
            .in0(N__31934),
            .in1(N__30618),
            .in2(N__30694),
            .in3(N__32007),
            .lcout(\c0.data_in_frame_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50520),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i21_LC_10_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i21_LC_10_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i21_LC_10_27_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i21_LC_10_27_7  (
            .in0(N__32008),
            .in1(N__31935),
            .in2(N__31834),
            .in3(N__31758),
            .lcout(\c0.data_in_frame_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50520),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_10_28_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_10_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_10_28_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_10_28_0  (
            .in0(N__34020),
            .in1(N__34035),
            .in2(_gnd_net_),
            .in3(N__51993),
            .lcout(\c0.n2_adj_2298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14792_2_lut_3_lut_LC_10_28_1 .C_ON=1'b0;
    defparam \c0.i14792_2_lut_3_lut_LC_10_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14792_2_lut_3_lut_LC_10_28_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i14792_2_lut_3_lut_LC_10_28_1  (
            .in0(N__45920),
            .in1(N__31741),
            .in2(_gnd_net_),
            .in3(N__31671),
            .lcout(n17230),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__7__2229_LC_10_28_3 .C_ON=1'b0;
    defparam \c0.data_out_1__7__2229_LC_10_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__7__2229_LC_10_28_3 .LUT_INIT=16'b1000110011011100;
    LogicCell40 \c0.data_out_1__7__2229_LC_10_28_3  (
            .in0(N__45544),
            .in1(N__31573),
            .in2(N__45982),
            .in3(N__46449),
            .lcout(data_out_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50529),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15355_2_lut_LC_10_28_5 .C_ON=1'b0;
    defparam \c0.i15355_2_lut_LC_10_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15355_2_lut_LC_10_28_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.i15355_2_lut_LC_10_28_5  (
            .in0(N__51994),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31572),
            .lcout(\c0.n17585 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i10_4_lut_LC_10_28_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i10_4_lut_LC_10_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i10_4_lut_LC_10_28_6 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i10_4_lut_LC_10_28_6  (
            .in0(N__33904),
            .in1(N__52257),
            .in2(N__39787),
            .in3(N__51995),
            .lcout(\c0.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i0_LC_10_28_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i0_LC_10_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i0_LC_10_28_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx2.r_Clock_Count__i0_LC_10_28_7  (
            .in0(N__31551),
            .in1(N__31420),
            .in2(_gnd_net_),
            .in3(N__31403),
            .lcout(r_Clock_Count_0_adj_2454),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50529),
            .ce(),
            .sr(_gnd_net_));
    defparam i14960_3_lut_LC_10_29_0.C_ON=1'b0;
    defparam i14960_3_lut_LC_10_29_0.SEQ_MODE=4'b0000;
    defparam i14960_3_lut_LC_10_29_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 i14960_3_lut_LC_10_29_0 (
            .in0(N__32169),
            .in1(N__31377),
            .in2(_gnd_net_),
            .in3(N__32067),
            .lcout(n17398),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__0__2180_LC_10_29_1 .C_ON=1'b0;
    defparam \c0.data_out_8__0__2180_LC_10_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__0__2180_LC_10_29_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_out_8__0__2180_LC_10_29_1  (
            .in0(N__46855),
            .in1(N__46567),
            .in2(_gnd_net_),
            .in3(N__36271),
            .lcout(data_out_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50540),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i52_4_lut_LC_10_29_2 .C_ON=1'b0;
    defparam \c0.i52_4_lut_LC_10_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i52_4_lut_LC_10_29_2 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.i52_4_lut_LC_10_29_2  (
            .in0(N__32038),
            .in1(N__43149),
            .in2(N__34114),
            .in3(N__52457),
            .lcout(),
            .ltout(\c0.n29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i1_LC_10_29_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i1_LC_10_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i1_LC_10_29_3 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \c0.tx.r_Tx_Data_i1_LC_10_29_3  (
            .in0(N__35605),
            .in1(N__32082),
            .in2(N__32086),
            .in3(N__35520),
            .lcout(r_Tx_Data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50540),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i5_LC_10_29_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i5_LC_10_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i5_LC_10_29_4 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \c0.tx.r_Tx_Data_i5_LC_10_29_4  (
            .in0(N__35519),
            .in1(N__32068),
            .in2(N__35616),
            .in3(N__34093),
            .lcout(r_Tx_Data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50540),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15210_3_lut_LC_10_29_6 .C_ON=1'b0;
    defparam \c0.i15210_3_lut_LC_10_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15210_3_lut_LC_10_29_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \c0.i15210_3_lut_LC_10_29_6  (
            .in0(N__42701),
            .in1(N__40478),
            .in2(_gnd_net_),
            .in3(N__42467),
            .lcout(\c0.n17518 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_10_29_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_10_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_10_29_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_10_29_7  (
            .in0(N__33987),
            .in1(N__32059),
            .in2(_gnd_net_),
            .in3(N__52062),
            .lcout(\c0.n1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10915_2_lut_LC_10_30_0 .C_ON=1'b0;
    defparam \c0.i10915_2_lut_LC_10_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10915_2_lut_LC_10_30_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i10915_2_lut_LC_10_30_0  (
            .in0(_gnd_net_),
            .in1(N__39915),
            .in2(_gnd_net_),
            .in3(N__52042),
            .lcout(),
            .ltout(\c0.n9_adj_2143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i50_4_lut_LC_10_30_1 .C_ON=1'b0;
    defparam \c0.i50_4_lut_LC_10_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i50_4_lut_LC_10_30_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \c0.i50_4_lut_LC_10_30_1  (
            .in0(N__43147),
            .in1(N__32107),
            .in2(N__32041),
            .in3(N__52296),
            .lcout(\c0.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_10_30_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_10_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_10_30_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_10_30_2  (
            .in0(N__36820),
            .in1(N__39817),
            .in2(_gnd_net_),
            .in3(N__52040),
            .lcout(),
            .ltout(\c0.n5_adj_2326_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15562_LC_10_30_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15562_LC_10_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15562_LC_10_30_3 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15562_LC_10_30_3  (
            .in0(N__32032),
            .in1(N__52415),
            .in2(N__32020),
            .in3(N__52294),
            .lcout(\c0.n18023 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i7_LC_10_30_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i7_LC_10_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i7_LC_10_30_4 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \c0.tx.r_Tx_Data_i7_LC_10_30_4  (
            .in0(N__32170),
            .in1(N__32128),
            .in2(N__35524),
            .in3(N__35615),
            .lcout(r_Tx_Data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50549),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_10_30_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_10_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_10_30_6 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_10_30_6  (
            .in0(N__52295),
            .in1(N__40000),
            .in2(N__38128),
            .in3(N__52041),
            .lcout(n10_adj_2423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15344_2_lut_LC_10_30_7 .C_ON=1'b0;
    defparam \c0.i15344_2_lut_LC_10_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15344_2_lut_LC_10_30_7 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \c0.i15344_2_lut_LC_10_30_7  (
            .in0(N__52039),
            .in1(N__35290),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n17592 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__1__2243_LC_10_31_0 .C_ON=1'b0;
    defparam \c0.data_out_0__1__2243_LC_10_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__1__2243_LC_10_31_0 .LUT_INIT=16'b1010101000111010;
    LogicCell40 \c0.data_out_0__1__2243_LC_10_31_0  (
            .in0(N__32121),
            .in1(N__46421),
            .in2(N__45951),
            .in3(N__45536),
            .lcout(data_out_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50558),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18011_bdd_4_lut_LC_10_31_1 .C_ON=1'b0;
    defparam \c0.n18011_bdd_4_lut_LC_10_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18011_bdd_4_lut_LC_10_31_1 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n18011_bdd_4_lut_LC_10_31_1  (
            .in0(N__35260),
            .in1(N__34153),
            .in2(N__38146),
            .in3(N__52455),
            .lcout(\c0.n18014 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18041_bdd_4_lut_LC_10_31_4 .C_ON=1'b0;
    defparam \c0.n18041_bdd_4_lut_LC_10_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18041_bdd_4_lut_LC_10_31_4 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n18041_bdd_4_lut_LC_10_31_4  (
            .in0(N__52454),
            .in1(N__32485),
            .in2(N__32152),
            .in3(N__34168),
            .lcout(),
            .ltout(n18044_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_773_LC_10_31_5.C_ON=1'b0;
    defparam i24_4_lut_adj_773_LC_10_31_5.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_773_LC_10_31_5.LUT_INIT=16'b0011000010111000;
    LogicCell40 i24_4_lut_adj_773_LC_10_31_5 (
            .in0(N__32137),
            .in1(N__43119),
            .in2(N__32131),
            .in3(N__52456),
            .lcout(n10_adj_2414),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15336_3_lut_4_lut_LC_10_32_0 .C_ON=1'b0;
    defparam \c0.i15336_3_lut_4_lut_LC_10_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15336_3_lut_4_lut_LC_10_32_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.i15336_3_lut_4_lut_LC_10_32_0  (
            .in0(N__42603),
            .in1(N__40341),
            .in2(N__40195),
            .in3(N__40242),
            .lcout(\c0.n17445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18077_bdd_4_lut_LC_10_32_2 .C_ON=1'b0;
    defparam \c0.n18077_bdd_4_lut_LC_10_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18077_bdd_4_lut_LC_10_32_2 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n18077_bdd_4_lut_LC_10_32_2  (
            .in0(N__43146),
            .in1(N__35419),
            .in2(N__32122),
            .in3(N__40366),
            .lcout(\c0.n18080 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_10_32_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_10_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_10_32_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_10_32_4  (
            .in0(N__32097),
            .in1(N__38380),
            .in2(_gnd_net_),
            .in3(N__52060),
            .lcout(\c0.n2_adj_2137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__4__2232_LC_10_32_6 .C_ON=1'b0;
    defparam \c0.data_out_1__4__2232_LC_10_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__4__2232_LC_10_32_6 .LUT_INIT=16'b0011011100000100;
    LogicCell40 \c0.data_out_1__4__2232_LC_10_32_6  (
            .in0(N__46437),
            .in1(N__46139),
            .in2(N__42660),
            .in3(N__32479),
            .lcout(\c0.data_out_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50568),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i0_LC_11_17_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i0_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_state_i0_LC_11_17_1 .LUT_INIT=16'b1000111111001111;
    LogicCell40 \c0.FRAME_MATCHER_state_i0_LC_11_17_1  (
            .in0(N__34248),
            .in1(N__32467),
            .in2(N__32458),
            .in3(N__32419),
            .lcout(FRAME_MATCHER_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50429),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_418_LC_11_17_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_418_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_418_LC_11_17_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_418_LC_11_17_2  (
            .in0(N__32190),
            .in1(N__34246),
            .in2(_gnd_net_),
            .in3(N__32389),
            .lcout(\c0.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_405_LC_11_17_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_405_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_405_LC_11_17_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i1_2_lut_adj_405_LC_11_17_4  (
            .in0(N__32191),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32325),
            .lcout(\c0.n6_adj_2140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_654_LC_11_17_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_654_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_654_LC_11_17_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \c0.i1_2_lut_adj_654_LC_11_17_5  (
            .in0(N__32326),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33425),
            .lcout(),
            .ltout(\c0.n16814_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_663_LC_11_17_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_663_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_663_LC_11_17_6 .LUT_INIT=16'b1000000001000000;
    LogicCell40 \c0.i3_4_lut_adj_663_LC_11_17_6  (
            .in0(N__33533),
            .in1(N__32218),
            .in2(N__32206),
            .in3(N__34247),
            .lcout(\c0.n10052 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_3_lut_LC_11_17_7 .C_ON=1'b0;
    defparam \c0.tx2.i1_3_lut_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_3_lut_LC_11_17_7 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.tx2.i1_3_lut_LC_11_17_7  (
            .in0(N__51701),
            .in1(N__51535),
            .in2(_gnd_net_),
            .in3(N__47578),
            .lcout(\c0.tx2.n89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i31_LC_11_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i31_LC_11_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i31_LC_11_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i31_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__32194),
            .in2(_gnd_net_),
            .in3(N__34662),
            .lcout(\c0.FRAME_MATCHER_state_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50438),
            .ce(),
            .sr(N__33292));
    defparam \c0.FRAME_MATCHER_i_i0_LC_11_19_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i0_LC_11_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i0_LC_11_19_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i0_LC_11_19_0  (
            .in0(N__33208),
            .in1(N__32959),
            .in2(_gnd_net_),
            .in3(N__32725),
            .lcout(\c0.FRAME_MATCHER_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50444),
            .ce(),
            .sr(N__32626));
    defparam \c0.i15337_2_lut_LC_11_19_1 .C_ON=1'b0;
    defparam \c0.i15337_2_lut_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15337_2_lut_LC_11_19_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i15337_2_lut_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__35089),
            .in2(_gnd_net_),
            .in3(N__52080),
            .lcout(\c0.n17589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_717_LC_11_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_717_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_717_LC_11_19_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_717_LC_11_19_5  (
            .in0(N__34430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32588),
            .lcout(\c0.n16455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_723_LC_11_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_723_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_723_LC_11_19_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_723_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__32609),
            .in2(_gnd_net_),
            .in3(N__32589),
            .lcout(\c0.n16449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15485_LC_11_20_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15485_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15485_LC_11_20_0 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15485_LC_11_20_0  (
            .in0(N__48456),
            .in1(N__38848),
            .in2(N__32530),
            .in3(N__48207),
            .lcout(\c0.n17927 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15641_LC_11_20_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15641_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15641_LC_11_20_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15641_LC_11_20_1  (
            .in0(N__34849),
            .in1(N__51631),
            .in2(N__34369),
            .in3(N__47642),
            .lcout(),
            .ltout(\c0.n18119_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18119_bdd_4_lut_LC_11_20_2 .C_ON=1'b0;
    defparam \c0.n18119_bdd_4_lut_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18119_bdd_4_lut_LC_11_20_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18119_bdd_4_lut_LC_11_20_2  (
            .in0(N__51632),
            .in1(N__35830),
            .in2(N__32515),
            .in3(N__34855),
            .lcout(),
            .ltout(\c0.n18122_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i2_LC_11_20_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i2_LC_11_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i2_LC_11_20_3 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.tx2.r_Tx_Data_i2_LC_11_20_3  (
            .in0(N__34375),
            .in1(N__51763),
            .in2(N__32512),
            .in3(N__51633),
            .lcout(\c0.tx2.r_Tx_Data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50456),
            .ce(N__51451),
            .sr(_gnd_net_));
    defparam \c0.i14902_3_lut_LC_11_21_0 .C_ON=1'b0;
    defparam \c0.i14902_3_lut_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14902_3_lut_LC_11_21_0 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \c0.i14902_3_lut_LC_11_21_0  (
            .in0(N__40147),
            .in1(N__37430),
            .in2(_gnd_net_),
            .in3(N__35034),
            .lcout(\c0.n17340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11148_2_lut_3_lut_LC_11_21_2 .C_ON=1'b0;
    defparam \c0.i11148_2_lut_3_lut_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11148_2_lut_3_lut_LC_11_21_2 .LUT_INIT=16'b1111111011111110;
    LogicCell40 \c0.i11148_2_lut_3_lut_LC_11_21_2  (
            .in0(N__33358),
            .in1(N__33321),
            .in2(N__33433),
            .in3(_gnd_net_),
            .lcout(\c0.n13496 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_685_LC_11_21_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_685_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_685_LC_11_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_685_LC_11_21_3  (
            .in0(N__35810),
            .in1(N__35869),
            .in2(N__37116),
            .in3(N__40146),
            .lcout(\c0.n9919 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i60_LC_11_21_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i60_LC_11_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i60_LC_11_21_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \c0.data_out_frame2_0___i60_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(N__51147),
            .in2(N__33564),
            .in3(N__48844),
            .lcout(data_out_frame2_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50466),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_535_LC_11_21_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_535_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_535_LC_11_21_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_535_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(N__33557),
            .in2(_gnd_net_),
            .in3(N__36076),
            .lcout(\c0.n9916 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i52_LC_11_22_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i52_LC_11_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i52_LC_11_22_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i52_LC_11_22_0  (
            .in0(N__36736),
            .in1(N__34915),
            .in2(_gnd_net_),
            .in3(N__51277),
            .lcout(data_out_frame2_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50478),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15309_3_lut_LC_11_22_1 .C_ON=1'b0;
    defparam \c0.i15309_3_lut_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15309_3_lut_LC_11_22_1 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \c0.i15309_3_lut_LC_11_22_1  (
            .in0(N__48489),
            .in1(N__48065),
            .in2(_gnd_net_),
            .in3(N__37105),
            .lcout(\c0.n17579 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i98_LC_11_22_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i98_LC_11_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i98_LC_11_22_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i98_LC_11_22_2  (
            .in0(N__36249),
            .in1(N__41570),
            .in2(_gnd_net_),
            .in3(N__51278),
            .lcout(data_out_frame2_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50478),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_652_LC_11_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_652_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_652_LC_11_22_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i1_2_lut_adj_652_LC_11_22_3  (
            .in0(_gnd_net_),
            .in1(N__33532),
            .in2(_gnd_net_),
            .in3(N__33429),
            .lcout(),
            .ltout(\c0.n2_adj_2330_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_636_LC_11_22_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_636_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_636_LC_11_22_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_636_LC_11_22_4  (
            .in0(N__33357),
            .in1(N__33319),
            .in2(N__33295),
            .in3(N__34280),
            .lcout(\c0.n5545 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_527_LC_11_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_527_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_527_LC_11_22_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_527_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__35873),
            .in2(_gnd_net_),
            .in3(N__40152),
            .lcout(\c0.n16946 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_641_LC_11_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_641_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_641_LC_11_22_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_641_LC_11_22_6  (
            .in0(_gnd_net_),
            .in1(N__41569),
            .in2(_gnd_net_),
            .in3(N__47371),
            .lcout(\c0.n16963 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_488_LC_11_22_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_488_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_488_LC_11_22_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_488_LC_11_22_7  (
            .in0(N__49011),
            .in1(N__49743),
            .in2(N__43728),
            .in3(N__33586),
            .lcout(\c0.n17073 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_564_LC_11_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_564_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_564_LC_11_23_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_564_LC_11_23_0  (
            .in0(N__35063),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45362),
            .lcout(\c0.n9754 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15505_LC_11_23_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15505_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15505_LC_11_23_1 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15505_LC_11_23_1  (
            .in0(N__47231),
            .in1(N__48043),
            .in2(N__48564),
            .in3(N__36069),
            .lcout(\c0.n17951 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i130_LC_11_23_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i130_LC_11_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i130_LC_11_23_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i130_LC_11_23_3  (
            .in0(N__36245),
            .in1(N__39127),
            .in2(_gnd_net_),
            .in3(N__51276),
            .lcout(data_out_frame2_16_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50491),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i112_LC_11_23_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i112_LC_11_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i112_LC_11_23_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i112_LC_11_23_4  (
            .in0(N__51275),
            .in1(N__44012),
            .in2(_gnd_net_),
            .in3(N__43724),
            .lcout(data_out_frame2_13_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50491),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_694_LC_11_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_694_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_694_LC_11_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_694_LC_11_23_5  (
            .in0(N__35237),
            .in1(N__44345),
            .in2(_gnd_net_),
            .in3(N__41345),
            .lcout(\c0.n17091 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15465_LC_11_23_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15465_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15465_LC_11_23_6 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15465_LC_11_23_6  (
            .in0(N__48044),
            .in1(N__38779),
            .in2(N__49744),
            .in3(N__48465),
            .lcout(\c0.n17891 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_637_LC_11_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_637_LC_11_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_637_LC_11_23_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_637_LC_11_23_7  (
            .in0(N__35238),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44346),
            .lcout(\c0.n16936 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i145_LC_11_24_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i145_LC_11_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i145_LC_11_24_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_out_frame2_0___i145_LC_11_24_0  (
            .in0(N__34806),
            .in1(_gnd_net_),
            .in2(N__39547),
            .in3(N__51213),
            .lcout(data_out_frame2_18_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50501),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17987_bdd_4_lut_4_lut_LC_11_24_1 .C_ON=1'b0;
    defparam \c0.n17987_bdd_4_lut_4_lut_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.n17987_bdd_4_lut_4_lut_LC_11_24_1 .LUT_INIT=16'b1010101010011000;
    LogicCell40 \c0.n17987_bdd_4_lut_4_lut_LC_11_24_1  (
            .in0(N__39301),
            .in1(N__48224),
            .in2(N__35814),
            .in3(N__47712),
            .lcout(\c0.n17990 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15475_LC_11_24_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15475_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15475_LC_11_24_3 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15475_LC_11_24_3  (
            .in0(N__48578),
            .in1(N__48223),
            .in2(N__49469),
            .in3(N__47181),
            .lcout(\c0.n17915 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i97_LC_11_24_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i97_LC_11_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i97_LC_11_24_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i97_LC_11_24_4  (
            .in0(N__39545),
            .in1(N__47360),
            .in2(_gnd_net_),
            .in3(N__51214),
            .lcout(data_out_frame2_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50501),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i146_LC_11_24_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i146_LC_11_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i146_LC_11_24_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \c0.data_out_frame2_0___i146_LC_11_24_5  (
            .in0(_gnd_net_),
            .in1(N__51212),
            .in2(N__33643),
            .in3(N__36250),
            .lcout(data_out_frame2_18_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50501),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15470_LC_11_24_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15470_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15470_LC_11_24_6 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15470_LC_11_24_6  (
            .in0(N__48225),
            .in1(N__33639),
            .in2(N__49216),
            .in3(N__48579),
            .lcout(),
            .ltout(\c0.n17909_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17909_bdd_4_lut_LC_11_24_7 .C_ON=1'b0;
    defparam \c0.n17909_bdd_4_lut_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.n17909_bdd_4_lut_LC_11_24_7 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n17909_bdd_4_lut_LC_11_24_7  (
            .in0(N__39126),
            .in1(N__37867),
            .in2(N__33631),
            .in3(N__48493),
            .lcout(\c0.n17912 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18107_bdd_4_lut_LC_11_25_2 .C_ON=1'b0;
    defparam \c0.n18107_bdd_4_lut_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18107_bdd_4_lut_LC_11_25_2 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n18107_bdd_4_lut_LC_11_25_2  (
            .in0(N__33628),
            .in1(N__33619),
            .in2(N__33613),
            .in3(N__51645),
            .lcout(\c0.n18110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_11_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_11_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_11_25_4 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_11_25_4  (
            .in0(N__47815),
            .in1(N__33601),
            .in2(N__35908),
            .in3(N__47713),
            .lcout(),
            .ltout(\c0.n22_adj_2359_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i1_LC_11_25_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i1_LC_11_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i1_LC_11_25_5 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.tx2.r_Tx_Data_i1_LC_11_25_5  (
            .in0(N__51646),
            .in1(N__33595),
            .in2(N__33589),
            .in3(N__51762),
            .lcout(\c0.tx2.r_Tx_Data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50512),
            .ce(N__51404),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15567_LC_11_26_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15567_LC_11_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15567_LC_11_26_0 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15567_LC_11_26_0  (
            .in0(N__52451),
            .in1(N__33937),
            .in2(N__33895),
            .in3(N__52290),
            .lcout(),
            .ltout(\c0.n18029_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18029_bdd_4_lut_LC_11_26_1 .C_ON=1'b0;
    defparam \c0.n18029_bdd_4_lut_LC_11_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18029_bdd_4_lut_LC_11_26_1 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n18029_bdd_4_lut_LC_11_26_1  (
            .in0(N__33925),
            .in1(N__33916),
            .in2(N__33907),
            .in3(N__52452),
            .lcout(n18032),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_11_26_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_11_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_11_26_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_11_26_2  (
            .in0(N__40508),
            .in1(N__46856),
            .in2(_gnd_net_),
            .in3(N__52064),
            .lcout(\c0.n8_adj_2138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_15528_LC_11_26_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_15528_LC_11_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_15528_LC_11_26_5 .LUT_INIT=16'b1011110010110000;
    LogicCell40 \c0.byte_transmit_counter2_1__bdd_4_lut_15528_LC_11_26_5  (
            .in0(N__35143),
            .in1(N__47660),
            .in2(N__48629),
            .in3(N__36028),
            .lcout(\c0.n17897 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_11_26_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_11_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_11_26_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_11_26_6  (
            .in0(N__34141),
            .in1(N__46201),
            .in2(_gnd_net_),
            .in3(N__52063),
            .lcout(\c0.n5_adj_2299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__0__2172_LC_11_27_0 .C_ON=1'b0;
    defparam \c0.data_out_9__0__2172_LC_11_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__0__2172_LC_11_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_9__0__2172_LC_11_27_0  (
            .in0(N__39760),
            .in1(N__40087),
            .in2(_gnd_net_),
            .in3(N__37993),
            .lcout(\c0.data_out_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50530),
            .ce(N__46589),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__4__2160_LC_11_27_1 .C_ON=1'b0;
    defparam \c0.data_out_10__4__2160_LC_11_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__4__2160_LC_11_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_10__4__2160_LC_11_27_1  (
            .in0(N__38034),
            .in1(N__33958),
            .in2(_gnd_net_),
            .in3(N__35305),
            .lcout(\c0.data_out_10_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50530),
            .ce(N__46589),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_11_27_5 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_11_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_11_27_5 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_11_27_5  (
            .in0(N__33834),
            .in1(N__33790),
            .in2(_gnd_net_),
            .in3(N__33731),
            .lcout(n1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__2__2226_LC_11_28_0 .C_ON=1'b0;
    defparam \c0.data_out_2__2__2226_LC_11_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__2__2226_LC_11_28_0 .LUT_INIT=16'b1100110001011100;
    LogicCell40 \c0.data_out_2__2__2226_LC_11_28_0  (
            .in0(N__46485),
            .in1(N__35272),
            .in2(N__45990),
            .in3(N__45547),
            .lcout(data_out_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50541),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__5__2215_LC_11_28_1 .C_ON=1'b0;
    defparam \c0.data_out_3__5__2215_LC_11_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__5__2215_LC_11_28_1 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \c0.data_out_3__5__2215_LC_11_28_1  (
            .in0(N__45545),
            .in1(N__34036),
            .in2(N__45976),
            .in3(N__46487),
            .lcout(data_out_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50541),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__5__2223_LC_11_28_2 .C_ON=1'b0;
    defparam \c0.data_out_2__5__2223_LC_11_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__5__2223_LC_11_28_2 .LUT_INIT=16'b1101000111110000;
    LogicCell40 \c0.data_out_2__5__2223_LC_11_28_2  (
            .in0(N__46486),
            .in1(N__45546),
            .in2(N__34024),
            .in3(N__45911),
            .lcout(data_out_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50541),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_501_LC_11_28_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_501_LC_11_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_501_LC_11_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_501_LC_11_28_3  (
            .in0(N__46654),
            .in1(N__40504),
            .in2(N__34009),
            .in3(N__36827),
            .lcout(\c0.n10_adj_2276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_664_LC_11_28_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_664_LC_11_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_664_LC_11_28_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_664_LC_11_28_4  (
            .in0(N__34196),
            .in1(N__46853),
            .in2(N__39706),
            .in3(N__40408),
            .lcout(\c0.n16990 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__5__2183_LC_11_28_7 .C_ON=1'b0;
    defparam \c0.data_out_7__5__2183_LC_11_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__5__2183_LC_11_28_7 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \c0.data_out_7__5__2183_LC_11_28_7  (
            .in0(N__36514),
            .in1(N__34355),
            .in2(N__34140),
            .in3(N__42798),
            .lcout(\c0.data_out_7_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50541),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__6__2230_LC_11_29_0 .C_ON=1'b0;
    defparam \c0.data_out_1__6__2230_LC_11_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__6__2230_LC_11_29_0 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.data_out_1__6__2230_LC_11_29_0  (
            .in0(N__46447),
            .in1(N__45943),
            .in2(N__33991),
            .in3(N__45487),
            .lcout(data_out_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50550),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__0__2228_LC_11_29_3 .C_ON=1'b0;
    defparam \c0.data_out_2__0__2228_LC_11_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__0__2228_LC_11_29_3 .LUT_INIT=16'b1000110011011100;
    LogicCell40 \c0.data_out_2__0__2228_LC_11_29_3  (
            .in0(N__45486),
            .in1(N__33972),
            .in2(N__45989),
            .in3(N__46448),
            .lcout(data_out_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50550),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_550_LC_11_29_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_550_LC_11_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_550_LC_11_29_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_550_LC_11_29_4  (
            .in0(N__46854),
            .in1(N__34198),
            .in2(_gnd_net_),
            .in3(N__40414),
            .lcout(\c0.n9509 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__2__2170_LC_11_29_5 .C_ON=1'b0;
    defparam \c0.data_out_9__2__2170_LC_11_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__2__2170_LC_11_29_5 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \c0.data_out_9__2__2170_LC_11_29_5  (
            .in0(N__38097),
            .in1(N__37972),
            .in2(N__42761),
            .in3(N__42822),
            .lcout(data_out_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50550),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_544_LC_11_29_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_544_LC_11_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_544_LC_11_29_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_544_LC_11_29_6  (
            .in0(N__38025),
            .in1(N__34197),
            .in2(_gnd_net_),
            .in3(N__34133),
            .lcout(\c0.n9505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i53_4_lut_LC_11_29_7 .C_ON=1'b0;
    defparam \c0.i53_4_lut_LC_11_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i53_4_lut_LC_11_29_7 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \c0.i53_4_lut_LC_11_29_7  (
            .in0(N__45191),
            .in1(N__52289),
            .in2(N__34087),
            .in3(N__52061),
            .lcout(\c0.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__4__2184_LC_11_30_1 .C_ON=1'b0;
    defparam \c0.data_out_7__4__2184_LC_11_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__4__2184_LC_11_30_1 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \c0.data_out_7__4__2184_LC_11_30_1  (
            .in0(N__42864),
            .in1(N__34348),
            .in2(N__36828),
            .in3(N__36535),
            .lcout(\c0.data_out_7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50559),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_769_LC_11_30_2.C_ON=1'b0;
    defparam i24_4_lut_adj_769_LC_11_30_2.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_769_LC_11_30_2.LUT_INIT=16'b0010001011100010;
    LogicCell40 i24_4_lut_adj_769_LC_11_30_2 (
            .in0(N__34102),
            .in1(N__43148),
            .in2(N__39970),
            .in3(N__52405),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i5_3_lut_LC_11_30_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i5_3_lut_LC_11_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i5_3_lut_LC_11_30_3 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_1_i5_3_lut_LC_11_30_3  (
            .in0(N__40550),
            .in1(N__39705),
            .in2(N__52097),
            .in3(_gnd_net_),
            .lcout(\c0.n5_adj_2142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__0__2220_LC_11_30_4 .C_ON=1'b0;
    defparam \c0.data_out_3__0__2220_LC_11_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__0__2220_LC_11_30_4 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_out_3__0__2220_LC_11_30_4  (
            .in0(N__45492),
            .in1(N__42131),
            .in2(N__45988),
            .in3(N__34074),
            .lcout(data_out_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50559),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15297_2_lut_LC_11_30_5 .C_ON=1'b0;
    defparam \c0.i15297_2_lut_LC_11_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15297_2_lut_LC_11_30_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.i15297_2_lut_LC_11_30_5  (
            .in0(N__52076),
            .in1(N__34060),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n17588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15417_2_lut_3_lut_4_lut_LC_11_30_6 .C_ON=1'b0;
    defparam \c0.i15417_2_lut_3_lut_4_lut_LC_11_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15417_2_lut_3_lut_4_lut_LC_11_30_6 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \c0.i15417_2_lut_3_lut_4_lut_LC_11_30_6  (
            .in0(N__45491),
            .in1(N__42680),
            .in2(N__45987),
            .in3(N__46466),
            .lcout(\c0.n10054 ),
            .ltout(\c0.n10054_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__6__2182_LC_11_30_7 .C_ON=1'b0;
    defparam \c0.data_out_7__6__2182_LC_11_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__6__2182_LC_11_30_7 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \c0.data_out_7__6__2182_LC_11_30_7  (
            .in0(N__42865),
            .in1(N__36493),
            .in2(N__34039),
            .in3(N__38029),
            .lcout(\c0.data_out_7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50559),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_11_31_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_11_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_11_31_0 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_11_31_0  (
            .in0(_gnd_net_),
            .in1(N__52054),
            .in2(N__47049),
            .in3(N__46689),
            .lcout(\c0.n5_adj_2208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__7__2181_LC_11_31_1 .C_ON=1'b0;
    defparam \c0.data_out_7__7__2181_LC_11_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__7__2181_LC_11_31_1 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \c0.data_out_7__7__2181_LC_11_31_1  (
            .in0(N__36472),
            .in1(N__34195),
            .in2(N__34356),
            .in3(N__42863),
            .lcout(\c0.data_out_7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50569),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_11_31_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_11_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_11_31_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_11_31_2  (
            .in0(N__34194),
            .in1(N__52056),
            .in2(_gnd_net_),
            .in3(N__40270),
            .lcout(),
            .ltout(\c0.n5_adj_2188_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15616_LC_11_31_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15616_LC_11_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15616_LC_11_31_3 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15616_LC_11_31_3  (
            .in0(N__35668),
            .in1(N__52465),
            .in2(N__34171),
            .in3(N__52231),
            .lcout(\c0.n18041 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_522_LC_11_31_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_522_LC_11_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_522_LC_11_31_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_522_LC_11_31_4  (
            .in0(N__47045),
            .in1(N__42937),
            .in2(_gnd_net_),
            .in3(N__40241),
            .lcout(\c0.n16981 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15370_2_lut_LC_11_31_5 .C_ON=1'b0;
    defparam \c0.i15370_2_lut_LC_11_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15370_2_lut_LC_11_31_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15370_2_lut_LC_11_31_5  (
            .in0(N__52055),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40474),
            .lcout(),
            .ltout(\c0.n17543_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15552_LC_11_31_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15552_LC_11_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15552_LC_11_31_6 .LUT_INIT=16'b1101100010101010;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15552_LC_11_31_6  (
            .in0(N__52230),
            .in1(N__34162),
            .in2(N__34156),
            .in3(N__52453),
            .lcout(\c0.n18011 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__1__2187_LC_11_32_0 .C_ON=1'b0;
    defparam \c0.data_out_7__1__2187_LC_11_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__1__2187_LC_11_32_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \c0.data_out_7__1__2187_LC_11_32_0  (
            .in0(N__46434),
            .in1(N__45956),
            .in2(N__36319),
            .in3(N__34147),
            .lcout(\c0.data_out_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50577),
            .ce(N__34357),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__2__2186_LC_11_32_3 .C_ON=1'b0;
    defparam \c0.data_out_7__2__2186_LC_11_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__2__2186_LC_11_32_3 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \c0.data_out_7__2__2186_LC_11_32_3  (
            .in0(N__42725),
            .in1(N__40335),
            .in2(N__45640),
            .in3(N__46435),
            .lcout(\c0.data_out_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50577),
            .ce(N__34357),
            .sr(_gnd_net_));
    defparam \c0.i15208_2_lut_LC_11_32_4 .C_ON=1'b0;
    defparam \c0.i15208_2_lut_LC_11_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15208_2_lut_LC_11_32_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15208_2_lut_LC_11_32_4  (
            .in0(_gnd_net_),
            .in1(N__36562),
            .in2(_gnd_net_),
            .in3(N__45954),
            .lcout(),
            .ltout(\c0.n17456_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__3__2185_LC_11_32_5 .C_ON=1'b0;
    defparam \c0.data_out_7__3__2185_LC_11_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__3__2185_LC_11_32_5 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \c0.data_out_7__3__2185_LC_11_32_5  (
            .in0(N__42726),
            .in1(N__45069),
            .in2(N__34360),
            .in3(N__46436),
            .lcout(\c0.data_out_7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50577),
            .ce(N__34357),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__0__2188_LC_11_32_6 .C_ON=1'b0;
    defparam \c0.data_out_7__0__2188_LC_11_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__0__2188_LC_11_32_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \c0.data_out_7__0__2188_LC_11_32_6  (
            .in0(N__46433),
            .in1(N__45955),
            .in2(N__36346),
            .in3(N__40162),
            .lcout(\c0.data_out_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50577),
            .ce(N__34357),
            .sr(_gnd_net_));
    defparam i14716_2_lut_3_lut_LC_11_32_7.C_ON=1'b0;
    defparam i14716_2_lut_3_lut_LC_11_32_7.SEQ_MODE=4'b0000;
    defparam i14716_2_lut_3_lut_LC_11_32_7.LUT_INIT=16'b1111111110001000;
    LogicCell40 i14716_2_lut_3_lut_LC_11_32_7 (
            .in0(N__45953),
            .in1(N__46432),
            .in2(_gnd_net_),
            .in3(N__34321),
            .lcout(n17154),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i139_LC_12_16_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i139_LC_12_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i139_LC_12_16_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i139_LC_12_16_1  (
            .in0(N__36620),
            .in1(N__34392),
            .in2(_gnd_net_),
            .in3(N__51223),
            .lcout(data_out_frame2_17_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50445),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7942_2_lut_LC_12_17_3 .C_ON=1'b0;
    defparam \c0.i7942_2_lut_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7942_2_lut_LC_12_17_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i7942_2_lut_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__34683),
            .in2(_gnd_net_),
            .in3(N__34262),
            .lcout(\c0.n10297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2353__i0_LC_12_18_0 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2353__i0_LC_12_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2353__i0_LC_12_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2353__i0_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__34219),
            .in2(N__48096),
            .in3(_gnd_net_),
            .lcout(\c0.byte_transmit_counter2_0 ),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(\c0.n15615 ),
            .clk(N__50446),
            .ce(N__34690),
            .sr(N__34672));
    defparam \c0.byte_transmit_counter2_2353__i1_LC_12_18_1 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2353__i1_LC_12_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2353__i1_LC_12_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2353__i1_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(N__48354),
            .in2(_gnd_net_),
            .in3(N__34207),
            .lcout(\c0.byte_transmit_counter2_1 ),
            .ltout(),
            .carryin(\c0.n15615 ),
            .carryout(\c0.n15616 ),
            .clk(N__50446),
            .ce(N__34690),
            .sr(N__34672));
    defparam \c0.byte_transmit_counter2_2353__i2_LC_12_18_2 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2353__i2_LC_12_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2353__i2_LC_12_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2353__i2_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__47658),
            .in2(_gnd_net_),
            .in3(N__34204),
            .lcout(\c0.byte_transmit_counter2_2 ),
            .ltout(),
            .carryin(\c0.n15616 ),
            .carryout(\c0.n15617 ),
            .clk(N__50446),
            .ce(N__34690),
            .sr(N__34672));
    defparam \c0.byte_transmit_counter2_2353__i3_LC_12_18_3 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2353__i3_LC_12_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2353__i3_LC_12_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2353__i3_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__51576),
            .in2(_gnd_net_),
            .in3(N__34201),
            .lcout(\c0.byte_transmit_counter2_3 ),
            .ltout(),
            .carryin(\c0.n15617 ),
            .carryout(\c0.n15618 ),
            .clk(N__50446),
            .ce(N__34690),
            .sr(N__34672));
    defparam \c0.byte_transmit_counter2_2353__i4_LC_12_18_4 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2353__i4_LC_12_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2353__i4_LC_12_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2353__i4_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(N__51714),
            .in2(_gnd_net_),
            .in3(N__34759),
            .lcout(\c0.byte_transmit_counter2_4 ),
            .ltout(),
            .carryin(\c0.n15618 ),
            .carryout(\c0.n15619 ),
            .clk(N__50446),
            .ce(N__34690),
            .sr(N__34672));
    defparam \c0.byte_transmit_counter2_2353__i5_LC_12_18_5 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2353__i5_LC_12_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2353__i5_LC_12_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2353__i5_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(N__34752),
            .in2(_gnd_net_),
            .in3(N__34738),
            .lcout(\c0.byte_transmit_counter2_5 ),
            .ltout(),
            .carryin(\c0.n15619 ),
            .carryout(\c0.n15620 ),
            .clk(N__50446),
            .ce(N__34690),
            .sr(N__34672));
    defparam \c0.byte_transmit_counter2_2353__i6_LC_12_18_6 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2353__i6_LC_12_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2353__i6_LC_12_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2353__i6_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(N__34728),
            .in2(_gnd_net_),
            .in3(N__34714),
            .lcout(\c0.byte_transmit_counter2_6 ),
            .ltout(),
            .carryin(\c0.n15620 ),
            .carryout(\c0.n15621 ),
            .clk(N__50446),
            .ce(N__34690),
            .sr(N__34672));
    defparam \c0.byte_transmit_counter2_2353__i7_LC_12_18_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2353__i7_LC_12_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2353__i7_LC_12_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2353__i7_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(N__34704),
            .in2(_gnd_net_),
            .in3(N__34711),
            .lcout(\c0.byte_transmit_counter2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50446),
            .ce(N__34690),
            .sr(N__34672));
    defparam \c0.FRAME_MATCHER_state_i9_LC_12_19_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i9_LC_12_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i9_LC_12_19_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i9_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(N__34431),
            .in2(_gnd_net_),
            .in3(N__34651),
            .lcout(\c0.FRAME_MATCHER_state_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50457),
            .ce(),
            .sr(N__34411));
    defparam \c0.n17927_bdd_4_lut_LC_12_20_1 .C_ON=1'b0;
    defparam \c0.n17927_bdd_4_lut_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.n17927_bdd_4_lut_LC_12_20_1 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \c0.n17927_bdd_4_lut_LC_12_20_1  (
            .in0(N__48459),
            .in1(N__34405),
            .in2(N__34399),
            .in3(N__37043),
            .lcout(),
            .ltout(\c0.n17930_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_12_20_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_12_20_2 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_12_20_2  (
            .in0(N__47817),
            .in1(N__36919),
            .in2(N__34378),
            .in3(N__47645),
            .lcout(\c0.n22_adj_2358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17933_bdd_4_lut_LC_12_20_3 .C_ON=1'b0;
    defparam \c0.n17933_bdd_4_lut_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.n17933_bdd_4_lut_LC_12_20_3 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n17933_bdd_4_lut_LC_12_20_3  (
            .in0(N__48458),
            .in1(N__43380),
            .in2(N__49283),
            .in3(N__35971),
            .lcout(\c0.n17936 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_551_LC_12_20_5 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_551_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_551_LC_12_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_551_LC_12_20_5  (
            .in0(N__44646),
            .in1(N__36987),
            .in2(N__41968),
            .in3(N__39049),
            .lcout(\c0.n28_adj_2294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_12_20_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_12_20_6 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_12_20_6  (
            .in0(N__35959),
            .in1(N__48460),
            .in2(N__37672),
            .in3(N__48066),
            .lcout(\c0.n6_adj_2201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17939_bdd_4_lut_LC_12_20_7 .C_ON=1'b0;
    defparam \c0.n17939_bdd_4_lut_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.n17939_bdd_4_lut_LC_12_20_7 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \c0.n17939_bdd_4_lut_LC_12_20_7  (
            .in0(N__48457),
            .in1(N__34924),
            .in2(N__43908),
            .in3(N__38514),
            .lcout(\c0.n17942 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14863_4_lut_LC_12_21_1 .C_ON=1'b0;
    defparam \c0.i14863_4_lut_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14863_4_lut_LC_12_21_1 .LUT_INIT=16'b1100110001010000;
    LogicCell40 \c0.i14863_4_lut_LC_12_21_1  (
            .in0(N__48492),
            .in1(N__35779),
            .in2(N__34843),
            .in3(N__47643),
            .lcout(),
            .ltout(\c0.n17301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14865_3_lut_LC_12_21_2 .C_ON=1'b0;
    defparam \c0.i14865_3_lut_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14865_3_lut_LC_12_21_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \c0.i14865_3_lut_LC_12_21_2  (
            .in0(_gnd_net_),
            .in1(N__39229),
            .in2(N__34828),
            .in3(N__51617),
            .lcout(),
            .ltout(\c0.n17303_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i0_LC_12_21_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i0_LC_12_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i0_LC_12_21_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i0_LC_12_21_3  (
            .in0(N__51618),
            .in1(N__34765),
            .in2(N__34825),
            .in3(N__51739),
            .lcout(\c0.tx2.r_Tx_Data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50479),
            .ce(N__51452),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_12_21_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_12_21_4 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_LC_12_21_4  (
            .in0(N__34807),
            .in1(N__48490),
            .in2(N__36943),
            .in3(N__48052),
            .lcout(),
            .ltout(\c0.n18101_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18101_bdd_4_lut_LC_12_21_5 .C_ON=1'b0;
    defparam \c0.n18101_bdd_4_lut_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18101_bdd_4_lut_LC_12_21_5 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n18101_bdd_4_lut_LC_12_21_5  (
            .in0(N__48491),
            .in1(N__34792),
            .in2(N__34771),
            .in3(N__43847),
            .lcout(),
            .ltout(\c0.n18104_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_12_21_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_12_21_6 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_12_21_6  (
            .in0(N__47644),
            .in1(N__35884),
            .in2(N__34768),
            .in3(N__47816),
            .lcout(\c0.n22_adj_2337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_642_LC_12_22_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_642_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_642_LC_12_22_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_642_LC_12_22_0  (
            .in0(N__35167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43690),
            .lcout(\c0.n17106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15495_LC_12_22_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15495_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15495_LC_12_22_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15495_LC_12_22_1  (
            .in0(N__48051),
            .in1(N__40871),
            .in2(N__48580),
            .in3(N__35166),
            .lcout(\c0.n17939 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_4_lut_LC_12_22_2 .C_ON=1'b0;
    defparam \c0.i6_2_lut_4_lut_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_4_lut_LC_12_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_2_lut_4_lut_LC_12_22_2  (
            .in0(N__41344),
            .in1(N__40979),
            .in2(N__36756),
            .in3(N__39598),
            .lcout(\c0.n18_adj_2251 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_595_LC_12_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_595_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_595_LC_12_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_595_LC_12_22_3  (
            .in0(N__38522),
            .in1(N__34914),
            .in2(_gnd_net_),
            .in3(N__38580),
            .lcout(\c0.n17118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_626_LC_12_22_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_626_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_626_LC_12_22_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_626_LC_12_22_6  (
            .in0(N__43771),
            .in1(N__45367),
            .in2(N__37738),
            .in3(N__35062),
            .lcout(\c0.n17061 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_453_LC_12_22_7 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_453_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_453_LC_12_22_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_453_LC_12_22_7  (
            .in0(N__37304),
            .in1(N__41017),
            .in2(N__34891),
            .in3(N__34876),
            .lcout(\c0.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_451_LC_12_23_0 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_451_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_451_LC_12_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_451_LC_12_23_0  (
            .in0(N__41343),
            .in1(N__47224),
            .in2(N__44806),
            .in3(N__38752),
            .lcout(\c0.n22_adj_2194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_532_LC_12_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_532_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_532_LC_12_23_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_532_LC_12_23_1  (
            .in0(N__37303),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44282),
            .lcout(\c0.n9901 ),
            .ltout(\c0.n9901_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_473_LC_12_23_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_473_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_473_LC_12_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_473_LC_12_23_2  (
            .in0(N__34867),
            .in1(N__35874),
            .in2(N__34858),
            .in3(N__41704),
            .lcout(\c0.n19_adj_2254 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i122_LC_12_23_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i122_LC_12_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i122_LC_12_23_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i122_LC_12_23_3  (
            .in0(N__51196),
            .in1(N__37911),
            .in2(_gnd_net_),
            .in3(N__47188),
            .lcout(data_out_frame2_15_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50502),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i44_LC_12_23_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i44_LC_12_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i44_LC_12_23_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i44_LC_12_23_4  (
            .in0(N__37953),
            .in1(N__35064),
            .in2(_gnd_net_),
            .in3(N__51198),
            .lcout(data_out_frame2_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50502),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_526_LC_12_23_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_526_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_526_LC_12_23_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_526_LC_12_23_5  (
            .in0(N__47313),
            .in1(N__41238),
            .in2(N__38724),
            .in3(N__37606),
            .lcout(\c0.n9692 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_605_LC_12_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_605_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_605_LC_12_23_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_605_LC_12_23_6  (
            .in0(_gnd_net_),
            .in1(N__35159),
            .in2(_gnd_net_),
            .in3(N__43573),
            .lcout(\c0.n9707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i58_LC_12_23_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i58_LC_12_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i58_LC_12_23_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i58_LC_12_23_7  (
            .in0(N__51197),
            .in1(N__37912),
            .in2(_gnd_net_),
            .in3(N__38600),
            .lcout(data_out_frame2_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50502),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14893_3_lut_LC_12_24_0 .C_ON=1'b0;
    defparam \c0.i14893_3_lut_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14893_3_lut_LC_12_24_0 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \c0.i14893_3_lut_LC_12_24_0  (
            .in0(N__48694),
            .in1(N__37454),
            .in2(_gnd_net_),
            .in3(N__35038),
            .lcout(),
            .ltout(\c0.n17331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i7_LC_12_24_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i7_LC_12_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i7_LC_12_24_1 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.data_out_frame2_0___i7_LC_12_24_1  (
            .in0(N__37455),
            .in1(N__37552),
            .in2(N__34981),
            .in3(N__34976),
            .lcout(\c0.data_out_frame2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50513),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17891_bdd_4_lut_LC_12_24_2 .C_ON=1'b0;
    defparam \c0.n17891_bdd_4_lut_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.n17891_bdd_4_lut_LC_12_24_2 .LUT_INIT=16'b1010101011100100;
    LogicCell40 \c0.n17891_bdd_4_lut_LC_12_24_2  (
            .in0(N__34930),
            .in1(N__37731),
            .in2(N__45256),
            .in3(N__48391),
            .lcout(\c0.n17894 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i129_LC_12_24_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i129_LC_12_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i129_LC_12_24_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.data_out_frame2_0___i129_LC_12_24_3  (
            .in0(_gnd_net_),
            .in1(N__51073),
            .in2(N__39533),
            .in3(N__43831),
            .lcout(data_out_frame2_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50513),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i125_LC_12_24_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i125_LC_12_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i125_LC_12_24_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i125_LC_12_24_4  (
            .in0(N__37767),
            .in1(N__44160),
            .in2(_gnd_net_),
            .in3(N__51211),
            .lcout(data_out_frame2_15_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50513),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i83_LC_12_24_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i83_LC_12_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i83_LC_12_24_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i83_LC_12_24_5  (
            .in0(N__51210),
            .in1(N__44487),
            .in2(_gnd_net_),
            .in3(N__35165),
            .lcout(data_out_frame2_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50513),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i12_3_lut_LC_12_24_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i12_3_lut_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i12_3_lut_LC_12_24_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i12_3_lut_LC_12_24_6  (
            .in0(N__37580),
            .in1(N__47962),
            .in2(_gnd_net_),
            .in3(N__37756),
            .lcout(\c0.n12_adj_2305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11219217_i1_3_lut_LC_12_24_7 .C_ON=1'b0;
    defparam \c0.i11219217_i1_3_lut_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i11219217_i1_3_lut_LC_12_24_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.i11219217_i1_3_lut_LC_12_24_7  (
            .in0(N__35134),
            .in1(N__35404),
            .in2(_gnd_net_),
            .in3(N__51613),
            .lcout(\c0.n15_adj_2356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15538_LC_12_25_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15538_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15538_LC_12_25_2 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15538_LC_12_25_2  (
            .in0(N__47963),
            .in1(N__48392),
            .in2(N__38570),
            .in3(N__41140),
            .lcout(),
            .ltout(\c0.n17993_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17993_bdd_4_lut_LC_12_25_3 .C_ON=1'b0;
    defparam \c0.n17993_bdd_4_lut_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.n17993_bdd_4_lut_LC_12_25_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n17993_bdd_4_lut_LC_12_25_3  (
            .in0(N__48393),
            .in1(N__41868),
            .in2(N__35128),
            .in3(N__44854),
            .lcout(),
            .ltout(\c0.n17393_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15606_LC_12_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15606_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15606_LC_12_25_4 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15606_LC_12_25_4  (
            .in0(N__35125),
            .in1(N__51614),
            .in2(N__35119),
            .in3(N__47631),
            .lcout(),
            .ltout(\c0.n17963_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17963_bdd_4_lut_LC_12_25_5 .C_ON=1'b0;
    defparam \c0.n17963_bdd_4_lut_LC_12_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.n17963_bdd_4_lut_LC_12_25_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n17963_bdd_4_lut_LC_12_25_5  (
            .in0(N__51615),
            .in1(N__35116),
            .in2(N__35107),
            .in3(N__44581),
            .lcout(),
            .ltout(\c0.n17966_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i5_LC_12_25_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i5_LC_12_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i5_LC_12_25_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \c0.tx2.r_Tx_Data_i5_LC_12_25_6  (
            .in0(N__51761),
            .in1(N__51616),
            .in2(N__35104),
            .in3(N__36115),
            .lcout(\c0.tx2.r_Tx_Data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50521),
            .ce(N__51411),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__5__2239_LC_12_26_0 .C_ON=1'b0;
    defparam \c0.data_out_0__5__2239_LC_12_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__5__2239_LC_12_26_0 .LUT_INIT=16'b1111101100001000;
    LogicCell40 \c0.data_out_0__5__2239_LC_12_26_0  (
            .in0(N__42156),
            .in1(N__45978),
            .in2(N__45537),
            .in3(N__35085),
            .lcout(data_out_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50531),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i66_LC_12_26_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i66_LC_12_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i66_LC_12_26_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i66_LC_12_26_1  (
            .in0(N__36231),
            .in1(N__47270),
            .in2(_gnd_net_),
            .in3(N__51178),
            .lcout(data_out_frame2_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50531),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i86_LC_12_26_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i86_LC_12_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i86_LC_12_26_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i86_LC_12_26_3  (
            .in0(N__40619),
            .in1(N__38569),
            .in2(_gnd_net_),
            .in3(N__51179),
            .lcout(data_out_frame2_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50531),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i9_3_lut_LC_12_26_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i9_3_lut_LC_12_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i9_3_lut_LC_12_26_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i9_3_lut_LC_12_26_4  (
            .in0(N__37838),
            .in1(N__48107),
            .in2(_gnd_net_),
            .in3(N__42072),
            .lcout(\c0.n9_adj_2347 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__3__2241_LC_12_26_5 .C_ON=1'b0;
    defparam \c0.data_out_0__3__2241_LC_12_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__3__2241_LC_12_26_5 .LUT_INIT=16'b1000110011011100;
    LogicCell40 \c0.data_out_0__3__2241_LC_12_26_5  (
            .in0(N__45510),
            .in1(N__35286),
            .in2(N__45999),
            .in3(N__46492),
            .lcout(data_out_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50531),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i149_LC_12_26_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i149_LC_12_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i149_LC_12_26_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i149_LC_12_26_7  (
            .in0(N__37348),
            .in1(N__37236),
            .in2(_gnd_net_),
            .in3(N__51177),
            .lcout(data_out_frame2_18_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50531),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_27_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_27_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_27_0  (
            .in0(N__35247),
            .in1(N__52065),
            .in2(_gnd_net_),
            .in3(N__35271),
            .lcout(\c0.n2_adj_2291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15249_3_lut_LC_12_27_2 .C_ON=1'b0;
    defparam \c0.i15249_3_lut_LC_12_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15249_3_lut_LC_12_27_2 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \c0.i15249_3_lut_LC_12_27_2  (
            .in0(N__45206),
            .in1(N__42752),
            .in2(_gnd_net_),
            .in3(N__40480),
            .lcout(\c0.n17514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__2__2218_LC_12_27_4 .C_ON=1'b0;
    defparam \c0.data_out_3__2__2218_LC_12_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__2__2218_LC_12_27_4 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.data_out_3__2__2218_LC_12_27_4  (
            .in0(N__35248),
            .in1(N__45977),
            .in2(N__42155),
            .in3(N__45514),
            .lcout(data_out_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50542),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i8_3_lut_LC_12_27_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i8_3_lut_LC_12_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i8_3_lut_LC_12_27_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i8_3_lut_LC_12_27_6  (
            .in0(N__48121),
            .in1(N__35236),
            .in2(_gnd_net_),
            .in3(N__49343),
            .lcout(),
            .ltout(\c0.n8_adj_2348_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17897_bdd_4_lut_LC_12_27_7 .C_ON=1'b0;
    defparam \c0.n17897_bdd_4_lut_LC_12_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.n17897_bdd_4_lut_LC_12_27_7 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n17897_bdd_4_lut_LC_12_27_7  (
            .in0(N__35185),
            .in1(N__35173),
            .in2(N__35407),
            .in3(N__47632),
            .lcout(\c0.n17900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4030_2_lut_LC_12_28_0 .C_ON=1'b0;
    defparam \c0.i4030_2_lut_LC_12_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4030_2_lut_LC_12_28_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i4030_2_lut_LC_12_28_0  (
            .in0(_gnd_net_),
            .in1(N__45936),
            .in2(_gnd_net_),
            .in3(N__46481),
            .lcout(n2547),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_667_LC_12_28_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_667_LC_12_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_667_LC_12_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_667_LC_12_28_2  (
            .in0(N__47139),
            .in1(N__52511),
            .in2(N__46702),
            .in3(N__39786),
            .lcout(\c0.n16975 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_15631_LC_12_28_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_15631_LC_12_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_15631_LC_12_28_5 .LUT_INIT=16'b1100111110100000;
    LogicCell40 \c0.tx2.r_Bit_Index_0__bdd_4_lut_15631_LC_12_28_5  (
            .in0(N__47530),
            .in1(N__45565),
            .in2(N__35392),
            .in3(N__35350),
            .lcout(\c0.tx2.n17903 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_643_LC_12_28_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_643_LC_12_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_643_LC_12_28_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_643_LC_12_28_7  (
            .in0(N__43011),
            .in1(N__39877),
            .in2(_gnd_net_),
            .in3(N__40412),
            .lcout(\c0.n32_adj_2297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__3__2177_LC_12_29_0 .C_ON=1'b0;
    defparam \c0.data_out_8__3__2177_LC_12_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__3__2177_LC_12_29_0 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_out_8__3__2177_LC_12_29_0  (
            .in0(N__42753),
            .in1(N__36390),
            .in2(N__42861),
            .in3(N__43012),
            .lcout(\c0.data_out_8_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50560),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_683_LC_12_29_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_683_LC_12_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_683_LC_12_29_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_683_LC_12_29_1  (
            .in0(N__42284),
            .in1(N__38101),
            .in2(_gnd_net_),
            .in3(N__42400),
            .lcout(\c0.n17055 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_539_LC_12_29_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_539_LC_12_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_539_LC_12_29_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_539_LC_12_29_2  (
            .in0(N__38102),
            .in1(N__46804),
            .in2(_gnd_net_),
            .in3(N__46898),
            .lcout(),
            .ltout(\c0.n16978_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_507_LC_12_29_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_507_LC_12_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_507_LC_12_29_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_507_LC_12_29_3  (
            .in0(N__35304),
            .in1(N__35659),
            .in2(N__35293),
            .in3(N__46719),
            .lcout(\c0.n20_adj_2282 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__4__2176_LC_12_29_5 .C_ON=1'b0;
    defparam \c0.data_out_8__4__2176_LC_12_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__4__2176_LC_12_29_5 .LUT_INIT=16'b1111101100001000;
    LogicCell40 \c0.data_out_8__4__2176_LC_12_29_5  (
            .in0(N__36372),
            .in1(N__42843),
            .in2(N__42762),
            .in3(N__42958),
            .lcout(data_out_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50560),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_689_LC_12_29_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_689_LC_12_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_689_LC_12_29_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_689_LC_12_29_7  (
            .in0(_gnd_net_),
            .in1(N__35701),
            .in2(_gnd_net_),
            .in3(N__42957),
            .lcout(\c0.n9728 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_499_LC_12_30_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_499_LC_12_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_499_LC_12_30_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_499_LC_12_30_0  (
            .in0(N__45114),
            .in1(N__42469),
            .in2(N__40524),
            .in3(N__42936),
            .lcout(\c0.n16969 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_513_LC_12_30_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_513_LC_12_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_513_LC_12_30_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_513_LC_12_30_1  (
            .in0(_gnd_net_),
            .in1(N__40336),
            .in2(_gnd_net_),
            .in3(N__45070),
            .lcout(\c0.n16912 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_3_lut_LC_12_30_3 .C_ON=1'b0;
    defparam \c0.i22_3_lut_LC_12_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i22_3_lut_LC_12_30_3 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.i22_3_lut_LC_12_30_3  (
            .in0(N__38096),
            .in1(N__39871),
            .in2(N__52098),
            .in3(_gnd_net_),
            .lcout(\c0.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18035_bdd_4_lut_LC_12_30_4 .C_ON=1'b0;
    defparam \c0.n18035_bdd_4_lut_LC_12_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18035_bdd_4_lut_LC_12_30_4 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n18035_bdd_4_lut_LC_12_30_4  (
            .in0(N__35641),
            .in1(N__35677),
            .in2(N__35635),
            .in3(N__52406),
            .lcout(),
            .ltout(n18038_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_771_LC_12_30_5.C_ON=1'b0;
    defparam i24_4_lut_adj_771_LC_12_30_5.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_771_LC_12_30_5.LUT_INIT=16'b0100010011110000;
    LogicCell40 i24_4_lut_adj_771_LC_12_30_5 (
            .in0(N__52407),
            .in1(N__38191),
            .in2(N__35620),
            .in3(N__43153),
            .lcout(),
            .ltout(n10_adj_2413_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i6_LC_12_30_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i6_LC_12_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i6_LC_12_30_6 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \c0.tx.r_Tx_Data_i6_LC_12_30_6  (
            .in0(N__35602),
            .in1(N__35433),
            .in2(N__35527),
            .in3(N__35523),
            .lcout(r_Tx_Data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50570),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__1__2203_LC_12_31_0 .C_ON=1'b0;
    defparam \c0.data_out_5__1__2203_LC_12_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__1__2203_LC_12_31_0 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \c0.data_out_5__1__2203_LC_12_31_0  (
            .in0(N__46403),
            .in1(N__45785),
            .in2(N__42751),
            .in3(N__36645),
            .lcout(\c0.data_out_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50578),
            .ce(N__46131),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__1__2235_LC_12_31_2 .C_ON=1'b0;
    defparam \c0.data_out_1__1__2235_LC_12_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__1__2235_LC_12_31_2 .LUT_INIT=16'b1000110110001101;
    LogicCell40 \c0.data_out_1__1__2235_LC_12_31_2  (
            .in0(N__46402),
            .in1(N__45784),
            .in2(N__42750),
            .in3(_gnd_net_),
            .lcout(\c0.data_out_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50578),
            .ce(N__46131),
            .sr(_gnd_net_));
    defparam \c0.mux_1210_i1_3_lut_LC_12_31_3 .C_ON=1'b0;
    defparam \c0.mux_1210_i1_3_lut_LC_12_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.mux_1210_i1_3_lut_LC_12_31_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.mux_1210_i1_3_lut_LC_12_31_3  (
            .in0(N__45782),
            .in1(N__42712),
            .in2(_gnd_net_),
            .in3(N__46401),
            .lcout(n2652),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_LC_12_31_5 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_LC_12_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_LC_12_31_5 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \c0.i6_2_lut_3_lut_LC_12_31_5  (
            .in0(N__45781),
            .in1(N__42711),
            .in2(_gnd_net_),
            .in3(N__46400),
            .lcout(\c0.n10181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__6__2190_LC_12_31_7 .C_ON=1'b0;
    defparam \c0.data_out_6__6__2190_LC_12_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__6__2190_LC_12_31_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_6__6__2190_LC_12_31_7  (
            .in0(N__45783),
            .in1(N__36669),
            .in2(N__37789),
            .in3(N__46404),
            .lcout(\c0.data_out_6_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50578),
            .ce(N__46131),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_12_32_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_12_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_12_32_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_12_32_0  (
            .in0(N__38033),
            .in1(N__35700),
            .in2(_gnd_net_),
            .in3(N__52071),
            .lcout(\c0.n5_adj_2300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15362_2_lut_LC_12_32_1 .C_ON=1'b0;
    defparam \c0.i15362_2_lut_LC_12_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15362_2_lut_LC_12_32_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15362_2_lut_LC_12_32_1  (
            .in0(N__52072),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40322),
            .lcout(),
            .ltout(\c0.n17555_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15572_LC_12_32_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15572_LC_12_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15572_LC_12_32_2 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15572_LC_12_32_2  (
            .in0(N__35686),
            .in1(N__52464),
            .in2(N__35680),
            .in3(N__52303),
            .lcout(\c0.n18035 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__6__2198_LC_12_32_3 .C_ON=1'b0;
    defparam \c0.data_out_5__6__2198_LC_12_32_3 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__6__2198_LC_12_32_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.data_out_5__6__2198_LC_12_32_3  (
            .in0(_gnd_net_),
            .in1(N__36870),
            .in2(_gnd_net_),
            .in3(N__45997),
            .lcout(\c0.data_out_7__2__N_447 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50584),
            .ce(N__46137),
            .sr(N__41896));
    defparam \c0.data_out_5__7__2197_LC_12_32_5 .C_ON=1'b0;
    defparam \c0.data_out_5__7__2197_LC_12_32_5 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__7__2197_LC_12_32_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.data_out_5__7__2197_LC_12_32_5  (
            .in0(_gnd_net_),
            .in1(N__36849),
            .in2(_gnd_net_),
            .in3(N__45998),
            .lcout(\c0.data_out_7__3__N_441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50584),
            .ce(N__46137),
            .sr(N__41896));
    defparam \c0.i15281_2_lut_LC_12_32_6 .C_ON=1'b0;
    defparam \c0.i15281_2_lut_LC_12_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15281_2_lut_LC_12_32_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15281_2_lut_LC_12_32_6  (
            .in0(_gnd_net_),
            .in1(N__45057),
            .in2(_gnd_net_),
            .in3(N__52070),
            .lcout(\c0.n17569 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_645_LC_13_18_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_645_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_645_LC_13_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_645_LC_13_18_1  (
            .in0(N__36961),
            .in1(N__40875),
            .in2(N__35941),
            .in3(N__43584),
            .lcout(\c0.n20_adj_2333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15324_2_lut_3_lut_LC_13_18_4 .C_ON=1'b0;
    defparam \c0.i15324_2_lut_3_lut_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15324_2_lut_3_lut_LC_13_18_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \c0.i15324_2_lut_3_lut_LC_13_18_4  (
            .in0(N__35875),
            .in1(N__48353),
            .in2(_gnd_net_),
            .in3(N__48009),
            .lcout(\c0.n17578 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_470_LC_13_19_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_470_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_470_LC_13_19_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_470_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__40978),
            .in2(_gnd_net_),
            .in3(N__39597),
            .lcout(\c0.n17121 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_572_LC_13_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_572_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_572_LC_13_19_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_572_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__43651),
            .in2(_gnd_net_),
            .in3(N__40803),
            .lcout(\c0.n9810 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_630_LC_13_19_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_630_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_630_LC_13_19_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_630_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__43464),
            .in2(_gnd_net_),
            .in3(N__37148),
            .lcout(\c0.n9859 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i67_LC_13_19_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i67_LC_13_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i67_LC_13_19_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i67_LC_13_19_7  (
            .in0(N__36441),
            .in1(N__38518),
            .in2(_gnd_net_),
            .in3(N__51183),
            .lcout(data_out_frame2_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50467),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_450_LC_13_20_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_450_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_450_LC_13_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_450_LC_13_20_0  (
            .in0(N__35818),
            .in1(N__37587),
            .in2(_gnd_net_),
            .in3(N__37771),
            .lcout(\c0.n17124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i131_LC_13_20_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i131_LC_13_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i131_LC_13_20_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i131_LC_13_20_1  (
            .in0(N__36439),
            .in1(N__37053),
            .in2(_gnd_net_),
            .in3(N__51136),
            .lcout(data_out_frame2_16_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50480),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i99_LC_13_20_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i99_LC_13_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i99_LC_13_20_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i99_LC_13_20_2  (
            .in0(N__51135),
            .in1(N__36440),
            .in2(_gnd_net_),
            .in3(N__49272),
            .lcout(data_out_frame2_12_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50480),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_13_20_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_13_20_3 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_13_20_3  (
            .in0(N__47961),
            .in1(N__48513),
            .in2(N__37126),
            .in3(N__44737),
            .lcout(\c0.n6_adj_2335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_13_20_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_13_20_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_13_20_4  (
            .in0(N__40977),
            .in1(N__47960),
            .in2(_gnd_net_),
            .in3(N__44442),
            .lcout(\c0.n5_adj_2317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i49_LC_13_20_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i49_LC_13_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i49_LC_13_20_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i49_LC_13_20_5  (
            .in0(N__41755),
            .in1(N__37150),
            .in2(_gnd_net_),
            .in3(N__51137),
            .lcout(data_out_frame2_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50480),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_486_LC_13_20_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_486_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_486_LC_13_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_486_LC_13_20_6  (
            .in0(N__49702),
            .in1(N__43902),
            .in2(N__38470),
            .in3(N__35950),
            .lcout(\c0.n15_adj_2269 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i76_LC_13_20_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i76_LC_13_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i76_LC_13_20_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i76_LC_13_20_7  (
            .in0(N__37957),
            .in1(N__37302),
            .in2(_gnd_net_),
            .in3(N__51138),
            .lcout(data_out_frame2_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50480),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_624_LC_13_21_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_624_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_624_LC_13_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_624_LC_13_21_1  (
            .in0(N__37847),
            .in1(N__49271),
            .in2(N__37668),
            .in3(N__43646),
            .lcout(\c0.n16957 ),
            .ltout(\c0.n16957_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_570_LC_13_21_2 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_570_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_570_LC_13_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_570_LC_13_21_2  (
            .in0(N__35937),
            .in1(N__35892),
            .in2(N__35917),
            .in3(N__37693),
            .lcout(\c0.n21_adj_2304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i162_LC_13_21_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i162_LC_13_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i162_LC_13_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i162_LC_13_21_3  (
            .in0(N__35914),
            .in1(N__41938),
            .in2(N__36892),
            .in3(N__37060),
            .lcout(\c0.data_out_frame2_20_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50492),
            .ce(N__51184),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i161_LC_13_21_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i161_LC_13_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i161_LC_13_21_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.data_out_frame2_0___i161_LC_13_21_5  (
            .in0(N__35893),
            .in1(N__38683),
            .in2(_gnd_net_),
            .in3(N__40828),
            .lcout(\c0.data_out_frame2_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50492),
            .ce(N__51184),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_562_LC_13_21_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_562_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_562_LC_13_21_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_562_LC_13_21_6  (
            .in0(_gnd_net_),
            .in1(N__37664),
            .in2(_gnd_net_),
            .in3(N__37848),
            .lcout(\c0.n9886 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_448_LC_13_22_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_448_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_448_LC_13_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_448_LC_13_22_1  (
            .in0(N__43477),
            .in1(N__49431),
            .in2(N__41067),
            .in3(N__36016),
            .lcout(),
            .ltout(\c0.n16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i167_LC_13_22_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i167_LC_13_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i167_LC_13_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i167_LC_13_22_2  (
            .in0(N__36007),
            .in1(N__37081),
            .in2(N__35995),
            .in3(N__36967),
            .lcout(\c0.data_out_frame2_20_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50503),
            .ce(N__50965),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_696_LC_13_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_696_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_696_LC_13_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_696_LC_13_22_3  (
            .in0(N__44284),
            .in1(N__37736),
            .in2(_gnd_net_),
            .in3(N__49007),
            .lcout(\c0.n17112 ),
            .ltout(\c0.n17112_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_580_LC_13_22_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_580_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_580_LC_13_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_580_LC_13_22_4  (
            .in0(N__38664),
            .in1(N__38455),
            .in2(N__35992),
            .in3(N__39403),
            .lcout(),
            .ltout(\c0.n14_adj_2308_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i158_LC_13_22_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i158_LC_13_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i158_LC_13_22_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i158_LC_13_22_5  (
            .in0(N__38545),
            .in1(N__37165),
            .in2(N__35989),
            .in3(N__47415),
            .lcout(\c0.data_out_frame2_19_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50503),
            .ce(N__50965),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_620_LC_13_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_620_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_620_LC_13_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_620_LC_13_22_6  (
            .in0(N__37652),
            .in1(N__43647),
            .in2(_gnd_net_),
            .in3(N__40782),
            .lcout(\c0.n17067 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i63_LC_13_23_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i63_LC_13_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i63_LC_13_23_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i63_LC_13_23_0  (
            .in0(N__50939),
            .in1(N__49106),
            .in2(_gnd_net_),
            .in3(N__44354),
            .lcout(data_out_frame2_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50514),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15490_LC_13_23_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15490_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15490_LC_13_23_1 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15490_LC_13_23_1  (
            .in0(N__48584),
            .in1(N__48042),
            .in2(N__39159),
            .in3(N__39589),
            .lcout(\c0.n17933 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i116_LC_13_23_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i116_LC_13_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i116_LC_13_23_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i116_LC_13_23_2  (
            .in0(N__50937),
            .in1(_gnd_net_),
            .in2(N__36735),
            .in3(N__47237),
            .lcout(data_out_frame2_14_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50514),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i111_LC_13_23_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i111_LC_13_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i111_LC_13_23_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i111_LC_13_23_3  (
            .in0(N__48935),
            .in1(N__49651),
            .in2(_gnd_net_),
            .in3(N__50941),
            .lcout(data_out_frame2_13_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50514),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_518_LC_13_23_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_518_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_518_LC_13_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_518_LC_13_23_4  (
            .in0(N__39334),
            .in1(N__37594),
            .in2(N__49658),
            .in3(N__37206),
            .lcout(\c0.n17133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_588_LC_13_23_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_588_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_588_LC_13_23_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_588_LC_13_23_5  (
            .in0(N__40717),
            .in1(N__36075),
            .in2(N__44736),
            .in3(N__39014),
            .lcout(\c0.n9865 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i59_LC_13_23_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i59_LC_13_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i59_LC_13_23_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i59_LC_13_23_6  (
            .in0(N__50938),
            .in1(_gnd_net_),
            .in2(N__36621),
            .in3(N__40983),
            .lcout(data_out_frame2_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50514),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i109_LC_13_23_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i109_LC_13_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i109_LC_13_23_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i109_LC_13_23_7  (
            .in0(N__39203),
            .in1(N__36043),
            .in2(_gnd_net_),
            .in3(N__50940),
            .lcout(data_out_frame2_13_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50514),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_589_LC_13_24_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_589_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_589_LC_13_24_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_589_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__39151),
            .in2(_gnd_net_),
            .in3(N__36042),
            .lcout(\c0.n9814 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i11_3_lut_LC_13_24_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i11_3_lut_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i11_3_lut_LC_13_24_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i11_3_lut_LC_13_24_1  (
            .in0(N__36041),
            .in1(N__38439),
            .in2(_gnd_net_),
            .in3(N__48030),
            .lcout(\c0.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i101_LC_13_24_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i101_LC_13_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i101_LC_13_24_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_out_frame2_0___i101_LC_13_24_2  (
            .in0(N__38440),
            .in1(_gnd_net_),
            .in2(N__37353),
            .in3(N__50923),
            .lcout(data_out_frame2_12_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50522),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i133_LC_13_24_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i133_LC_13_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i133_LC_13_24_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i133_LC_13_24_3  (
            .in0(N__50921),
            .in1(N__37344),
            .in2(_gnd_net_),
            .in3(N__40781),
            .lcout(data_out_frame2_16_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50522),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i123_LC_13_24_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i123_LC_13_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i123_LC_13_24_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i123_LC_13_24_4  (
            .in0(N__36619),
            .in1(N__39152),
            .in2(_gnd_net_),
            .in3(N__50924),
            .lcout(data_out_frame2_15_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50522),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17981_bdd_4_lut_LC_13_24_5 .C_ON=1'b0;
    defparam \c0.n17981_bdd_4_lut_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.n17981_bdd_4_lut_LC_13_24_5 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \c0.n17981_bdd_4_lut_LC_13_24_5  (
            .in0(N__36130),
            .in1(N__48586),
            .in2(N__36108),
            .in3(N__41406),
            .lcout(),
            .ltout(\c0.n17984_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_13_24_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_13_24_6 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_13_24_6  (
            .in0(N__38905),
            .in1(N__47804),
            .in2(N__36118),
            .in3(N__47706),
            .lcout(\c0.n22_adj_2354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i142_LC_13_24_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i142_LC_13_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i142_LC_13_24_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_out_frame2_0___i142_LC_13_24_7  (
            .in0(N__50922),
            .in1(_gnd_net_),
            .in2(N__36109),
            .in3(N__44557),
            .lcout(data_out_frame2_17_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50522),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i0_LC_13_25_0.C_ON=1'b1;
    defparam rand_data_2350__i0_LC_13_25_0.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i0_LC_13_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i0_LC_13_25_0 (
            .in0(_gnd_net_),
            .in1(N__39522),
            .in2(_gnd_net_),
            .in3(N__36094),
            .lcout(rand_data_0),
            .ltout(),
            .carryin(bfn_13_25_0_),
            .carryout(n15528),
            .clk(N__50532),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i1_LC_13_25_1.C_ON=1'b1;
    defparam rand_data_2350__i1_LC_13_25_1.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i1_LC_13_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i1_LC_13_25_1 (
            .in0(_gnd_net_),
            .in1(N__36224),
            .in2(_gnd_net_),
            .in3(N__36091),
            .lcout(rand_data_1),
            .ltout(),
            .carryin(n15528),
            .carryout(n15529),
            .clk(N__50532),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i2_LC_13_25_2.C_ON=1'b1;
    defparam rand_data_2350__i2_LC_13_25_2.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i2_LC_13_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i2_LC_13_25_2 (
            .in0(_gnd_net_),
            .in1(N__36418),
            .in2(_gnd_net_),
            .in3(N__36088),
            .lcout(rand_data_2),
            .ltout(),
            .carryin(n15529),
            .carryout(n15530),
            .clk(N__50532),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i3_LC_13_25_3.C_ON=1'b1;
    defparam rand_data_2350__i3_LC_13_25_3.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i3_LC_13_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i3_LC_13_25_3 (
            .in0(_gnd_net_),
            .in1(N__49780),
            .in2(_gnd_net_),
            .in3(N__36085),
            .lcout(rand_data_3),
            .ltout(),
            .carryin(n15530),
            .carryout(n15531),
            .clk(N__50532),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i4_LC_13_25_4.C_ON=1'b1;
    defparam rand_data_2350__i4_LC_13_25_4.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i4_LC_13_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i4_LC_13_25_4 (
            .in0(_gnd_net_),
            .in1(N__37343),
            .in2(_gnd_net_),
            .in3(N__36082),
            .lcout(rand_data_4),
            .ltout(),
            .carryin(n15531),
            .carryout(n15532),
            .clk(N__50532),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i5_LC_13_25_5.C_ON=1'b1;
    defparam rand_data_2350__i5_LC_13_25_5.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i5_LC_13_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i5_LC_13_25_5 (
            .in0(_gnd_net_),
            .in1(N__41444),
            .in2(_gnd_net_),
            .in3(N__36079),
            .lcout(rand_data_5),
            .ltout(),
            .carryin(n15532),
            .carryout(n15533),
            .clk(N__50532),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i6_LC_13_25_6.C_ON=1'b1;
    defparam rand_data_2350__i6_LC_13_25_6.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i6_LC_13_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i6_LC_13_25_6 (
            .in0(_gnd_net_),
            .in1(N__49878),
            .in2(_gnd_net_),
            .in3(N__36160),
            .lcout(rand_data_6),
            .ltout(),
            .carryin(n15533),
            .carryout(n15534),
            .clk(N__50532),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i7_LC_13_25_7.C_ON=1'b1;
    defparam rand_data_2350__i7_LC_13_25_7.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i7_LC_13_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i7_LC_13_25_7 (
            .in0(_gnd_net_),
            .in1(N__51304),
            .in2(_gnd_net_),
            .in3(N__36157),
            .lcout(rand_data_7),
            .ltout(),
            .carryin(n15534),
            .carryout(n15535),
            .clk(N__50532),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i8_LC_13_26_0.C_ON=1'b1;
    defparam rand_data_2350__i8_LC_13_26_0.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i8_LC_13_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i8_LC_13_26_0 (
            .in0(_gnd_net_),
            .in1(N__48732),
            .in2(_gnd_net_),
            .in3(N__36154),
            .lcout(rand_data_8),
            .ltout(),
            .carryin(bfn_13_26_0_),
            .carryout(n15536),
            .clk(N__50543),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i9_LC_13_26_1.C_ON=1'b1;
    defparam rand_data_2350__i9_LC_13_26_1.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i9_LC_13_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i9_LC_13_26_1 (
            .in0(_gnd_net_),
            .in1(N__37896),
            .in2(_gnd_net_),
            .in3(N__36151),
            .lcout(rand_data_9),
            .ltout(),
            .carryin(n15536),
            .carryout(n15537),
            .clk(N__50543),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i10_LC_13_26_2.C_ON=1'b1;
    defparam rand_data_2350__i10_LC_13_26_2.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i10_LC_13_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i10_LC_13_26_2 (
            .in0(_gnd_net_),
            .in1(N__36596),
            .in2(_gnd_net_),
            .in3(N__36148),
            .lcout(rand_data_10),
            .ltout(),
            .carryin(n15537),
            .carryout(n15538),
            .clk(N__50543),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i11_LC_13_26_3.C_ON=1'b1;
    defparam rand_data_2350__i11_LC_13_26_3.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i11_LC_13_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i11_LC_13_26_3 (
            .in0(_gnd_net_),
            .in1(N__48815),
            .in2(_gnd_net_),
            .in3(N__36145),
            .lcout(rand_data_11),
            .ltout(),
            .carryin(n15538),
            .carryout(n15539),
            .clk(N__50543),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i12_LC_13_26_4.C_ON=1'b1;
    defparam rand_data_2350__i12_LC_13_26_4.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i12_LC_13_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i12_LC_13_26_4 (
            .in0(_gnd_net_),
            .in1(N__44139),
            .in2(_gnd_net_),
            .in3(N__36142),
            .lcout(rand_data_12),
            .ltout(),
            .carryin(n15539),
            .carryout(n15540),
            .clk(N__50543),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i13_LC_13_26_5.C_ON=1'b1;
    defparam rand_data_2350__i13_LC_13_26_5.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i13_LC_13_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i13_LC_13_26_5 (
            .in0(_gnd_net_),
            .in1(N__44547),
            .in2(_gnd_net_),
            .in3(N__36139),
            .lcout(rand_data_13),
            .ltout(),
            .carryin(n15540),
            .carryout(n15541),
            .clk(N__50543),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i14_LC_13_26_6.C_ON=1'b1;
    defparam rand_data_2350__i14_LC_13_26_6.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i14_LC_13_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i14_LC_13_26_6 (
            .in0(_gnd_net_),
            .in1(N__49073),
            .in2(_gnd_net_),
            .in3(N__36136),
            .lcout(rand_data_14),
            .ltout(),
            .carryin(n15541),
            .carryout(n15542),
            .clk(N__50543),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i15_LC_13_26_7.C_ON=1'b1;
    defparam rand_data_2350__i15_LC_13_26_7.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i15_LC_13_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i15_LC_13_26_7 (
            .in0(_gnd_net_),
            .in1(N__44918),
            .in2(_gnd_net_),
            .in3(N__36133),
            .lcout(rand_data_15),
            .ltout(),
            .carryin(n15542),
            .carryout(n15543),
            .clk(N__50543),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i16_LC_13_27_0.C_ON=1'b1;
    defparam rand_data_2350__i16_LC_13_27_0.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i16_LC_13_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i16_LC_13_27_0 (
            .in0(_gnd_net_),
            .in1(N__41733),
            .in2(_gnd_net_),
            .in3(N__36187),
            .lcout(rand_data_16),
            .ltout(),
            .carryin(bfn_13_27_0_),
            .carryout(n15544),
            .clk(N__50551),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i17_LC_13_27_1.C_ON=1'b1;
    defparam rand_data_2350__i17_LC_13_27_1.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i17_LC_13_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i17_LC_13_27_1 (
            .in0(_gnd_net_),
            .in1(N__39358),
            .in2(_gnd_net_),
            .in3(N__36184),
            .lcout(rand_data_17),
            .ltout(),
            .carryin(n15544),
            .carryout(n15545),
            .clk(N__50551),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i18_LC_13_27_2.C_ON=1'b1;
    defparam rand_data_2350__i18_LC_13_27_2.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i18_LC_13_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i18_LC_13_27_2 (
            .in0(_gnd_net_),
            .in1(N__44462),
            .in2(_gnd_net_),
            .in3(N__36181),
            .lcout(rand_data_18),
            .ltout(),
            .carryin(n15545),
            .carryout(n15546),
            .clk(N__50551),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i19_LC_13_27_3.C_ON=1'b1;
    defparam rand_data_2350__i19_LC_13_27_3.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i19_LC_13_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i19_LC_13_27_3 (
            .in0(_gnd_net_),
            .in1(N__36708),
            .in2(_gnd_net_),
            .in3(N__36178),
            .lcout(rand_data_19),
            .ltout(),
            .carryin(n15546),
            .carryout(n15547),
            .clk(N__50551),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i20_LC_13_27_4.C_ON=1'b1;
    defparam rand_data_2350__i20_LC_13_27_4.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i20_LC_13_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i20_LC_13_27_4 (
            .in0(_gnd_net_),
            .in1(N__39073),
            .in2(_gnd_net_),
            .in3(N__36175),
            .lcout(rand_data_20),
            .ltout(),
            .carryin(n15547),
            .carryout(n15548),
            .clk(N__50551),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i21_LC_13_27_5.C_ON=1'b1;
    defparam rand_data_2350__i21_LC_13_27_5.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i21_LC_13_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i21_LC_13_27_5 (
            .in0(_gnd_net_),
            .in1(N__40618),
            .in2(_gnd_net_),
            .in3(N__36172),
            .lcout(rand_data_21),
            .ltout(),
            .carryin(n15548),
            .carryout(n15549),
            .clk(N__50551),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i22_LC_13_27_6.C_ON=1'b1;
    defparam rand_data_2350__i22_LC_13_27_6.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i22_LC_13_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i22_LC_13_27_6 (
            .in0(_gnd_net_),
            .in1(N__41185),
            .in2(_gnd_net_),
            .in3(N__36169),
            .lcout(rand_data_22),
            .ltout(),
            .carryin(n15549),
            .carryout(n15550),
            .clk(N__50551),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i23_LC_13_27_7.C_ON=1'b1;
    defparam rand_data_2350__i23_LC_13_27_7.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i23_LC_13_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i23_LC_13_27_7 (
            .in0(_gnd_net_),
            .in1(N__44068),
            .in2(_gnd_net_),
            .in3(N__36166),
            .lcout(rand_data_23),
            .ltout(),
            .carryin(n15550),
            .carryout(n15551),
            .clk(N__50551),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i24_LC_13_28_0.C_ON=1'b1;
    defparam rand_data_2350__i24_LC_13_28_0.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i24_LC_13_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i24_LC_13_28_0 (
            .in0(_gnd_net_),
            .in1(N__44761),
            .in2(_gnd_net_),
            .in3(N__36163),
            .lcout(rand_data_24),
            .ltout(),
            .carryin(bfn_13_28_0_),
            .carryout(n15552),
            .clk(N__50561),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i25_LC_13_28_1.C_ON=1'b1;
    defparam rand_data_2350__i25_LC_13_28_1.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i25_LC_13_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i25_LC_13_28_1 (
            .in0(_gnd_net_),
            .in1(N__44666),
            .in2(_gnd_net_),
            .in3(N__36292),
            .lcout(rand_data_25),
            .ltout(),
            .carryin(n15552),
            .carryout(n15553),
            .clk(N__50561),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i26_LC_13_28_2.C_ON=1'b1;
    defparam rand_data_2350__i26_LC_13_28_2.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i26_LC_13_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i26_LC_13_28_2 (
            .in0(_gnd_net_),
            .in1(N__39622),
            .in2(_gnd_net_),
            .in3(N__36289),
            .lcout(rand_data_26),
            .ltout(),
            .carryin(n15553),
            .carryout(n15554),
            .clk(N__50561),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i27_LC_13_28_3.C_ON=1'b1;
    defparam rand_data_2350__i27_LC_13_28_3.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i27_LC_13_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i27_LC_13_28_3 (
            .in0(_gnd_net_),
            .in1(N__37936),
            .in2(_gnd_net_),
            .in3(N__36286),
            .lcout(rand_data_27),
            .ltout(),
            .carryin(n15554),
            .carryout(n15555),
            .clk(N__50561),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i28_LC_13_28_4.C_ON=1'b1;
    defparam rand_data_2350__i28_LC_13_28_4.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i28_LC_13_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i28_LC_13_28_4 (
            .in0(_gnd_net_),
            .in1(N__39198),
            .in2(_gnd_net_),
            .in3(N__36283),
            .lcout(rand_data_28),
            .ltout(),
            .carryin(n15555),
            .carryout(n15556),
            .clk(N__50561),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i29_LC_13_28_5.C_ON=1'b1;
    defparam rand_data_2350__i29_LC_13_28_5.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i29_LC_13_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i29_LC_13_28_5 (
            .in0(_gnd_net_),
            .in1(N__45279),
            .in2(_gnd_net_),
            .in3(N__36280),
            .lcout(rand_data_29),
            .ltout(),
            .carryin(n15556),
            .carryout(n15557),
            .clk(N__50561),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i30_LC_13_28_6.C_ON=1'b1;
    defparam rand_data_2350__i30_LC_13_28_6.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i30_LC_13_28_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i30_LC_13_28_6 (
            .in0(_gnd_net_),
            .in1(N__48912),
            .in2(_gnd_net_),
            .in3(N__36277),
            .lcout(rand_data_30),
            .ltout(),
            .carryin(n15557),
            .carryout(n15558),
            .clk(N__50561),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2350__i31_LC_13_28_7.C_ON=1'b0;
    defparam rand_data_2350__i31_LC_13_28_7.SEQ_MODE=4'b1000;
    defparam rand_data_2350__i31_LC_13_28_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2350__i31_LC_13_28_7 (
            .in0(_gnd_net_),
            .in1(N__43990),
            .in2(_gnd_net_),
            .in3(N__36274),
            .lcout(rand_data_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50561),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i0_LC_13_29_0.C_ON=1'b1;
    defparam rand_setpoint_2351__i0_LC_13_29_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i0_LC_13_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i0_LC_13_29_0 (
            .in0(_gnd_net_),
            .in1(N__39532),
            .in2(N__36267),
            .in3(_gnd_net_),
            .lcout(rand_setpoint_0),
            .ltout(),
            .carryin(bfn_13_29_0_),
            .carryout(n15559),
            .clk(N__50571),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i1_LC_13_29_1.C_ON=1'b1;
    defparam rand_setpoint_2351__i1_LC_13_29_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i1_LC_13_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i1_LC_13_29_1 (
            .in0(_gnd_net_),
            .in1(N__36232),
            .in2(N__40569),
            .in3(N__36190),
            .lcout(rand_setpoint_1),
            .ltout(),
            .carryin(n15559),
            .carryout(n15560),
            .clk(N__50571),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i2_LC_13_29_2.C_ON=1'b1;
    defparam rand_setpoint_2351__i2_LC_13_29_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i2_LC_13_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i2_LC_13_29_2 (
            .in0(_gnd_net_),
            .in1(N__36424),
            .in2(N__38163),
            .in3(N__36394),
            .lcout(rand_setpoint_2),
            .ltout(),
            .carryin(n15560),
            .carryout(n15561),
            .clk(N__50571),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i3_LC_13_29_3.C_ON=1'b1;
    defparam rand_setpoint_2351__i3_LC_13_29_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i3_LC_13_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i3_LC_13_29_3 (
            .in0(_gnd_net_),
            .in1(N__49784),
            .in2(N__36391),
            .in3(N__36376),
            .lcout(rand_setpoint_3),
            .ltout(),
            .carryin(n15561),
            .carryout(n15562),
            .clk(N__50571),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i4_LC_13_29_4.C_ON=1'b1;
    defparam rand_setpoint_2351__i4_LC_13_29_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i4_LC_13_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i4_LC_13_29_4 (
            .in0(_gnd_net_),
            .in1(N__37354),
            .in2(N__36373),
            .in3(N__36358),
            .lcout(rand_setpoint_4),
            .ltout(),
            .carryin(n15562),
            .carryout(n15563),
            .clk(N__50571),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i5_LC_13_29_5.C_ON=1'b1;
    defparam rand_setpoint_2351__i5_LC_13_29_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i5_LC_13_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i5_LC_13_29_5 (
            .in0(_gnd_net_),
            .in1(N__41465),
            .in2(N__40104),
            .in3(N__36355),
            .lcout(rand_setpoint_5),
            .ltout(),
            .carryin(n15563),
            .carryout(n15564),
            .clk(N__50571),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i6_LC_13_29_6.C_ON=1'b1;
    defparam rand_setpoint_2351__i6_LC_13_29_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i6_LC_13_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i6_LC_13_29_6 (
            .in0(_gnd_net_),
            .in1(N__49897),
            .in2(N__40044),
            .in3(N__36352),
            .lcout(rand_setpoint_6),
            .ltout(),
            .carryin(n15564),
            .carryout(n15565),
            .clk(N__50571),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i7_LC_13_29_7.C_ON=1'b1;
    defparam rand_setpoint_2351__i7_LC_13_29_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i7_LC_13_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i7_LC_13_29_7 (
            .in0(_gnd_net_),
            .in1(N__38205),
            .in2(N__51327),
            .in3(N__36349),
            .lcout(rand_setpoint_7),
            .ltout(),
            .carryin(n15565),
            .carryout(n15566),
            .clk(N__50571),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i8_LC_13_30_0.C_ON=1'b1;
    defparam rand_setpoint_2351__i8_LC_13_30_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i8_LC_13_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i8_LC_13_30_0 (
            .in0(_gnd_net_),
            .in1(N__48744),
            .in2(N__36339),
            .in3(N__36322),
            .lcout(rand_setpoint_8),
            .ltout(),
            .carryin(bfn_13_30_0_),
            .carryout(n15567),
            .clk(N__50579),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i9_LC_13_30_1.C_ON=1'b1;
    defparam rand_setpoint_2351__i9_LC_13_30_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i9_LC_13_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i9_LC_13_30_1 (
            .in0(_gnd_net_),
            .in1(N__37901),
            .in2(N__36312),
            .in3(N__36295),
            .lcout(rand_setpoint_9),
            .ltout(),
            .carryin(n15567),
            .carryout(n15568),
            .clk(N__50579),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i10_LC_13_30_2.C_ON=1'b1;
    defparam rand_setpoint_2351__i10_LC_13_30_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i10_LC_13_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i10_LC_13_30_2 (
            .in0(_gnd_net_),
            .in1(N__36609),
            .in2(N__46017),
            .in3(N__36565),
            .lcout(rand_setpoint_10),
            .ltout(),
            .carryin(n15568),
            .carryout(n15569),
            .clk(N__50579),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i11_LC_13_30_3.C_ON=1'b1;
    defparam rand_setpoint_2351__i11_LC_13_30_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i11_LC_13_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i11_LC_13_30_3 (
            .in0(_gnd_net_),
            .in1(N__48828),
            .in2(N__36555),
            .in3(N__36538),
            .lcout(rand_setpoint_11),
            .ltout(),
            .carryin(n15569),
            .carryout(n15570),
            .clk(N__50579),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i12_LC_13_30_4.C_ON=1'b1;
    defparam rand_setpoint_2351__i12_LC_13_30_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i12_LC_13_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i12_LC_13_30_4 (
            .in0(_gnd_net_),
            .in1(N__36528),
            .in2(N__44164),
            .in3(N__36517),
            .lcout(rand_setpoint_12),
            .ltout(),
            .carryin(n15570),
            .carryout(n15571),
            .clk(N__50579),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i13_LC_13_30_5.C_ON=1'b1;
    defparam rand_setpoint_2351__i13_LC_13_30_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i13_LC_13_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i13_LC_13_30_5 (
            .in0(_gnd_net_),
            .in1(N__36507),
            .in2(N__44566),
            .in3(N__36496),
            .lcout(rand_setpoint_13),
            .ltout(),
            .carryin(n15571),
            .carryout(n15572),
            .clk(N__50579),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i14_LC_13_30_6.C_ON=1'b1;
    defparam rand_setpoint_2351__i14_LC_13_30_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i14_LC_13_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i14_LC_13_30_6 (
            .in0(_gnd_net_),
            .in1(N__49095),
            .in2(N__36492),
            .in3(N__36475),
            .lcout(rand_setpoint_14),
            .ltout(),
            .carryin(n15572),
            .carryout(n15573),
            .clk(N__50579),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i15_LC_13_30_7.C_ON=1'b1;
    defparam rand_setpoint_2351__i15_LC_13_30_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i15_LC_13_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i15_LC_13_30_7 (
            .in0(_gnd_net_),
            .in1(N__36465),
            .in2(N__44943),
            .in3(N__36454),
            .lcout(rand_setpoint_15),
            .ltout(),
            .carryin(n15573),
            .carryout(n15574),
            .clk(N__50579),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i16_LC_13_31_0.C_ON=1'b1;
    defparam rand_setpoint_2351__i16_LC_13_31_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i16_LC_13_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i16_LC_13_31_0 (
            .in0(_gnd_net_),
            .in1(N__41752),
            .in2(N__42882),
            .in3(N__36451),
            .lcout(rand_setpoint_16),
            .ltout(),
            .carryin(bfn_13_31_0_),
            .carryout(n15575),
            .clk(N__50585),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i17_LC_13_31_1.C_ON=1'b1;
    defparam rand_setpoint_2351__i17_LC_13_31_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i17_LC_13_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i17_LC_13_31_1 (
            .in0(_gnd_net_),
            .in1(N__39374),
            .in2(N__38272),
            .in3(N__36448),
            .lcout(rand_setpoint_17),
            .ltout(),
            .carryin(n15575),
            .carryout(n15576),
            .clk(N__50585),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i18_LC_13_31_2.C_ON=1'b1;
    defparam rand_setpoint_2351__i18_LC_13_31_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i18_LC_13_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i18_LC_13_31_2 (
            .in0(_gnd_net_),
            .in1(N__44470),
            .in2(N__38299),
            .in3(N__36445),
            .lcout(rand_setpoint_18),
            .ltout(),
            .carryin(n15576),
            .carryout(n15577),
            .clk(N__50585),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i19_LC_13_31_3.C_ON=1'b1;
    defparam rand_setpoint_2351__i19_LC_13_31_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i19_LC_13_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i19_LC_13_31_3 (
            .in0(_gnd_net_),
            .in1(N__36718),
            .in2(N__38332),
            .in3(N__36679),
            .lcout(rand_setpoint_19),
            .ltout(),
            .carryin(n15577),
            .carryout(n15578),
            .clk(N__50585),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i20_LC_13_31_4.C_ON=1'b1;
    defparam rand_setpoint_2351__i20_LC_13_31_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i20_LC_13_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i20_LC_13_31_4 (
            .in0(_gnd_net_),
            .in1(N__39082),
            .in2(N__38362),
            .in3(N__36676),
            .lcout(rand_setpoint_20),
            .ltout(),
            .carryin(n15578),
            .carryout(n15579),
            .clk(N__50585),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i21_LC_13_31_5.C_ON=1'b1;
    defparam rand_setpoint_2351__i21_LC_13_31_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i21_LC_13_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i21_LC_13_31_5 (
            .in0(_gnd_net_),
            .in1(N__40634),
            .in2(N__46518),
            .in3(N__36673),
            .lcout(rand_setpoint_21),
            .ltout(),
            .carryin(n15579),
            .carryout(n15580),
            .clk(N__50585),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i22_LC_13_31_6.C_ON=1'b1;
    defparam rand_setpoint_2351__i22_LC_13_31_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i22_LC_13_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i22_LC_13_31_6 (
            .in0(_gnd_net_),
            .in1(N__41203),
            .in2(N__36670),
            .in3(N__36655),
            .lcout(rand_setpoint_22),
            .ltout(),
            .carryin(n15580),
            .carryout(n15581),
            .clk(N__50585),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i23_LC_13_31_7.C_ON=1'b1;
    defparam rand_setpoint_2351__i23_LC_13_31_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i23_LC_13_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i23_LC_13_31_7 (
            .in0(_gnd_net_),
            .in1(N__44081),
            .in2(N__40290),
            .in3(N__36652),
            .lcout(rand_setpoint_23),
            .ltout(),
            .carryin(n15581),
            .carryout(n15582),
            .clk(N__50585),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i24_LC_13_32_0.C_ON=1'b1;
    defparam rand_setpoint_2351__i24_LC_13_32_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i24_LC_13_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i24_LC_13_32_0 (
            .in0(_gnd_net_),
            .in1(N__44782),
            .in2(N__38224),
            .in3(N__36649),
            .lcout(rand_setpoint_24),
            .ltout(),
            .carryin(bfn_13_32_0_),
            .carryout(n15583),
            .clk(N__50589),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i25_LC_13_32_1.C_ON=1'b1;
    defparam rand_setpoint_2351__i25_LC_13_32_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i25_LC_13_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i25_LC_13_32_1 (
            .in0(_gnd_net_),
            .in1(N__44686),
            .in2(N__36646),
            .in3(N__36631),
            .lcout(rand_setpoint_25),
            .ltout(),
            .carryin(n15583),
            .carryout(n15584),
            .clk(N__50589),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i26_LC_13_32_2.C_ON=1'b1;
    defparam rand_setpoint_2351__i26_LC_13_32_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i26_LC_13_32_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i26_LC_13_32_2 (
            .in0(_gnd_net_),
            .in1(N__38253),
            .in2(N__39636),
            .in3(N__36628),
            .lcout(rand_setpoint_26),
            .ltout(),
            .carryin(n15584),
            .carryout(n15585),
            .clk(N__50589),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i27_LC_13_32_3.C_ON=1'b1;
    defparam rand_setpoint_2351__i27_LC_13_32_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i27_LC_13_32_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i27_LC_13_32_3 (
            .in0(_gnd_net_),
            .in1(N__37945),
            .in2(N__38641),
            .in3(N__36625),
            .lcout(rand_setpoint_27),
            .ltout(),
            .carryin(n15585),
            .carryout(n15586),
            .clk(N__50589),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i28_LC_13_32_4.C_ON=1'b1;
    defparam rand_setpoint_2351__i28_LC_13_32_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i28_LC_13_32_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i28_LC_13_32_4 (
            .in0(_gnd_net_),
            .in1(N__39202),
            .in2(N__38626),
            .in3(N__36877),
            .lcout(rand_setpoint_28),
            .ltout(),
            .carryin(n15586),
            .carryout(n15587),
            .clk(N__50589),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i29_LC_13_32_5.C_ON=1'b1;
    defparam rand_setpoint_2351__i29_LC_13_32_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i29_LC_13_32_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i29_LC_13_32_5 (
            .in0(_gnd_net_),
            .in1(N__45292),
            .in2(N__38241),
            .in3(N__36874),
            .lcout(rand_setpoint_29),
            .ltout(),
            .carryin(n15587),
            .carryout(n15588),
            .clk(N__50589),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i30_LC_13_32_6.C_ON=1'b1;
    defparam rand_setpoint_2351__i30_LC_13_32_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i30_LC_13_32_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2351__i30_LC_13_32_6 (
            .in0(_gnd_net_),
            .in1(N__48934),
            .in2(N__36871),
            .in3(N__36856),
            .lcout(rand_setpoint_30),
            .ltout(),
            .carryin(n15588),
            .carryout(n15589),
            .clk(N__50589),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2351__i31_LC_13_32_7.C_ON=1'b0;
    defparam rand_setpoint_2351__i31_LC_13_32_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2351__i31_LC_13_32_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 rand_setpoint_2351__i31_LC_13_32_7 (
            .in0(N__44002),
            .in1(N__36850),
            .in2(_gnd_net_),
            .in3(N__36853),
            .lcout(rand_setpoint_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50589),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_537_LC_14_17_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_537_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_537_LC_14_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_537_LC_14_17_0  (
            .in0(N__52513),
            .in1(N__40351),
            .in2(_gnd_net_),
            .in3(N__36838),
            .lcout(\c0.n17064 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_14_18_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_14_18_0 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_14_18_0  (
            .in0(N__47821),
            .in1(N__48955),
            .in2(N__38791),
            .in3(N__47659),
            .lcout(),
            .ltout(\c0.n22_adj_2357_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i3_LC_14_18_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i3_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i3_LC_14_18_1 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.tx2.r_Tx_Data_i3_LC_14_18_1  (
            .in0(N__51609),
            .in1(N__36769),
            .in2(N__36796),
            .in3(N__51738),
            .lcout(\c0.tx2.r_Tx_Data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50468),
            .ce(N__51447),
            .sr(_gnd_net_));
    defparam \c0.n18125_bdd_4_lut_LC_14_18_4 .C_ON=1'b0;
    defparam \c0.n18125_bdd_4_lut_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18125_bdd_4_lut_LC_14_18_4 .LUT_INIT=16'b1010101011011000;
    LogicCell40 \c0.n18125_bdd_4_lut_LC_14_18_4  (
            .in0(N__38386),
            .in1(N__36781),
            .in2(N__40744),
            .in3(N__51608),
            .lcout(\c0.n18128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_644_LC_14_19_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_644_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_644_LC_14_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_644_LC_14_19_1  (
            .in0(N__40799),
            .in1(N__49198),
            .in2(N__36763),
            .in3(N__41242),
            .lcout(\c0.n18_adj_2331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_573_LC_14_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_573_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_573_LC_14_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_573_LC_14_19_2  (
            .in0(N__49557),
            .in1(N__43465),
            .in2(_gnd_net_),
            .in3(N__37149),
            .lcout(\c0.n17100 ),
            .ltout(\c0.n17100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_LC_14_19_3 .C_ON=1'b0;
    defparam \c0.i5_2_lut_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_LC_14_19_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i5_2_lut_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36955),
            .in3(N__41934),
            .lcout(),
            .ltout(\c0.n16_adj_2332_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i153_LC_14_19_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i153_LC_14_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i153_LC_14_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i153_LC_14_19_4  (
            .in0(N__38419),
            .in1(N__37195),
            .in2(N__36952),
            .in3(N__36949),
            .lcout(\c0.data_out_frame2_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50481),
            .ce(N__51185),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_481_LC_14_20_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_481_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_481_LC_14_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_481_LC_14_20_0  (
            .in0(N__39670),
            .in1(N__43189),
            .in2(N__42010),
            .in3(N__39496),
            .lcout(),
            .ltout(\c0.n12_adj_2263_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i163_LC_14_20_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i163_LC_14_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i163_LC_14_20_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i163_LC_14_20_1  (
            .in0(N__36928),
            .in1(N__41068),
            .in2(N__36922),
            .in3(N__38833),
            .lcout(\c0.data_out_frame2_20_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50493),
            .ce(N__51182),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_590_LC_14_20_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_590_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_590_LC_14_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_590_LC_14_20_3  (
            .in0(N__39435),
            .in1(N__37588),
            .in2(N__37054),
            .in3(N__37624),
            .lcout(),
            .ltout(\c0.n16_adj_2312_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i157_LC_14_20_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i157_LC_14_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i157_LC_14_20_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i157_LC_14_20_4  (
            .in0(N__36907),
            .in1(N__36888),
            .in2(N__36895),
            .in3(N__38401),
            .lcout(\c0.data_out_frame2_19_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50493),
            .ce(N__51182),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_584_LC_14_20_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_584_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_584_LC_14_20_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_584_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__43309),
            .in2(_gnd_net_),
            .in3(N__39669),
            .lcout(\c0.n17097 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_14_20_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_14_20_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_14_20_6  (
            .in0(N__39668),
            .in1(N__48092),
            .in2(_gnd_net_),
            .in3(N__37147),
            .lcout(\c0.n5_adj_2334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_480_LC_14_21_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_480_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_480_LC_14_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_480_LC_14_21_1  (
            .in0(N__37117),
            .in1(N__38541),
            .in2(N__49476),
            .in3(N__38976),
            .lcout(\c0.n17052 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_4_lut_LC_14_21_2 .C_ON=1'b0;
    defparam \c0.i7_3_lut_4_lut_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_4_lut_LC_14_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_3_lut_4_lut_LC_14_21_2  (
            .in0(N__37737),
            .in1(N__40148),
            .in2(N__37077),
            .in3(N__49015),
            .lcout(\c0.n20_adj_2202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_593_LC_14_21_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_593_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_593_LC_14_21_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_593_LC_14_21_3  (
            .in0(N__37042),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38462),
            .lcout(\c0.n9839 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_LC_14_21_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_LC_14_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_LC_14_21_4  (
            .in0(N__41110),
            .in1(N__43524),
            .in2(_gnd_net_),
            .in3(N__38679),
            .lcout(\c0.n14_adj_2264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17957_bdd_4_lut_LC_14_21_5 .C_ON=1'b0;
    defparam \c0.n17957_bdd_4_lut_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.n17957_bdd_4_lut_LC_14_21_5 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \c0.n17957_bdd_4_lut_LC_14_21_5  (
            .in0(N__48512),
            .in1(N__37156),
            .in2(N__37305),
            .in3(N__40725),
            .lcout(\c0.n17960 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_490_LC_14_21_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_490_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_490_LC_14_21_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_490_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__37041),
            .in2(_gnd_net_),
            .in3(N__44434),
            .lcout(\c0.n17031 ),
            .ltout(\c0.n17031_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_493_LC_14_21_7 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_493_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_493_LC_14_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_493_LC_14_21_7  (
            .in0(N__37003),
            .in1(N__37692),
            .in2(N__36991),
            .in3(N__37264),
            .lcout(\c0.n26_adj_2273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_447_LC_14_22_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_447_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_447_LC_14_22_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_447_LC_14_22_0  (
            .in0(N__38773),
            .in1(N__45628),
            .in2(_gnd_net_),
            .in3(N__36988),
            .lcout(\c0.n17085 ),
            .ltout(\c0.n17085_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_445_LC_14_22_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_445_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_445_LC_14_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_445_LC_14_22_1  (
            .in0(N__37309),
            .in1(N__44307),
            .in2(N__37267),
            .in3(N__37263),
            .lcout(\c0.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15523_LC_14_22_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15523_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15523_LC_14_22_2 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15523_LC_14_22_2  (
            .in0(N__37243),
            .in1(N__48142),
            .in2(N__48583),
            .in3(N__37222),
            .lcout(\c0.n17969 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_607_LC_14_22_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_607_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_607_LC_14_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_607_LC_14_22_3  (
            .in0(N__37849),
            .in1(N__37174),
            .in2(_gnd_net_),
            .in3(N__37213),
            .lcout(\c0.n17088 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_606_LC_14_22_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_606_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_606_LC_14_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_606_LC_14_22_4  (
            .in0(N__45363),
            .in1(N__37191),
            .in2(N__49290),
            .in3(N__41160),
            .lcout(\c0.n9579 ),
            .ltout(\c0.n9579_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_579_LC_14_22_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_579_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_579_LC_14_22_5 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \c0.i2_2_lut_adj_579_LC_14_22_5  (
            .in0(_gnd_net_),
            .in1(N__38774),
            .in2(N__37168),
            .in3(_gnd_net_),
            .lcout(\c0.n10_adj_2307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15621_LC_14_22_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15621_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15621_LC_14_22_6 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15621_LC_14_22_6  (
            .in0(N__38892),
            .in1(N__48141),
            .in2(N__48582),
            .in3(N__41159),
            .lcout(\c0.n18071 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15514_LC_14_22_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15514_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15514_LC_14_22_7 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15514_LC_14_22_7  (
            .in0(N__48140),
            .in1(N__41831),
            .in2(N__48581),
            .in3(N__41263),
            .lcout(\c0.n17957 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i90_LC_14_23_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i90_LC_14_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i90_LC_14_23_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_out_frame2_0___i90_LC_14_23_0  (
            .in0(N__41535),
            .in1(N__50936),
            .in2(_gnd_net_),
            .in3(N__37910),
            .lcout(data_out_frame2_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50523),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i68_LC_14_23_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i68_LC_14_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i68_LC_14_23_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i68_LC_14_23_1  (
            .in0(N__50932),
            .in1(N__49802),
            .in2(_gnd_net_),
            .in3(N__40724),
            .lcout(data_out_frame2_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50523),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i81_LC_14_23_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i81_LC_14_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i81_LC_14_23_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i81_LC_14_23_2  (
            .in0(N__41753),
            .in1(N__50935),
            .in2(_gnd_net_),
            .in3(N__43572),
            .lcout(data_out_frame2_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50523),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_525_LC_14_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_525_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_525_LC_14_23_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_525_LC_14_23_3  (
            .in0(_gnd_net_),
            .in1(N__41534),
            .in2(_gnd_net_),
            .in3(N__40860),
            .lcout(\c0.n16908 ),
            .ltout(\c0.n16908_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_475_LC_14_23_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_475_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_475_LC_14_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_475_LC_14_23_4  (
            .in0(N__49698),
            .in1(N__38890),
            .in2(N__37597),
            .in3(N__41264),
            .lcout(\c0.n17022 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_684_LC_14_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_684_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_684_LC_14_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_684_LC_14_23_5  (
            .in0(N__39275),
            .in1(N__39128),
            .in2(_gnd_net_),
            .in3(N__49423),
            .lcout(\c0.n6_adj_2286 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i104_LC_14_23_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i104_LC_14_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i104_LC_14_23_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i104_LC_14_23_6  (
            .in0(N__51328),
            .in1(N__50934),
            .in2(_gnd_net_),
            .in3(N__43756),
            .lcout(data_out_frame2_12_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50523),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i92_LC_14_23_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i92_LC_14_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i92_LC_14_23_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_out_frame2_0___i92_LC_14_23_7  (
            .in0(N__50933),
            .in1(_gnd_net_),
            .in2(N__41269),
            .in3(N__48829),
            .lcout(data_out_frame2_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50523),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i117_LC_14_24_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i117_LC_14_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i117_LC_14_24_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i117_LC_14_24_0  (
            .in0(N__39090),
            .in1(N__37579),
            .in2(_gnd_net_),
            .in3(N__51104),
            .lcout(data_out_frame2_14_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50533),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15414_3_lut_LC_14_24_1 .C_ON=1'b0;
    defparam \c0.i15414_3_lut_LC_14_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15414_3_lut_LC_14_24_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \c0.i15414_3_lut_LC_14_24_1  (
            .in0(N__37555),
            .in1(N__37453),
            .in2(_gnd_net_),
            .in3(N__37383),
            .lcout(n10197),
            .ltout(n10197_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i69_LC_14_24_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i69_LC_14_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i69_LC_14_24_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_out_frame2_0___i69_LC_14_24_2  (
            .in0(N__37349),
            .in1(_gnd_net_),
            .in2(N__37312),
            .in3(N__49324),
            .lcout(data_out_frame2_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50533),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i82_LC_14_24_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i82_LC_14_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i82_LC_14_24_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i82_LC_14_24_3  (
            .in0(N__51102),
            .in1(N__39368),
            .in2(_gnd_net_),
            .in3(N__47409),
            .lcout(data_out_frame2_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50533),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i119_LC_14_24_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i119_LC_14_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i119_LC_14_24_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i119_LC_14_24_4  (
            .in0(N__41204),
            .in1(N__43678),
            .in2(_gnd_net_),
            .in3(N__51105),
            .lcout(data_out_frame2_14_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50533),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_575_LC_14_24_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_575_LC_14_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_575_LC_14_24_5 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \c0.i2_3_lut_adj_575_LC_14_24_5  (
            .in0(N__49323),
            .in1(N__37766),
            .in2(N__39495),
            .in3(_gnd_net_),
            .lcout(\c0.n9749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i102_LC_14_24_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i102_LC_14_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i102_LC_14_24_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i102_LC_14_24_6  (
            .in0(N__37732),
            .in1(N__41454),
            .in2(_gnd_net_),
            .in3(N__51103),
            .lcout(data_out_frame2_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50533),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_629_LC_14_24_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_629_LC_14_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_629_LC_14_24_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_629_LC_14_24_7  (
            .in0(N__40774),
            .in1(N__41859),
            .in2(N__43267),
            .in3(N__41689),
            .lcout(\c0.n17049 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i75_LC_14_25_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i75_LC_14_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i75_LC_14_25_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i75_LC_14_25_1  (
            .in0(N__39635),
            .in1(N__43884),
            .in2(_gnd_net_),
            .in3(N__50927),
            .lcout(data_out_frame2_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50544),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15224_3_lut_LC_14_25_2 .C_ON=1'b0;
    defparam \c0.i15224_3_lut_LC_14_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15224_3_lut_LC_14_25_2 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \c0.i15224_3_lut_LC_14_25_2  (
            .in0(N__48165),
            .in1(N__49536),
            .in2(_gnd_net_),
            .in3(N__48585),
            .lcout(\c0.n17561 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_631_LC_14_25_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_631_LC_14_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_631_LC_14_25_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_631_LC_14_25_3  (
            .in0(_gnd_net_),
            .in1(N__49535),
            .in2(_gnd_net_),
            .in3(N__48705),
            .lcout(\c0.n9589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i43_LC_14_25_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i43_LC_14_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i43_LC_14_25_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i43_LC_14_25_4  (
            .in0(N__50925),
            .in1(N__39634),
            .in2(_gnd_net_),
            .in3(N__37651),
            .lcout(data_out_frame2_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50544),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_576_LC_14_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_576_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_576_LC_14_25_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_576_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(N__37623),
            .in2(_gnd_net_),
            .in3(N__39038),
            .lcout(),
            .ltout(\c0.n6_adj_2306_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_577_LC_14_25_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_577_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_577_LC_14_25_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_577_LC_14_25_6  (
            .in0(N__38893),
            .in1(N__45248),
            .in2(N__37960),
            .in3(N__49503),
            .lcout(\c0.n16987 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i42_LC_14_25_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i42_LC_14_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i42_LC_14_25_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i42_LC_14_25_7  (
            .in0(N__44687),
            .in1(N__39013),
            .in2(_gnd_net_),
            .in3(N__50926),
            .lcout(data_out_frame2_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50544),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i108_LC_14_26_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i108_LC_14_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i108_LC_14_26_0 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.data_out_frame2_0___i108_LC_14_26_0  (
            .in0(N__37946),
            .in1(N__39274),
            .in2(N__51246),
            .in3(_gnd_net_),
            .lcout(data_out_frame2_13_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50552),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_444_LC_14_26_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_444_LC_14_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_444_LC_14_26_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_444_LC_14_26_1  (
            .in0(_gnd_net_),
            .in1(N__43682),
            .in2(_gnd_net_),
            .in3(N__48706),
            .lcout(\c0.n10_adj_2191 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i138_LC_14_26_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i138_LC_14_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i138_LC_14_26_2 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.data_out_frame2_0___i138_LC_14_26_2  (
            .in0(N__37897),
            .in1(N__37863),
            .in2(N__51247),
            .in3(_gnd_net_),
            .lcout(data_out_frame2_17_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50552),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i85_LC_14_26_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i85_LC_14_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i85_LC_14_26_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.data_out_frame2_0___i85_LC_14_26_5  (
            .in0(_gnd_net_),
            .in1(N__51161),
            .in2(N__39083),
            .in3(N__37837),
            .lcout(data_out_frame2_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50552),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i168_LC_14_27_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i168_LC_14_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i168_LC_14_27_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i168_LC_14_27_0  (
            .in0(N__41608),
            .in1(N__43766),
            .in2(N__37807),
            .in3(N__37798),
            .lcout(\c0.data_out_frame2_20_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50562),
            .ce(N__51181),
            .sr(_gnd_net_));
    defparam \c0.i15256_3_lut_LC_14_27_5 .C_ON=1'b0;
    defparam \c0.i15256_3_lut_LC_14_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15256_3_lut_LC_14_27_5 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \c0.i15256_3_lut_LC_14_27_5  (
            .in0(N__42396),
            .in1(N__42754),
            .in2(_gnd_net_),
            .in3(N__40228),
            .lcout(\c0.n17528 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15245_3_lut_LC_14_27_6 .C_ON=1'b0;
    defparam \c0.i15245_3_lut_LC_14_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15245_3_lut_LC_14_27_6 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \c0.i15245_3_lut_LC_14_27_6  (
            .in0(N__45205),
            .in1(_gnd_net_),
            .in2(N__42763),
            .in3(N__52140),
            .lcout(\c0.n17507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__2__2162_LC_14_28_0 .C_ON=1'b0;
    defparam \c0.data_out_10__2__2162_LC_14_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__2__2162_LC_14_28_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__2__2162_LC_14_28_0  (
            .in0(N__38107),
            .in1(N__46803),
            .in2(N__38065),
            .in3(N__46911),
            .lcout(\c0.data_out_10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50572),
            .ce(N__46620),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_533_LC_14_28_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_533_LC_14_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_533_LC_14_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_533_LC_14_28_2  (
            .in0(N__39957),
            .in1(N__39721),
            .in2(N__38064),
            .in3(N__42464),
            .lcout(),
            .ltout(\c0.n12_adj_2289_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__1__2163_LC_14_28_3 .C_ON=1'b0;
    defparam \c0.data_out_10__1__2163_LC_14_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__1__2163_LC_14_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__1__2163_LC_14_28_3  (
            .in0(N__46697),
            .in1(N__47140),
            .in2(N__38041),
            .in3(N__39730),
            .lcout(\c0.data_out_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50572),
            .ce(N__46620),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__0__2164_LC_14_28_5 .C_ON=1'b0;
    defparam \c0.data_out_10__0__2164_LC_14_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__0__2164_LC_14_28_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__0__2164_LC_14_28_5  (
            .in0(N__38038),
            .in1(N__42288),
            .in2(N__42217),
            .in3(N__39729),
            .lcout(\c0.data_out_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50572),
            .ce(N__46620),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_524_LC_14_29_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_524_LC_14_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_524_LC_14_29_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_524_LC_14_29_0  (
            .in0(N__39832),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39898),
            .lcout(\c0.n9496 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_494_LC_14_29_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_494_LC_14_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_494_LC_14_29_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_494_LC_14_29_1  (
            .in0(_gnd_net_),
            .in1(N__40479),
            .in2(_gnd_net_),
            .in3(N__40025),
            .lcout(\c0.n6_adj_2274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_LC_14_29_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_LC_14_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_LC_14_29_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_LC_14_29_2  (
            .in0(N__40024),
            .in1(N__40077),
            .in2(_gnd_net_),
            .in3(N__52136),
            .lcout(\c0.n9716 ),
            .ltout(\c0.n9716_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_693_LC_14_29_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_693_LC_14_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_693_LC_14_29_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_693_LC_14_29_3  (
            .in0(N__46739),
            .in1(N__52544),
            .in2(N__37996),
            .in3(N__37989),
            .lcout(),
            .ltout(\c0.n10_adj_2162_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_LC_14_29_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_LC_14_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_LC_14_29_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_LC_14_29_4  (
            .in0(N__46646),
            .in1(N__45201),
            .in2(N__37975),
            .in3(N__45106),
            .lcout(data_out_9__2__N_367),
            .ltout(data_out_9__2__N_367_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_686_LC_14_29_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_686_LC_14_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_686_LC_14_29_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_686_LC_14_29_5  (
            .in0(N__39899),
            .in1(_gnd_net_),
            .in2(N__37963),
            .in3(N__39833),
            .lcout(\c0.n17094 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_648_LC_14_29_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_648_LC_14_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_648_LC_14_29_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_648_LC_14_29_6  (
            .in0(N__39813),
            .in1(N__40057),
            .in2(N__40413),
            .in3(N__46863),
            .lcout(\c0.n16998 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__7__2173_LC_14_29_7 .C_ON=1'b0;
    defparam \c0.data_out_8__7__2173_LC_14_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__7__2173_LC_14_29_7 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_8__7__2173_LC_14_29_7  (
            .in0(N__45107),
            .in1(N__42745),
            .in2(N__38209),
            .in3(N__42838),
            .lcout(data_out_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50580),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_14_30_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_14_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_14_30_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_14_30_0  (
            .in0(N__52091),
            .in1(N__46798),
            .in2(_gnd_net_),
            .in3(N__40023),
            .lcout(),
            .ltout(\c0.n8_adj_2169_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_14_30_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_14_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_14_30_1 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_14_30_1  (
            .in0(N__52301),
            .in1(N__46647),
            .in2(N__38194),
            .in3(N__52092),
            .lcout(n10_adj_2427),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_484_LC_14_30_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_484_LC_14_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_484_LC_14_30_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_484_LC_14_30_2  (
            .in0(N__46200),
            .in1(N__38179),
            .in2(N__38173),
            .in3(N__40269),
            .lcout(\c0.n10_adj_2268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__2__2178_LC_14_30_3 .C_ON=1'b0;
    defparam \c0.data_out_8__2__2178_LC_14_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__2__2178_LC_14_30_3 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_8__2__2178_LC_14_30_3  (
            .in0(N__42847),
            .in1(N__42760),
            .in2(N__38164),
            .in3(N__39875),
            .lcout(\c0.data_out_8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50586),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15347_2_lut_LC_14_30_4 .C_ON=1'b0;
    defparam \c0.i15347_2_lut_LC_14_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15347_2_lut_LC_14_30_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15347_2_lut_LC_14_30_4  (
            .in0(N__52090),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38115),
            .lcout(\c0.n17594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_14_30_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_14_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_14_30_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_14_30_5  (
            .in0(N__45099),
            .in1(N__46969),
            .in2(_gnd_net_),
            .in3(N__52089),
            .lcout(\c0.n8_adj_2176 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__2__2234_LC_14_30_6 .C_ON=1'b0;
    defparam \c0.data_out_1__2__2234_LC_14_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__2__2234_LC_14_30_6 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \c0.data_out_1__2__2234_LC_14_30_6  (
            .in0(N__46488),
            .in1(N__38116),
            .in2(N__46138),
            .in3(N__42727),
            .lcout(\c0.data_out_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50586),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__7__2221_LC_14_30_7 .C_ON=1'b0;
    defparam \c0.data_out_2__7__2221_LC_14_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__7__2221_LC_14_30_7 .LUT_INIT=16'b1000110011011100;
    LogicCell40 \c0.data_out_2__7__2221_LC_14_30_7  (
            .in0(N__45455),
            .in1(N__38379),
            .in2(N__46000),
            .in3(N__46489),
            .lcout(data_out_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50586),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__4__2192_LC_14_31_1 .C_ON=1'b0;
    defparam \c0.data_out_6__4__2192_LC_14_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__4__2192_LC_14_31_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_6__4__2192_LC_14_31_1  (
            .in0(N__38361),
            .in1(N__45803),
            .in2(N__38347),
            .in3(N__46420),
            .lcout(\c0.data_out_6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50590),
            .ce(N__46130),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__3__2193_LC_14_31_2 .C_ON=1'b0;
    defparam \c0.data_out_6__3__2193_LC_14_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__3__2193_LC_14_31_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \c0.data_out_6__3__2193_LC_14_31_2  (
            .in0(N__46417),
            .in1(N__38331),
            .in2(N__38317),
            .in3(N__45874),
            .lcout(\c0.data_out_6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50590),
            .ce(N__46130),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__2__2194_LC_14_31_3 .C_ON=1'b0;
    defparam \c0.data_out_6__2__2194_LC_14_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__2__2194_LC_14_31_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_6__2__2194_LC_14_31_3  (
            .in0(N__38298),
            .in1(N__45802),
            .in2(N__38284),
            .in3(N__46419),
            .lcout(\c0.data_out_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50590),
            .ce(N__46130),
            .sr(_gnd_net_));
    defparam \c0.i15246_2_lut_LC_14_31_6 .C_ON=1'b0;
    defparam \c0.i15246_2_lut_LC_14_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15246_2_lut_LC_14_31_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.i15246_2_lut_LC_14_31_6  (
            .in0(N__45801),
            .in1(N__38271),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n17506_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__1__2195_LC_14_31_7 .C_ON=1'b0;
    defparam \c0.data_out_6__1__2195_LC_14_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__1__2195_LC_14_31_7 .LUT_INIT=16'b1111001111010001;
    LogicCell40 \c0.data_out_6__1__2195_LC_14_31_7  (
            .in0(N__42758),
            .in1(N__46418),
            .in2(N__38257),
            .in3(N__52135),
            .lcout(\c0.data_out_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50590),
            .ce(N__46130),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__2__2202_LC_14_32_0 .C_ON=1'b0;
    defparam \c0.data_out_5__2__2202_LC_14_32_0 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__2__2202_LC_14_32_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.data_out_5__2__2202_LC_14_32_0  (
            .in0(N__45994),
            .in1(N__38254),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_out_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50595),
            .ce(N__46129),
            .sr(N__41889));
    defparam \c0.data_out_5__5__2199_LC_14_32_1 .C_ON=1'b0;
    defparam \c0.data_out_5__5__2199_LC_14_32_1 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__5__2199_LC_14_32_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.data_out_5__5__2199_LC_14_32_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38242),
            .in3(N__45992),
            .lcout(\c0.data_out_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50595),
            .ce(N__46129),
            .sr(N__41889));
    defparam \c0.data_out_5__0__2204_LC_14_32_2 .C_ON=1'b0;
    defparam \c0.data_out_5__0__2204_LC_14_32_2 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__0__2204_LC_14_32_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.data_out_5__0__2204_LC_14_32_2  (
            .in0(N__45993),
            .in1(N__38223),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_out_6__1__N_537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50595),
            .ce(N__46129),
            .sr(N__41889));
    defparam \c0.data_out_5__3__2201_LC_14_32_3 .C_ON=1'b0;
    defparam \c0.data_out_5__3__2201_LC_14_32_3 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__3__2201_LC_14_32_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.data_out_5__3__2201_LC_14_32_3  (
            .in0(_gnd_net_),
            .in1(N__45991),
            .in2(_gnd_net_),
            .in3(N__38640),
            .lcout(\c0.data_out_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50595),
            .ce(N__46129),
            .sr(N__41889));
    defparam \c0.data_out_5__4__2200_LC_14_32_4 .C_ON=1'b0;
    defparam \c0.data_out_5__4__2200_LC_14_32_4 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__4__2200_LC_14_32_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.data_out_5__4__2200_LC_14_32_4  (
            .in0(N__45995),
            .in1(N__38625),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_out_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50595),
            .ce(N__46129),
            .sr(N__41889));
    defparam \c0.i1_2_lut_adj_574_LC_15_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_574_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_574_LC_15_18_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_574_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__38611),
            .in2(_gnd_net_),
            .in3(N__38581),
            .lcout(\c0.n9763 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_639_LC_15_19_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_639_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_639_LC_15_19_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_639_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(N__39333),
            .in2(_gnd_net_),
            .in3(N__38523),
            .lcout(\c0.n17037 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_541_LC_15_19_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_541_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_541_LC_15_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_541_LC_15_19_1  (
            .in0(N__39442),
            .in1(N__38485),
            .in2(N__40692),
            .in3(N__43523),
            .lcout(\c0.n17040 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_586_LC_15_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_586_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_586_LC_15_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_586_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__42331),
            .in2(_gnd_net_),
            .in3(N__38469),
            .lcout(\c0.n16933 ),
            .ltout(\c0.n16933_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_591_LC_15_19_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_591_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_591_LC_15_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_591_LC_15_19_3  (
            .in0(N__38415),
            .in1(N__38862),
            .in2(N__38404),
            .in3(N__44242),
            .lcout(\c0.n17_adj_2313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_15_19_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_15_19_6 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_LC_15_19_6  (
            .in0(N__38395),
            .in1(N__51643),
            .in2(N__39244),
            .in3(N__47674),
            .lcout(\c0.n18125 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_611_LC_15_20_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_611_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_611_LC_15_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_611_LC_15_20_0  (
            .in0(N__43216),
            .in1(N__44441),
            .in2(N__38986),
            .in3(N__39593),
            .lcout(),
            .ltout(\c0.n15_adj_2320_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i155_LC_15_20_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i155_LC_15_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i155_LC_15_20_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i155_LC_15_20_1  (
            .in0(N__38839),
            .in1(N__38935),
            .in2(N__38866),
            .in3(N__38863),
            .lcout(\c0.data_out_frame2_19_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50504),
            .ce(N__51168),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_674_LC_15_20_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_674_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_674_LC_15_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_674_LC_15_20_2  (
            .in0(N__43463),
            .in1(N__47200),
            .in2(N__47320),
            .in3(N__49345),
            .lcout(\c0.n14_adj_2323 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_474_LC_15_20_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_474_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_474_LC_15_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_474_LC_15_20_4  (
            .in0(N__38832),
            .in1(N__47505),
            .in2(N__38821),
            .in3(N__40654),
            .lcout(),
            .ltout(\c0.n21_adj_2255_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i164_LC_15_20_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i164_LC_15_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i164_LC_15_20_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.data_out_frame2_0___i164_LC_15_20_5  (
            .in0(N__38806),
            .in1(_gnd_net_),
            .in2(N__38794),
            .in3(N__41788),
            .lcout(\c0.data_out_frame2_20_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50504),
            .ce(N__51168),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i118_LC_15_21_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i118_LC_15_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i118_LC_15_21_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i118_LC_15_21_0  (
            .in0(N__40641),
            .in1(N__38775),
            .in2(_gnd_net_),
            .in3(N__51001),
            .lcout(data_out_frame2_14_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50515),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_478_LC_15_21_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_478_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_478_LC_15_21_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_478_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__42327),
            .in2(_gnd_net_),
            .in3(N__38751),
            .lcout(\c0.n9555 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_503_LC_15_21_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_503_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_503_LC_15_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_503_LC_15_21_4  (
            .in0(N__38734),
            .in1(N__43318),
            .in2(N__38728),
            .in3(N__39385),
            .lcout(\c0.n17103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_LC_15_21_5 .C_ON=1'b0;
    defparam \c0.i13_4_lut_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_LC_15_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_LC_15_21_5  (
            .in0(N__38668),
            .in1(N__41487),
            .in2(N__47484),
            .in3(N__38650),
            .lcout(\c0.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_569_LC_15_21_6 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_569_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_569_LC_15_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_569_LC_15_21_6  (
            .in0(N__39048),
            .in1(N__39022),
            .in2(N__41413),
            .in3(N__47376),
            .lcout(\c0.n19_adj_2303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_609_LC_15_21_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_609_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_609_LC_15_21_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_609_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__41872),
            .in2(_gnd_net_),
            .in3(N__43278),
            .lcout(\c0.n9776 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_465_LC_15_22_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_465_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_465_LC_15_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_465_LC_15_22_0  (
            .in0(N__43411),
            .in1(N__38977),
            .in2(N__43795),
            .in3(N__39494),
            .lcout(),
            .ltout(\c0.n22_adj_2207_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i165_LC_15_22_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i165_LC_15_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i165_LC_15_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i165_LC_15_22_1  (
            .in0(N__41379),
            .in1(N__38965),
            .in2(N__38953),
            .in3(N__38950),
            .lcout(\c0.data_out_frame2_20_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50524),
            .ce(N__50995),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_603_LC_15_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_603_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_603_LC_15_22_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_603_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(N__41135),
            .in2(_gnd_net_),
            .in3(N__42073),
            .lcout(\c0.n9892 ),
            .ltout(\c0.n9892_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_682_LC_15_22_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_682_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_682_LC_15_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_682_LC_15_22_4  (
            .in0(N__39133),
            .in1(N__49427),
            .in2(N__38938),
            .in3(N__44241),
            .lcout(\c0.n17079 ),
            .ltout(\c0.n17079_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i166_LC_15_22_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i166_LC_15_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i166_LC_15_22_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i166_LC_15_22_5  (
            .in0(N__38926),
            .in1(N__41488),
            .in2(N__38917),
            .in3(N__38914),
            .lcout(\c0.data_out_frame2_20_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50524),
            .ce(N__50995),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i94_LC_15_23_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i94_LC_15_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i94_LC_15_23_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i94_LC_15_23_0  (
            .in0(N__50944),
            .in1(N__44568),
            .in2(_gnd_net_),
            .in3(N__41136),
            .lcout(data_out_frame2_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50534),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i88_LC_15_23_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i88_LC_15_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i88_LC_15_23_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i88_LC_15_23_1  (
            .in0(N__44092),
            .in1(N__38891),
            .in2(_gnd_net_),
            .in3(N__50947),
            .lcout(data_out_frame2_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50534),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i45_LC_15_23_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i45_LC_15_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i45_LC_15_23_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i45_LC_15_23_2  (
            .in0(N__50942),
            .in1(N__39214),
            .in2(_gnd_net_),
            .in3(N__43519),
            .lcout(data_out_frame2_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50534),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i79_LC_15_23_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i79_LC_15_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i79_LC_15_23_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i79_LC_15_23_3  (
            .in0(N__48936),
            .in1(N__43472),
            .in2(_gnd_net_),
            .in3(N__50946),
            .lcout(data_out_frame2_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50534),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_597_LC_15_23_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_597_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_597_LC_15_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_597_LC_15_23_4  (
            .in0(N__39163),
            .in1(N__39277),
            .in2(_gnd_net_),
            .in3(N__39132),
            .lcout(\c0.n17082 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i96_LC_15_23_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i96_LC_15_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i96_LC_15_23_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i96_LC_15_23_5  (
            .in0(N__44946),
            .in1(N__41161),
            .in2(_gnd_net_),
            .in3(N__50948),
            .lcout(data_out_frame2_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50534),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i55_LC_15_23_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i55_LC_15_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i55_LC_15_23_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i55_LC_15_23_6  (
            .in0(N__50943),
            .in1(_gnd_net_),
            .in2(N__41217),
            .in3(N__43266),
            .lcout(data_out_frame2_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50534),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i126_LC_15_23_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i126_LC_15_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i126_LC_15_23_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i126_LC_15_23_7  (
            .in0(N__44567),
            .in1(N__49735),
            .in2(_gnd_net_),
            .in3(N__50945),
            .lcout(data_out_frame2_15_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50534),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i50_LC_15_24_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i50_LC_15_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i50_LC_15_24_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i50_LC_15_24_0  (
            .in0(N__39376),
            .in1(N__50930),
            .in2(_gnd_net_),
            .in3(N__41514),
            .lcout(data_out_frame2_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50545),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i53_LC_15_24_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i53_LC_15_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i53_LC_15_24_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i53_LC_15_24_1  (
            .in0(N__50928),
            .in1(_gnd_net_),
            .in2(N__39094),
            .in3(N__39326),
            .lcout(data_out_frame2_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50545),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i61_LC_15_24_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i61_LC_15_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i61_LC_15_24_2 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \c0.data_out_frame2_0___i61_LC_15_24_2  (
            .in0(N__41041),
            .in1(N__50931),
            .in2(N__44173),
            .in3(_gnd_net_),
            .lcout(data_out_frame2_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50545),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_498_LC_15_24_3 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_498_LC_15_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_498_LC_15_24_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_498_LC_15_24_3  (
            .in0(N__39434),
            .in1(N__39396),
            .in2(N__47312),
            .in3(N__49227),
            .lcout(\c0.n25_adj_2275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i114_LC_15_24_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i114_LC_15_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i114_LC_15_24_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i114_LC_15_24_4  (
            .in0(N__39375),
            .in1(N__50929),
            .in2(_gnd_net_),
            .in3(N__49459),
            .lcout(data_out_frame2_14_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50545),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_15_24_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_15_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_15_24_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_15_24_5  (
            .in0(N__48120),
            .in1(N__41040),
            .in2(_gnd_net_),
            .in3(N__39325),
            .lcout(),
            .ltout(\c0.n5_adj_2141_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_15582_LC_15_24_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_15582_LC_15_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_15582_LC_15_24_6 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter2_1__bdd_4_lut_15582_LC_15_24_6  (
            .in0(N__48630),
            .in1(N__43489),
            .in2(N__39304),
            .in3(N__47705),
            .lcout(\c0.n17987 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17951_bdd_4_lut_LC_15_24_7 .C_ON=1'b0;
    defparam \c0.n17951_bdd_4_lut_LC_15_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.n17951_bdd_4_lut_LC_15_24_7 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \c0.n17951_bdd_4_lut_LC_15_24_7  (
            .in0(N__48568),
            .in1(N__39289),
            .in2(N__45361),
            .in3(N__39276),
            .lcout(\c0.n17954 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i70_LC_15_25_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i70_LC_15_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i70_LC_15_25_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i70_LC_15_25_1  (
            .in0(N__41464),
            .in1(N__41867),
            .in2(_gnd_net_),
            .in3(N__50952),
            .lcout(data_out_frame2_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50553),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i74_LC_15_25_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i74_LC_15_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i74_LC_15_25_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i74_LC_15_25_2  (
            .in0(N__50950),
            .in1(_gnd_net_),
            .in2(N__44694),
            .in3(N__41696),
            .lcout(data_out_frame2_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50553),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14884_3_lut_LC_15_25_3 .C_ON=1'b0;
    defparam \c0.i14884_3_lut_LC_15_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14884_3_lut_LC_15_25_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.i14884_3_lut_LC_15_25_3  (
            .in0(N__41956),
            .in1(N__48187),
            .in2(_gnd_net_),
            .in3(N__47372),
            .lcout(\c0.n17322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18053_bdd_4_lut_LC_15_25_5 .C_ON=1'b0;
    defparam \c0.n18053_bdd_4_lut_LC_15_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18053_bdd_4_lut_LC_15_25_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18053_bdd_4_lut_LC_15_25_5  (
            .in0(N__47715),
            .in1(N__39646),
            .in2(N__41764),
            .in3(N__43537),
            .lcout(\c0.n18056 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i57_LC_15_25_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i57_LC_15_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i57_LC_15_25_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i57_LC_15_25_6  (
            .in0(N__50949),
            .in1(N__48768),
            .in2(_gnd_net_),
            .in3(N__39660),
            .lcout(data_out_frame2_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50553),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i105_LC_15_25_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i105_LC_15_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i105_LC_15_25_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i105_LC_15_25_7  (
            .in0(N__41957),
            .in1(N__44784),
            .in2(_gnd_net_),
            .in3(N__50951),
            .lcout(data_out_frame2_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50553),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14908_3_lut_LC_15_26_0 .C_ON=1'b0;
    defparam \c0.i14908_3_lut_LC_15_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14908_3_lut_LC_15_26_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.i14908_3_lut_LC_15_26_0  (
            .in0(N__48164),
            .in1(N__49415),
            .in2(_gnd_net_),
            .in3(N__39477),
            .lcout(\c0.n17346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i107_LC_15_26_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i107_LC_15_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i107_LC_15_26_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i107_LC_15_26_1  (
            .in0(N__39637),
            .in1(N__43372),
            .in2(_gnd_net_),
            .in3(N__51192),
            .lcout(data_out_frame2_13_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50563),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_558_LC_15_26_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_558_LC_15_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_558_LC_15_26_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_558_LC_15_26_2  (
            .in0(_gnd_net_),
            .in1(N__42205),
            .in2(_gnd_net_),
            .in3(N__46199),
            .lcout(\c0.n16918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i115_LC_15_26_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i115_LC_15_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i115_LC_15_26_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i115_LC_15_26_3  (
            .in0(N__44480),
            .in1(N__39576),
            .in2(_gnd_net_),
            .in3(N__51193),
            .lcout(data_out_frame2_14_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50563),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i65_LC_15_26_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i65_LC_15_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i65_LC_15_26_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i65_LC_15_26_5  (
            .in0(N__49416),
            .in1(N__39546),
            .in2(_gnd_net_),
            .in3(N__51194),
            .lcout(data_out_frame2_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50563),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i73_LC_15_26_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i73_LC_15_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i73_LC_15_26_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i73_LC_15_26_6  (
            .in0(N__51191),
            .in1(N__44783),
            .in2(_gnd_net_),
            .in3(N__39478),
            .lcout(data_out_frame2_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50563),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i78_LC_15_26_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i78_LC_15_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i78_LC_15_26_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i78_LC_15_26_7  (
            .in0(N__45293),
            .in1(N__44842),
            .in2(_gnd_net_),
            .in3(N__51195),
            .lcout(data_out_frame2_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50563),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__7__2157_LC_15_27_6 .C_ON=1'b0;
    defparam \c0.data_out_10__7__2157_LC_15_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__7__2157_LC_15_27_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__7__2157_LC_15_27_6  (
            .in0(N__47023),
            .in1(N__46968),
            .in2(N__42982),
            .in3(N__39454),
            .lcout(\c0.data_out_10_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50573),
            .ce(N__46616),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_523_LC_15_28_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_523_LC_15_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_523_LC_15_28_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_523_LC_15_28_1  (
            .in0(N__47096),
            .in1(N__39812),
            .in2(N__39782),
            .in3(N__40056),
            .lcout(\c0.n16966 ),
            .ltout(\c0.n16966_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_530_LC_15_28_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_530_LC_15_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_530_LC_15_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_530_LC_15_28_2  (
            .in0(N__46967),
            .in1(N__45000),
            .in2(N__39745),
            .in3(N__46791),
            .lcout(),
            .ltout(\c0.n10_adj_2288_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_531_LC_15_28_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_531_LC_15_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_531_LC_15_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_531_LC_15_28_3  (
            .in0(N__39742),
            .in1(N__45144),
            .in2(N__39733),
            .in3(N__47004),
            .lcout(\c0.n17109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_552_LC_15_28_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_552_LC_15_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_552_LC_15_28_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_552_LC_15_28_5  (
            .in0(_gnd_net_),
            .in1(N__39720),
            .in2(_gnd_net_),
            .in3(N__39934),
            .lcout(\c0.n17070 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_15_28_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_15_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_15_28_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_15_28_6  (
            .in0(N__52066),
            .in1(N__45022),
            .in2(_gnd_net_),
            .in3(N__43020),
            .lcout(\c0.n8_adj_2153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_545_LC_15_28_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_545_LC_15_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_545_LC_15_28_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_545_LC_15_28_7  (
            .in0(_gnd_net_),
            .in1(N__39704),
            .in2(_gnd_net_),
            .in3(N__46966),
            .lcout(\c0.n17007 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_688_LC_15_29_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_688_LC_15_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_688_LC_15_29_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_688_LC_15_29_0  (
            .in0(N__40079),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40026),
            .lcout(\c0.n16949 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_15_29_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_15_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_15_29_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_15_29_1  (
            .in0(N__39932),
            .in1(N__40078),
            .in2(_gnd_net_),
            .in3(N__52082),
            .lcout(\c0.n8_adj_2166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_LC_15_29_2.C_ON=1'b0;
    defparam i1_2_lut_3_lut_LC_15_29_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_LC_15_29_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 i1_2_lut_3_lut_LC_15_29_2 (
            .in0(N__45930),
            .in1(N__42647),
            .in2(_gnd_net_),
            .in3(N__46475),
            .lcout(n4445),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__5__2175_LC_15_29_3 .C_ON=1'b0;
    defparam \c0.data_out_8__5__2175_LC_15_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__5__2175_LC_15_29_3 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_out_8__5__2175_LC_15_29_3  (
            .in0(N__42648),
            .in1(N__40105),
            .in2(N__42860),
            .in3(N__40080),
            .lcout(data_out_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50587),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_509_LC_15_29_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_509_LC_15_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_509_LC_15_29_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_509_LC_15_29_4  (
            .in0(N__42402),
            .in1(N__39933),
            .in2(N__40429),
            .in3(N__42466),
            .lcout(\c0.n19_adj_2283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_557_LC_15_29_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_557_LC_15_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_557_LC_15_29_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_557_LC_15_29_5  (
            .in0(N__39858),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43013),
            .lcout(\c0.n28_adj_2287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__6__2174_LC_15_29_6 .C_ON=1'b0;
    defparam \c0.data_out_8__6__2174_LC_15_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__6__2174_LC_15_29_6 .LUT_INIT=16'b1111101100001000;
    LogicCell40 \c0.data_out_8__6__2174_LC_15_29_6  (
            .in0(N__40045),
            .in1(N__42842),
            .in2(N__42708),
            .in3(N__40027),
            .lcout(data_out_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50587),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_529_LC_15_29_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_529_LC_15_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_529_LC_15_29_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_529_LC_15_29_7  (
            .in0(N__46822),
            .in1(N__39993),
            .in2(_gnd_net_),
            .in3(N__40425),
            .lcout(\c0.n17043 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_15_30_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_15_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_15_30_0 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_15_30_0  (
            .in0(N__52088),
            .in1(N__39976),
            .in2(N__39838),
            .in3(N__52288),
            .lcout(n10_adj_2425),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__5__2167_LC_15_30_2 .C_ON=1'b0;
    defparam \c0.data_out_9__5__2167_LC_15_30_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__5__2167_LC_15_30_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_9__5__2167_LC_15_30_2  (
            .in0(N__39837),
            .in1(N__39958),
            .in2(N__44973),
            .in3(N__40552),
            .lcout(\c0.data_out_9_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50591),
            .ce(N__46606),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__5__2159_LC_15_30_5 .C_ON=1'b0;
    defparam \c0.data_out_10__5__2159_LC_15_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__5__2159_LC_15_30_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__5__2159_LC_15_30_5  (
            .in0(N__42253),
            .in1(N__42202),
            .in2(N__39916),
            .in3(N__39876),
            .lcout(\c0.data_out_10_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50591),
            .ce(N__46606),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_553_LC_15_31_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_553_LC_15_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_553_LC_15_31_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_553_LC_15_31_2  (
            .in0(N__42228),
            .in1(N__40455),
            .in2(N__45214),
            .in3(N__52131),
            .lcout(\c0.n17025 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__1__2179_LC_15_31_3 .C_ON=1'b0;
    defparam \c0.data_out_8__1__2179_LC_15_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__1__2179_LC_15_31_3 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \c0.data_out_8__1__2179_LC_15_31_3  (
            .in0(N__40385),
            .in1(N__40573),
            .in2(N__42862),
            .in3(N__42759),
            .lcout(data_out_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50596),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_521_LC_15_31_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_521_LC_15_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_521_LC_15_31_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_521_LC_15_31_4  (
            .in0(N__40551),
            .in1(N__40259),
            .in2(N__40525),
            .in3(N__40454),
            .lcout(\c0.n9522 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_31_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_31_5 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_31_5  (
            .in0(N__40384),
            .in1(N__43112),
            .in2(N__52081),
            .in3(N__42921),
            .lcout(\c0.n18077 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15213_3_lut_4_lut_LC_15_32_0 .C_ON=1'b0;
    defparam \c0.i15213_3_lut_4_lut_LC_15_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15213_3_lut_4_lut_LC_15_32_0 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \c0.i15213_3_lut_4_lut_LC_15_32_0  (
            .in0(N__42653),
            .in1(N__40340),
            .in2(N__40188),
            .in3(N__45075),
            .lcout(),
            .ltout(\c0.n17532_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__7__2189_LC_15_32_1 .C_ON=1'b0;
    defparam \c0.data_out_6__7__2189_LC_15_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__7__2189_LC_15_32_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_6__7__2189_LC_15_32_1  (
            .in0(N__40294),
            .in1(N__45996),
            .in2(N__40273),
            .in3(N__46490),
            .lcout(\c0.data_out_6_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50599),
            .ce(N__46128),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_538_LC_15_32_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_538_LC_15_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_538_LC_15_32_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_538_LC_15_32_4  (
            .in0(_gnd_net_),
            .in1(N__42439),
            .in2(_gnd_net_),
            .in3(N__42371),
            .lcout(\c0.n9737 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15255_3_lut_4_lut_LC_15_32_6 .C_ON=1'b0;
    defparam \c0.i15255_3_lut_4_lut_LC_15_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15255_3_lut_4_lut_LC_15_32_6 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \c0.i15255_3_lut_4_lut_LC_15_32_6  (
            .in0(N__42652),
            .in1(N__40219),
            .in2(N__40187),
            .in3(N__45074),
            .lcout(\c0.n17534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15543_LC_16_18_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15543_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15543_LC_16_18_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15543_LC_16_18_1  (
            .in0(N__40669),
            .in1(N__48535),
            .in2(N__40924),
            .in3(N__48105),
            .lcout(\c0.n17999 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15284_3_lut_LC_16_19_2 .C_ON=1'b0;
    defparam \c0.i15284_3_lut_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15284_3_lut_LC_16_19_2 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \c0.i15284_3_lut_LC_16_19_2  (
            .in0(N__40153),
            .in1(N__48624),
            .in2(_gnd_net_),
            .in3(N__48106),
            .lcout(\c0.n17576 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_628_LC_16_19_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_628_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_628_LC_16_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_628_LC_16_19_3  (
            .in0(N__41347),
            .in1(N__44200),
            .in2(_gnd_net_),
            .in3(N__40729),
            .lcout(\c0.n9826 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_608_LC_16_20_0 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_608_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_608_LC_16_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_608_LC_16_20_0  (
            .in0(N__43848),
            .in1(N__43373),
            .in2(N__49855),
            .in3(N__49379),
            .lcout(\c0.n17016 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_601_LC_16_20_1 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_601_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_601_LC_16_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_601_LC_16_20_1  (
            .in0(N__43231),
            .in1(N__44044),
            .in2(N__40696),
            .in3(N__44887),
            .lcout(\c0.n25_adj_2316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i151_LC_16_20_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i151_LC_16_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i151_LC_16_20_2 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.data_out_frame2_0___i151_LC_16_20_2  (
            .in0(N__49917),
            .in1(N__40668),
            .in2(N__51248),
            .in3(_gnd_net_),
            .lcout(data_out_frame2_18_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50516),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_621_LC_16_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_621_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_621_LC_16_20_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_621_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(N__41832),
            .in2(_gnd_net_),
            .in3(N__44632),
            .lcout(\c0.n9843 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_516_LC_16_20_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_516_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_516_LC_16_20_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_516_LC_16_20_5  (
            .in0(N__44356),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43959),
            .lcout(\c0.n16994 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i54_LC_16_20_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i54_LC_16_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i54_LC_16_20_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \c0.data_out_frame2_0___i54_LC_16_20_7  (
            .in0(_gnd_net_),
            .in1(N__51170),
            .in2(N__44642),
            .in3(N__40645),
            .lcout(data_out_frame2_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50516),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_3_lut_LC_16_21_0 .C_ON=1'b0;
    defparam \c0.i14_3_lut_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14_3_lut_LC_16_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i14_3_lut_LC_16_21_0  (
            .in0(N__44308),
            .in1(N__40594),
            .in2(_gnd_net_),
            .in3(N__43336),
            .lcout(),
            .ltout(\c0.n32_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i160_LC_16_21_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i160_LC_16_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i160_LC_16_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i160_LC_16_21_1  (
            .in0(N__41353),
            .in1(N__41005),
            .in2(N__40582),
            .in3(N__40579),
            .lcout(\c0.data_out_frame2_19_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50525),
            .ce(N__51169),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_559_LC_16_21_2 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_559_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_559_LC_16_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_559_LC_16_21_2  (
            .in0(N__44735),
            .in1(N__43279),
            .in2(N__44443),
            .in3(N__49003),
            .lcout(\c0.n29_adj_2296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_598_LC_16_21_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_598_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_598_LC_16_21_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_598_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(N__41596),
            .in2(_gnd_net_),
            .in3(N__44734),
            .lcout(\c0.n16915 ),
            .ltout(\c0.n16915_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_568_LC_16_21_4 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_568_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_568_LC_16_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_568_LC_16_21_4  (
            .in0(N__40999),
            .in1(N__49629),
            .in2(N__40987),
            .in3(N__40984),
            .lcout(),
            .ltout(\c0.n20_adj_2302_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i159_LC_16_21_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i159_LC_16_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i159_LC_16_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_out_frame2_0___i159_LC_16_21_5  (
            .in0(_gnd_net_),
            .in1(N__40942),
            .in2(N__40936),
            .in3(N__40933),
            .lcout(\c0.data_out_frame2_19_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50525),
            .ce(N__51169),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_673_LC_16_22_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_673_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_673_LC_16_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_673_LC_16_22_0  (
            .in0(N__49576),
            .in1(N__41074),
            .in2(N__44614),
            .in3(N__41049),
            .lcout(\c0.n16972 ),
            .ltout(\c0.n16972_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_505_LC_16_22_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_505_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_505_LC_16_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_505_LC_16_22_1  (
            .in0(N__40912),
            .in1(N__49380),
            .in2(N__40879),
            .in3(N__40876),
            .lcout(\c0.n10_adj_2281 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17969_bdd_4_lut_LC_16_22_2 .C_ON=1'b0;
    defparam \c0.n17969_bdd_4_lut_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.n17969_bdd_4_lut_LC_16_22_2 .LUT_INIT=16'b1010101011100100;
    LogicCell40 \c0.n17969_bdd_4_lut_LC_16_22_2  (
            .in0(N__40813),
            .in1(N__40804),
            .in2(N__44110),
            .in3(N__48625),
            .lcout(),
            .ltout(\c0.n17972_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_16_22_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_16_22_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_16_22_3  (
            .in0(N__47761),
            .in1(N__40753),
            .in2(N__40747),
            .in3(N__47710),
            .lcout(\c0.n22_adj_2355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_555_LC_16_22_4 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_555_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_555_LC_16_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_555_LC_16_22_4  (
            .in0(N__41380),
            .in1(N__43182),
            .in2(N__41623),
            .in3(N__41359),
            .lcout(\c0.n30_adj_2295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_16_22_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_16_22_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_16_22_6  (
            .in0(N__41346),
            .in1(N__48167),
            .in2(_gnd_net_),
            .in3(N__44040),
            .lcout(\c0.n5_adj_2351 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_638_LC_16_23_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_638_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_638_LC_16_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_638_LC_16_23_0  (
            .in0(N__41268),
            .in1(N__42068),
            .in2(_gnd_net_),
            .in3(N__47451),
            .lcout(\c0.n9695 ),
            .ltout(\c0.n9695_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_617_LC_16_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_617_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_617_LC_16_23_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_617_LC_16_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41221),
            .in3(N__41509),
            .lcout(\c0.n6_adj_2325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i87_LC_16_23_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i87_LC_16_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i87_LC_16_23_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i87_LC_16_23_2  (
            .in0(N__51199),
            .in1(N__41218),
            .in2(_gnd_net_),
            .in3(N__42316),
            .lcout(data_out_frame2_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50546),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_634_LC_16_23_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_634_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_634_LC_16_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_634_LC_16_23_3  (
            .in0(N__41158),
            .in1(N__41131),
            .in2(_gnd_net_),
            .in3(N__44221),
            .lcout(\c0.n17019 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_542_LC_16_23_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_542_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_542_LC_16_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_542_LC_16_23_4  (
            .in0(N__41109),
            .in1(N__41086),
            .in2(N__41995),
            .in3(N__42315),
            .lcout(\c0.n10_adj_2292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6319_2_lut_LC_16_23_5 .C_ON=1'b0;
    defparam \c0.i6319_2_lut_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6319_2_lut_LC_16_23_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i6319_2_lut_LC_16_23_5  (
            .in0(N__48614),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48190),
            .lcout(\c0.n8621 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_534_LC_16_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_534_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_534_LC_16_23_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_534_LC_16_23_6  (
            .in0(N__41042),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44605),
            .lcout(\c0.n9913 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i103_LC_16_23_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i103_LC_16_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i103_LC_16_23_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i103_LC_16_23_7  (
            .in0(N__49906),
            .in1(N__43636),
            .in2(_gnd_net_),
            .in3(N__51200),
            .lcout(data_out_frame2_12_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50546),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i80_LC_16_24_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i80_LC_16_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i80_LC_16_24_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i80_LC_16_24_0  (
            .in0(N__51202),
            .in1(N__44013),
            .in2(_gnd_net_),
            .in3(N__44878),
            .lcout(data_out_frame2_9_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50554),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_LC_16_24_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_LC_16_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_LC_16_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_LC_16_24_1  (
            .in0(N__44877),
            .in1(N__47410),
            .in2(N__44852),
            .in3(N__47361),
            .lcout(\c0.n17034 ),
            .ltout(\c0.n17034_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_615_LC_16_24_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_615_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_615_LC_16_24_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_615_LC_16_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41611),
            .in3(N__41398),
            .lcout(\c0.n9688 ),
            .ltout(\c0.n9688_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_618_LC_16_24_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_618_LC_16_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_618_LC_16_24_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_618_LC_16_24_3  (
            .in0(N__43832),
            .in1(N__41595),
            .in2(N__41551),
            .in3(N__41548),
            .lcout(\c0.n17010 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i46_LC_16_24_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i46_LC_16_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i46_LC_16_24_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i46_LC_16_24_4  (
            .in0(N__51201),
            .in1(N__45301),
            .in2(_gnd_net_),
            .in3(N__44610),
            .lcout(data_out_frame2_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50554),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15480_LC_16_24_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15480_LC_16_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15480_LC_16_24_5 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15480_LC_16_24_5  (
            .in0(N__48171),
            .in1(N__41542),
            .in2(N__48653),
            .in3(N__47411),
            .lcout(\c0.n17921 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_514_LC_16_24_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_514_LC_16_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_514_LC_16_24_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_514_LC_16_24_6  (
            .in0(N__41513),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45252),
            .lcout(\c0.n17115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i134_LC_16_24_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i134_LC_16_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i134_LC_16_24_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i134_LC_16_24_7  (
            .in0(N__41399),
            .in1(N__41469),
            .in2(_gnd_net_),
            .in3(N__51203),
            .lcout(data_out_frame2_16_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50554),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_600_LC_16_25_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_600_LC_16_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_600_LC_16_25_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_600_LC_16_25_1  (
            .in0(N__45348),
            .in1(N__41866),
            .in2(N__50644),
            .in3(N__41833),
            .lcout(\c0.n24_adj_2315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_472_LC_16_25_2 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_472_LC_16_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_472_LC_16_25_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_472_LC_16_25_2  (
            .in0(N__45596),
            .in1(N__44841),
            .in2(N__49156),
            .in3(N__42066),
            .lcout(\c0.n20_adj_2252 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14885_3_lut_LC_16_25_3 .C_ON=1'b0;
    defparam \c0.i14885_3_lut_LC_16_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14885_3_lut_LC_16_25_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i14885_3_lut_LC_16_25_3  (
            .in0(N__49365),
            .in1(N__42023),
            .in2(_gnd_net_),
            .in3(N__48188),
            .lcout(),
            .ltout(\c0.n17323_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_LC_16_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_LC_16_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_LC_16_25_4 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter2_1__bdd_4_lut_LC_16_25_4  (
            .in0(N__48655),
            .in1(N__41773),
            .in2(N__41767),
            .in3(N__47714),
            .lcout(\c0.n18053 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i121_LC_16_25_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i121_LC_16_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i121_LC_16_25_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \c0.data_out_frame2_0___i121_LC_16_25_5  (
            .in0(_gnd_net_),
            .in1(N__48766),
            .in2(N__49378),
            .in3(N__51186),
            .lcout(data_out_frame2_15_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50564),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i113_LC_16_25_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i113_LC_16_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i113_LC_16_25_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i113_LC_16_25_6  (
            .in0(N__42024),
            .in1(N__41754),
            .in2(_gnd_net_),
            .in3(N__51190),
            .lcout(data_out_frame2_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50564),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17921_bdd_4_lut_LC_16_25_7 .C_ON=1'b0;
    defparam \c0.n17921_bdd_4_lut_LC_16_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.n17921_bdd_4_lut_LC_16_25_7 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.n17921_bdd_4_lut_LC_16_25_7  (
            .in0(N__41690),
            .in1(N__48654),
            .in2(N__47302),
            .in3(N__41668),
            .lcout(\c0.n17924 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i152_LC_16_26_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i152_LC_16_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i152_LC_16_26_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i152_LC_16_26_0  (
            .in0(N__51187),
            .in1(N__51339),
            .in2(_gnd_net_),
            .in3(N__41647),
            .lcout(data_out_frame2_18_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50574),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15592_LC_16_26_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15592_LC_16_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15592_LC_16_26_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15592_LC_16_26_1  (
            .in0(N__41646),
            .in1(N__48651),
            .in2(N__41638),
            .in3(N__48189),
            .lcout(),
            .ltout(\c0.n18059_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18059_bdd_4_lut_LC_16_26_2 .C_ON=1'b0;
    defparam \c0.n18059_bdd_4_lut_LC_16_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18059_bdd_4_lut_LC_16_26_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n18059_bdd_4_lut_LC_16_26_2  (
            .in0(N__48652),
            .in1(N__42033),
            .in2(N__42094),
            .in3(N__50637),
            .lcout(),
            .ltout(\c0.n18062_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_16_26_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_16_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_16_26_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_16_26_3  (
            .in0(N__42091),
            .in1(N__47787),
            .in2(N__42076),
            .in3(N__47716),
            .lcout(\c0.n22_adj_2352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i93_LC_16_26_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i93_LC_16_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i93_LC_16_26_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i93_LC_16_26_4  (
            .in0(N__51188),
            .in1(N__44165),
            .in2(_gnd_net_),
            .in3(N__42067),
            .lcout(data_out_frame2_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50574),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i144_LC_16_26_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i144_LC_16_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i144_LC_16_26_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i144_LC_16_26_5  (
            .in0(N__42034),
            .in1(N__44945),
            .in2(_gnd_net_),
            .in3(N__51189),
            .lcout(data_out_frame2_17_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50574),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_632_LC_16_26_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_632_LC_16_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_632_LC_16_26_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_632_LC_16_26_6  (
            .in0(_gnd_net_),
            .in1(N__42025),
            .in2(_gnd_net_),
            .in3(N__44395),
            .lcout(\c0.n9853 ),
            .ltout(\c0.n9853_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_633_LC_16_26_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_633_LC_16_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_633_LC_16_26_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_633_LC_16_26_7  (
            .in0(N__41994),
            .in1(N__49854),
            .in2(N__41971),
            .in3(N__41958),
            .lcout(\c0.n17046 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15331_2_lut_LC_16_27_5 .C_ON=1'b0;
    defparam \c0.i15331_2_lut_LC_16_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15331_2_lut_LC_16_27_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i15331_2_lut_LC_16_27_5  (
            .in0(_gnd_net_),
            .in1(N__45378),
            .in2(_gnd_net_),
            .in3(N__52096),
            .lcout(\c0.n17581 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15411_2_lut_3_lut_LC_16_28_0 .C_ON=1'b0;
    defparam \c0.i15411_2_lut_3_lut_LC_16_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15411_2_lut_3_lut_LC_16_28_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \c0.i15411_2_lut_3_lut_LC_16_28_0  (
            .in0(N__45931),
            .in1(N__45435),
            .in2(_gnd_net_),
            .in3(N__46480),
            .lcout(\c0.n10259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_16_28_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_16_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_16_28_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_16_28_1  (
            .in0(N__42289),
            .in1(N__42203),
            .in2(_gnd_net_),
            .in3(N__52084),
            .lcout(\c0.n5_adj_2350 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i10_4_lut_LC_16_28_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i10_4_lut_LC_16_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i10_4_lut_LC_16_28_2 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_3_i10_4_lut_LC_16_28_2  (
            .in0(N__52085),
            .in1(N__42259),
            .in2(N__52300),
            .in3(N__46821),
            .lcout(\c0.n10_adj_2154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_515_LC_16_28_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_515_LC_16_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_515_LC_16_28_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_515_LC_16_28_4  (
            .in0(N__42249),
            .in1(N__42340),
            .in2(N__42238),
            .in3(N__46878),
            .lcout(\c0.n12_adj_2285 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_647_LC_16_28_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_647_LC_16_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_647_LC_16_28_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_647_LC_16_28_6  (
            .in0(N__42204),
            .in1(N__46820),
            .in2(_gnd_net_),
            .in3(N__46192),
            .lcout(\c0.n17028 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__3__2225_LC_16_29_0 .C_ON=1'b0;
    defparam \c0.data_out_2__3__2225_LC_16_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__3__2225_LC_16_29_0 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \c0.data_out_2__3__2225_LC_16_29_0  (
            .in0(N__42172),
            .in1(N__42710),
            .in2(N__46133),
            .in3(N__46479),
            .lcout(\c0.data_out_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50592),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15290_2_lut_LC_16_29_1 .C_ON=1'b0;
    defparam \c0.i15290_2_lut_LC_16_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15290_2_lut_LC_16_29_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i15290_2_lut_LC_16_29_1  (
            .in0(_gnd_net_),
            .in1(N__52086),
            .in2(_gnd_net_),
            .in3(N__42171),
            .lcout(\c0.n17593 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__4__2216_LC_16_29_3 .C_ON=1'b0;
    defparam \c0.data_out_3__4__2216_LC_16_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__4__2216_LC_16_29_3 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_3__4__2216_LC_16_29_3  (
            .in0(N__45935),
            .in1(N__42910),
            .in2(N__42163),
            .in3(N__45454),
            .lcout(data_out_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50592),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15261_2_lut_LC_16_29_4 .C_ON=1'b0;
    defparam \c0.i15261_2_lut_LC_16_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15261_2_lut_LC_16_29_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.i15261_2_lut_LC_16_29_4  (
            .in0(N__52087),
            .in1(N__42465),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n17546_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15557_LC_16_29_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15557_LC_16_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15557_LC_16_29_5 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15557_LC_16_29_5  (
            .in0(N__42118),
            .in1(N__52461),
            .in2(N__42112),
            .in3(N__52302),
            .lcout(),
            .ltout(\c0.n18017_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18017_bdd_4_lut_LC_16_29_6 .C_ON=1'b0;
    defparam \c0.n18017_bdd_4_lut_LC_16_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.n18017_bdd_4_lut_LC_16_29_6 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18017_bdd_4_lut_LC_16_29_6  (
            .in0(N__52462),
            .in1(N__42109),
            .in2(N__43171),
            .in3(N__43168),
            .lcout(),
            .ltout(\c0.n18020_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_adj_426_LC_16_29_7 .C_ON=1'b0;
    defparam \c0.i24_4_lut_adj_426_LC_16_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_adj_426_LC_16_29_7 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.i24_4_lut_adj_426_LC_16_29_7  (
            .in0(N__43162),
            .in1(N__52463),
            .in2(N__43156),
            .in3(N__43152),
            .lcout(\c0.n10_adj_2155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__1__2171_LC_16_30_3 .C_ON=1'b0;
    defparam \c0.data_out_9__1__2171_LC_16_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__1__2171_LC_16_30_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_9__1__2171_LC_16_30_3  (
            .in0(N__43030),
            .in1(N__43021),
            .in2(_gnd_net_),
            .in3(N__42981),
            .lcout(\c0.data_out_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50597),
            .ce(N__46621),
            .sr(_gnd_net_));
    defparam \c0.i15289_2_lut_LC_16_30_7 .C_ON=1'b0;
    defparam \c0.i15289_2_lut_LC_16_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15289_2_lut_LC_16_30_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15289_2_lut_LC_16_30_7  (
            .in0(_gnd_net_),
            .in1(N__42909),
            .in2(_gnd_net_),
            .in3(N__52083),
            .lcout(\c0.n17591 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__0__2196_LC_16_31_0 .C_ON=1'b0;
    defparam \c0.data_out_6__0__2196_LC_16_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__0__2196_LC_16_31_0 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \c0.data_out_6__0__2196_LC_16_31_0  (
            .in0(N__42883),
            .in1(N__52498),
            .in2(N__46132),
            .in3(N__42851),
            .lcout(data_out_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50600),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15211_3_lut_LC_16_31_3 .C_ON=1'b0;
    defparam \c0.i15211_3_lut_LC_16_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15211_3_lut_LC_16_31_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \c0.i15211_3_lut_LC_16_31_3  (
            .in0(N__42709),
            .in1(N__42468),
            .in2(_gnd_net_),
            .in3(N__42401),
            .lcout(\c0.n17522 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_547_LC_16_31_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_547_LC_16_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_547_LC_16_31_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_547_LC_16_31_6  (
            .in0(_gnd_net_),
            .in1(N__52497),
            .in2(_gnd_net_),
            .in3(N__46690),
            .lcout(\c0.n9783 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15423_4_lut_LC_16_31_7 .C_ON=1'b0;
    defparam \c0.i15423_4_lut_LC_16_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15423_4_lut_LC_16_31_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i15423_4_lut_LC_16_31_7  (
            .in0(_gnd_net_),
            .in1(N__45875),
            .in2(_gnd_net_),
            .in3(N__45456),
            .lcout(n10055),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15587_LC_17_19_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15587_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15587_LC_17_19_0 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15587_LC_17_19_0  (
            .in0(N__42326),
            .in1(N__48104),
            .in2(N__48636),
            .in3(N__44231),
            .lcout(\c0.n18047 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15368_2_lut_LC_17_20_1 .C_ON=1'b0;
    defparam \c0.i15368_2_lut_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15368_2_lut_LC_17_20_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15368_2_lut_LC_17_20_1  (
            .in0(_gnd_net_),
            .in1(N__43525),
            .in2(_gnd_net_),
            .in3(N__48097),
            .lcout(\c0.n17495 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_594_LC_17_20_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_594_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_594_LC_17_20_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_594_LC_17_20_2  (
            .in0(N__43300),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49273),
            .lcout(\c0.n9671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18047_bdd_4_lut_LC_17_20_6 .C_ON=1'b0;
    defparam \c0.n18047_bdd_4_lut_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.n18047_bdd_4_lut_LC_17_20_6 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.n18047_bdd_4_lut_LC_17_20_6  (
            .in0(N__43473),
            .in1(N__48595),
            .in2(N__43305),
            .in3(N__43417),
            .lcout(\c0.n18050 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_502_LC_17_21_3 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_502_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_502_LC_17_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_502_LC_17_21_3  (
            .in0(N__43410),
            .in1(N__43915),
            .in2(N__43387),
            .in3(N__43335),
            .lcout(\c0.n27_adj_2277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i71_LC_17_21_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i71_LC_17_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i71_LC_17_21_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i71_LC_17_21_4  (
            .in0(N__43304),
            .in1(N__49918),
            .in2(_gnd_net_),
            .in3(N__51207),
            .lcout(data_out_frame2_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50535),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_17_21_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_17_21_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_17_21_5  (
            .in0(N__44355),
            .in1(N__43277),
            .in2(_gnd_net_),
            .in3(N__48221),
            .lcout(\c0.n5_adj_2321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15611_LC_17_21_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15611_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15611_LC_17_21_6 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15611_LC_17_21_6  (
            .in0(N__43237),
            .in1(N__51620),
            .in2(N__43597),
            .in3(N__47708),
            .lcout(\c0.n18083 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_548_LC_17_21_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_548_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_548_LC_17_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_548_LC_17_21_7  (
            .in0(N__43227),
            .in1(N__43215),
            .in2(N__45601),
            .in3(N__43204),
            .lcout(\c0.n16960 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_492_LC_17_22_0 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_492_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_492_LC_17_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_492_LC_17_22_0  (
            .in0(N__48865),
            .in1(N__44039),
            .in2(N__43958),
            .in3(N__45597),
            .lcout(\c0.n24_adj_2272 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_463_LC_17_22_1 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_463_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_463_LC_17_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_463_LC_17_22_1  (
            .in0(N__43907),
            .in1(N__43849),
            .in2(N__47248),
            .in3(N__43804),
            .lcout(\c0.n20_adj_2205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18071_bdd_4_lut_LC_17_22_4 .C_ON=1'b0;
    defparam \c0.n18071_bdd_4_lut_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18071_bdd_4_lut_LC_17_22_4 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \c0.n18071_bdd_4_lut_LC_17_22_4  (
            .in0(N__48594),
            .in1(N__43783),
            .in2(N__44283),
            .in3(N__44886),
            .lcout(),
            .ltout(\c0.n18074_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15626_LC_17_22_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15626_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15626_LC_17_22_5 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15626_LC_17_22_5  (
            .in0(N__43696),
            .in1(N__51619),
            .in2(N__43774),
            .in3(N__47709),
            .lcout(\c0.n18089 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15597_LC_17_22_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15597_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15597_LC_17_22_6 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15597_LC_17_22_6  (
            .in0(N__49194),
            .in1(N__44196),
            .in2(N__48637),
            .in3(N__48215),
            .lcout(),
            .ltout(\c0.n18065_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18065_bdd_4_lut_LC_17_22_7 .C_ON=1'b0;
    defparam \c0.n18065_bdd_4_lut_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.n18065_bdd_4_lut_LC_17_22_7 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n18065_bdd_4_lut_LC_17_22_7  (
            .in0(N__43767),
            .in1(N__43732),
            .in2(N__43699),
            .in3(N__48593),
            .lcout(\c0.n18068 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15577_LC_17_23_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15577_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15577_LC_17_23_0 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15577_LC_17_23_0  (
            .in0(N__44393),
            .in1(N__43686),
            .in2(N__48649),
            .in3(N__48214),
            .lcout(),
            .ltout(\c0.n18005_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18005_bdd_4_lut_LC_17_23_1 .C_ON=1'b0;
    defparam \c0.n18005_bdd_4_lut_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18005_bdd_4_lut_LC_17_23_1 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n18005_bdd_4_lut_LC_17_23_1  (
            .in0(N__49659),
            .in1(N__43626),
            .in2(N__43600),
            .in3(N__48623),
            .lcout(\c0.n18008 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14909_3_lut_LC_17_23_2 .C_ON=1'b0;
    defparam \c0.i14909_3_lut_LC_17_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14909_3_lut_LC_17_23_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.i14909_3_lut_LC_17_23_2  (
            .in0(N__49684),
            .in1(N__48213),
            .in2(_gnd_net_),
            .in3(N__43574),
            .lcout(\c0.n17347 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i132_LC_17_23_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i132_LC_17_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i132_LC_17_23_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i132_LC_17_23_3  (
            .in0(N__49813),
            .in1(N__48993),
            .in2(_gnd_net_),
            .in3(N__51205),
            .lcout(data_out_frame2_16_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50555),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i51_LC_17_23_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i51_LC_17_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i51_LC_17_23_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i51_LC_17_23_4  (
            .in0(N__51204),
            .in1(N__44488),
            .in2(_gnd_net_),
            .in3(N__44421),
            .lcout(data_out_frame2_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50555),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_687_LC_17_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_687_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_687_LC_17_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_687_LC_17_23_6  (
            .in0(N__44394),
            .in1(N__44347),
            .in2(_gnd_net_),
            .in3(N__43947),
            .lcout(\c0.n17127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i72_LC_17_23_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i72_LC_17_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i72_LC_17_23_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i72_LC_17_23_7  (
            .in0(N__51338),
            .in1(N__44272),
            .in2(_gnd_net_),
            .in3(N__51206),
            .lcout(data_out_frame2_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50555),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i95_LC_17_24_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i95_LC_17_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i95_LC_17_24_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i95_LC_17_24_1  (
            .in0(N__51128),
            .in1(_gnd_net_),
            .in2(N__49111),
            .in3(N__44230),
            .lcout(data_out_frame2_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50565),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i120_LC_17_24_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i120_LC_17_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i120_LC_17_24_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i120_LC_17_24_2  (
            .in0(N__44090),
            .in1(N__51129),
            .in2(_gnd_net_),
            .in3(N__44195),
            .lcout(data_out_frame2_14_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50565),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i141_LC_17_24_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i141_LC_17_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i141_LC_17_24_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i141_LC_17_24_3  (
            .in0(N__51126),
            .in1(N__44172),
            .in2(_gnd_net_),
            .in3(N__44106),
            .lcout(data_out_frame2_17_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50565),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i56_LC_17_24_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i56_LC_17_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i56_LC_17_24_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i56_LC_17_24_4  (
            .in0(N__44091),
            .in1(N__51131),
            .in2(_gnd_net_),
            .in3(N__44038),
            .lcout(data_out_frame2_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50565),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i48_LC_17_24_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i48_LC_17_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i48_LC_17_24_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i48_LC_17_24_5  (
            .in0(N__51127),
            .in1(N__44014),
            .in2(_gnd_net_),
            .in3(N__43948),
            .lcout(data_out_frame2_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50565),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i128_LC_17_24_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i128_LC_17_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i128_LC_17_24_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i128_LC_17_24_6  (
            .in0(N__44950),
            .in1(N__51130),
            .in2(_gnd_net_),
            .in3(N__49187),
            .lcout(data_out_frame2_15_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50565),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_613_LC_17_24_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_613_LC_17_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_613_LC_17_24_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_613_LC_17_24_7  (
            .in0(_gnd_net_),
            .in1(N__44882),
            .in2(_gnd_net_),
            .in3(N__44853),
            .lcout(\c0.n16926 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i41_LC_17_25_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i41_LC_17_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i41_LC_17_25_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i41_LC_17_25_0  (
            .in0(N__51243),
            .in1(N__44788),
            .in2(_gnd_net_),
            .in3(N__44716),
            .lcout(data_out_frame2_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50575),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i106_LC_17_25_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i106_LC_17_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i106_LC_17_25_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i106_LC_17_25_1  (
            .in0(N__44695),
            .in1(N__49596),
            .in2(_gnd_net_),
            .in3(N__51245),
            .lcout(data_out_frame2_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50575),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_17_25_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_17_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_17_25_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_17_25_2  (
            .in0(N__45617),
            .in1(N__48228),
            .in2(_gnd_net_),
            .in3(N__44647),
            .lcout(),
            .ltout(\c0.n5_adj_2349_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_17_25_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_17_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_17_25_3 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_17_25_3  (
            .in0(N__48229),
            .in1(N__44606),
            .in2(N__44584),
            .in3(N__48650),
            .lcout(\c0.n6_adj_2280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i62_LC_17_25_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i62_LC_17_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i62_LC_17_25_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_out_frame2_0___i62_LC_17_25_4  (
            .in0(N__51244),
            .in1(_gnd_net_),
            .in2(N__45624),
            .in3(N__44569),
            .lcout(data_out_frame2_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50575),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18089_bdd_4_lut_LC_17_25_6 .C_ON=1'b0;
    defparam \c0.n18089_bdd_4_lut_LC_17_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.n18089_bdd_4_lut_LC_17_25_6 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n18089_bdd_4_lut_LC_17_25_6  (
            .in0(N__44518),
            .in1(N__44509),
            .in2(N__44500),
            .in3(N__51621),
            .lcout(\c0.n18092 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_510_LC_17_25_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_510_LC_17_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_510_LC_17_25_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_510_LC_17_25_7  (
            .in0(_gnd_net_),
            .in1(N__45616),
            .in2(_gnd_net_),
            .in3(N__47198),
            .lcout(\c0.n9678 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i7_LC_17_26_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i7_LC_17_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i7_LC_17_26_3 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \c0.tx2.r_Tx_Data_i7_LC_17_26_3  (
            .in0(N__45577),
            .in1(N__51622),
            .in2(N__51775),
            .in3(N__45571),
            .lcout(\c0.tx2.r_Tx_Data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50581),
            .ce(N__51446),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__0__2244_LC_17_27_0 .C_ON=1'b0;
    defparam \c0.data_out_0__0__2244_LC_17_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__0__2244_LC_17_27_0 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_0__0__2244_LC_17_27_0  (
            .in0(N__45986),
            .in1(N__45516),
            .in2(N__45382),
            .in3(N__46491),
            .lcout(data_out_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50588),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i100_LC_17_27_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i100_LC_17_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i100_LC_17_27_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i100_LC_17_27_5  (
            .in0(N__49809),
            .in1(N__45336),
            .in2(_gnd_net_),
            .in3(N__51209),
            .lcout(data_out_frame2_12_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50588),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i110_LC_17_27_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i110_LC_17_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i110_LC_17_27_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i110_LC_17_27_6  (
            .in0(N__51208),
            .in1(N__45300),
            .in2(_gnd_net_),
            .in3(N__45238),
            .lcout(data_out_frame2_13_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50588),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__3__2169_LC_17_28_0 .C_ON=1'b0;
    defparam \c0.data_out_9__3__2169_LC_17_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__3__2169_LC_17_28_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_9__3__2169_LC_17_28_0  (
            .in0(N__45213),
            .in1(N__45151),
            .in2(N__45133),
            .in3(N__45118),
            .lcout(\c0.data_out_9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50593),
            .ce(N__46623),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_543_LC_17_28_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_543_LC_17_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_543_LC_17_28_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_543_LC_17_28_1  (
            .in0(_gnd_net_),
            .in1(N__45020),
            .in2(_gnd_net_),
            .in3(N__45079),
            .lcout(\c0.n17076 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__6__2166_LC_17_28_5 .C_ON=1'b0;
    defparam \c0.data_out_9__6__2166_LC_17_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__6__2166_LC_17_28_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.data_out_9__6__2166_LC_17_28_5  (
            .in0(N__45034),
            .in1(N__45021),
            .in2(_gnd_net_),
            .in3(N__45004),
            .lcout(\c0.data_out_9_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50593),
            .ce(N__46623),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__4__2168_LC_17_29_1 .C_ON=1'b0;
    defparam \c0.data_out_9__4__2168_LC_17_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__4__2168_LC_17_29_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_9__4__2168_LC_17_29_1  (
            .in0(N__44977),
            .in1(N__47029),
            .in2(N__47152),
            .in3(N__52549),
            .lcout(\c0.data_out_9_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50598),
            .ce(N__46624),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_506_LC_17_29_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_506_LC_17_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_506_LC_17_29_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_506_LC_17_29_2  (
            .in0(_gnd_net_),
            .in1(N__47097),
            .in2(_gnd_net_),
            .in3(N__47056),
            .lcout(\c0.n17058 ),
            .ltout(\c0.n17058_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_511_LC_17_29_3 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_511_LC_17_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_511_LC_17_29_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_511_LC_17_29_3  (
            .in0(N__47022),
            .in1(N__46926),
            .in2(N__47011),
            .in3(N__47008),
            .lcout(),
            .ltout(\c0.n21_adj_2284_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__7__2165_LC_17_29_4 .C_ON=1'b0;
    defparam \c0.data_out_9__7__2165_LC_17_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__7__2165_LC_17_29_4 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.data_out_9__7__2165_LC_17_29_4  (
            .in0(N__46993),
            .in1(_gnd_net_),
            .in2(N__46984),
            .in3(N__46981),
            .lcout(\c0.data_out_9_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50598),
            .ce(N__46624),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__3__2161_LC_17_29_6 .C_ON=1'b0;
    defparam \c0.data_out_10__3__2161_LC_17_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__3__2161_LC_17_29_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__3__2161_LC_17_29_6  (
            .in0(N__46927),
            .in1(N__46912),
            .in2(N__46882),
            .in3(N__46867),
            .lcout(\c0.data_out_10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50598),
            .ce(N__46624),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__6__2158_LC_17_30_1 .C_ON=1'b0;
    defparam \c0.data_out_10__6__2158_LC_17_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__6__2158_LC_17_30_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__6__2158_LC_17_30_1  (
            .in0(N__46799),
            .in1(N__46755),
            .in2(N__46726),
            .in3(N__46701),
            .lcout(\c0.data_out_10_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50601),
            .ce(N__46622),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__5__2191_LC_17_31_0 .C_ON=1'b0;
    defparam \c0.data_out_6__5__2191_LC_17_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__5__2191_LC_17_31_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_6__5__2191_LC_17_31_0  (
            .in0(N__46519),
            .in1(N__45879),
            .in2(N__46501),
            .in3(N__46423),
            .lcout(\c0.data_out_6_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50602),
            .ce(N__46106),
            .sr(_gnd_net_));
    defparam \c0.i15206_2_lut_LC_17_32_3 .C_ON=1'b0;
    defparam \c0.i15206_2_lut_LC_17_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15206_2_lut_LC_17_32_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15206_2_lut_LC_17_32_3  (
            .in0(N__46024),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45947),
            .lcout(\c0.n17450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17999_bdd_4_lut_LC_18_18_5 .C_ON=1'b0;
    defparam \c0.n17999_bdd_4_lut_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.n17999_bdd_4_lut_LC_18_18_5 .LUT_INIT=16'b1100110011100010;
    LogicCell40 \c0.n17999_bdd_4_lut_LC_18_18_5  (
            .in0(N__49847),
            .in1(N__47830),
            .in2(N__49042),
            .in3(N__48461),
            .lcout(\c0.n18002 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_18_19_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_18_19_2 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_18_19_2  (
            .in0(N__47814),
            .in1(N__47740),
            .in2(N__47734),
            .in3(N__47707),
            .lcout(\c0.n22_adj_2353 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i6_LC_18_20_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i6_LC_18_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i6_LC_18_20_0 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \c0.tx2.r_Tx_Data_i6_LC_18_20_0  (
            .in0(N__47422),
            .in1(N__51651),
            .in2(N__51774),
            .in3(N__47536),
            .lcout(\c0.tx2.r_Tx_Data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50536),
            .ce(N__51462),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_599_LC_18_21_0 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_599_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_599_LC_18_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_599_LC_18_21_0  (
            .in0(N__47518),
            .in1(N__47509),
            .in2(N__47488),
            .in3(N__47458),
            .lcout(\c0.n26_adj_2314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_18_21_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_18_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_18_21_6 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_18_21_6  (
            .in0(N__48166),
            .in1(N__48876),
            .in2(N__47440),
            .in3(N__48604),
            .lcout(),
            .ltout(\c0.n6_adj_2290_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18083_bdd_4_lut_LC_18_21_7 .C_ON=1'b0;
    defparam \c0.n18083_bdd_4_lut_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.n18083_bdd_4_lut_LC_18_21_7 .LUT_INIT=16'b1100110011100010;
    LogicCell40 \c0.n18083_bdd_4_lut_LC_18_21_7  (
            .in0(N__47839),
            .in1(N__47431),
            .in2(N__47425),
            .in3(N__51647),
            .lcout(\c0.n18086 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_614_LC_18_22_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_614_LC_18_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_614_LC_18_22_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_614_LC_18_22_1  (
            .in0(_gnd_net_),
            .in1(N__47416),
            .in2(_gnd_net_),
            .in3(N__47377),
            .lcout(),
            .ltout(\c0.n9895_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_4_lut_LC_18_22_2 .C_ON=1'b0;
    defparam \c0.i8_3_lut_4_lut_LC_18_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_4_lut_LC_18_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_3_lut_4_lut_LC_18_22_2  (
            .in0(N__47301),
            .in1(N__47247),
            .in2(N__47203),
            .in3(N__47199),
            .lcout(),
            .ltout(\c0.n23_adj_2318_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i156_LC_18_22_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i156_LC_18_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i156_LC_18_22_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i156_LC_18_22_3  (
            .in0(N__49144),
            .in1(N__49138),
            .in2(N__49126),
            .in3(N__49123),
            .lcout(\c0.data_out_frame2_19_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50556),
            .ce(N__51216),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i143_LC_18_23_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i143_LC_18_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i143_LC_18_23_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i143_LC_18_23_1  (
            .in0(N__49110),
            .in1(N__49038),
            .in2(_gnd_net_),
            .in3(N__51217),
            .lcout(data_out_frame2_17_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50566),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15500_LC_18_23_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15500_LC_18_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15500_LC_18_23_2 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15500_LC_18_23_2  (
            .in0(N__49755),
            .in1(N__48638),
            .in2(N__48222),
            .in3(N__49024),
            .lcout(),
            .ltout(\c0.n17945_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n17945_bdd_4_lut_LC_18_23_3 .C_ON=1'b0;
    defparam \c0.n17945_bdd_4_lut_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.n17945_bdd_4_lut_LC_18_23_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n17945_bdd_4_lut_LC_18_23_3  (
            .in0(N__48639),
            .in1(N__48780),
            .in2(N__49018),
            .in3(N__48989),
            .lcout(\c0.n17948 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i47_LC_18_23_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i47_LC_18_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i47_LC_18_23_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i47_LC_18_23_7  (
            .in0(N__48940),
            .in1(N__48872),
            .in2(_gnd_net_),
            .in3(N__51218),
            .lcout(data_out_frame2_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50566),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i140_LC_18_24_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i140_LC_18_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i140_LC_18_24_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i140_LC_18_24_0  (
            .in0(N__51219),
            .in1(N__48840),
            .in2(_gnd_net_),
            .in3(N__48781),
            .lcout(data_out_frame2_17_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50576),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i89_LC_18_24_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i89_LC_18_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i89_LC_18_24_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i89_LC_18_24_1  (
            .in0(N__48767),
            .in1(N__49686),
            .in2(_gnd_net_),
            .in3(N__51222),
            .lcout(data_out_frame2_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50576),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15313_3_lut_LC_18_24_2 .C_ON=1'b0;
    defparam \c0.i15313_3_lut_LC_18_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15313_3_lut_LC_18_24_2 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \c0.i15313_3_lut_LC_18_24_2  (
            .in0(N__48701),
            .in1(N__48640),
            .in2(_gnd_net_),
            .in3(N__48212),
            .lcout(\c0.n17563 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i135_LC_18_24_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i135_LC_18_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i135_LC_18_24_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i135_LC_18_24_3  (
            .in0(N__49916),
            .in1(N__49843),
            .in2(_gnd_net_),
            .in3(N__51220),
            .lcout(data_out_frame2_16_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50576),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i148_LC_18_24_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i148_LC_18_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i148_LC_18_24_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i148_LC_18_24_5  (
            .in0(N__49801),
            .in1(N__49756),
            .in2(_gnd_net_),
            .in3(N__51221),
            .lcout(data_out_frame2_18_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50576),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_563_LC_18_24_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_563_LC_18_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_563_LC_18_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_563_LC_18_24_7  (
            .in0(N__49742),
            .in1(N__49685),
            .in2(_gnd_net_),
            .in3(N__49663),
            .lcout(\c0.n16923 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_578_LC_18_25_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_578_LC_18_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_578_LC_18_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_578_LC_18_25_0  (
            .in0(N__50635),
            .in1(N__49595),
            .in2(_gnd_net_),
            .in3(N__49182),
            .lcout(\c0.n9910 ),
            .ltout(\c0.n9910_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_622_LC_18_25_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_622_LC_18_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_622_LC_18_25_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_622_LC_18_25_1  (
            .in0(N__49564),
            .in1(N__49540),
            .in2(N__49507),
            .in3(N__49504),
            .lcout(\c0.n16_adj_2327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_623_LC_18_25_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_623_LC_18_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_623_LC_18_25_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_623_LC_18_25_3  (
            .in0(N__49477),
            .in1(N__49432),
            .in2(N__49384),
            .in3(N__49344),
            .lcout(),
            .ltout(\c0.n17_adj_2328_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i154_LC_18_25_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i154_LC_18_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i154_LC_18_25_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i154_LC_18_25_4  (
            .in0(N__49300),
            .in1(N__49294),
            .in2(N__49237),
            .in3(N__49234),
            .lcout(\c0.data_out_frame2_19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50582),
            .ce(N__51215),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_619_LC_18_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_619_LC_18_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_619_LC_18_25_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_619_LC_18_25_5  (
            .in0(N__49183),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50636),
            .lcout(\c0.n16940 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_18_30_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_18_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_18_30_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_18_30_5  (
            .in0(N__52548),
            .in1(N__52512),
            .in2(_gnd_net_),
            .in3(N__52099),
            .lcout(),
            .ltout(\c0.n5_adj_2265_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_18_30_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_18_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_18_30_6 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_LC_18_30_6  (
            .in0(N__51781),
            .in1(N__52404),
            .in2(N__52306),
            .in3(N__52265),
            .lcout(\c0.n18095 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15367_2_lut_LC_18_31_5 .C_ON=1'b0;
    defparam \c0.i15367_2_lut_LC_18_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15367_2_lut_LC_18_31_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15367_2_lut_LC_18_31_5  (
            .in0(_gnd_net_),
            .in1(N__52141),
            .in2(_gnd_net_),
            .in3(N__52038),
            .lcout(\c0.n17632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i4_LC_19_24_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i4_LC_19_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i4_LC_19_24_3 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \c0.tx2.r_Tx_Data_i4_LC_19_24_3  (
            .in0(N__51770),
            .in1(N__51670),
            .in2(N__51655),
            .in3(N__51496),
            .lcout(\c0.tx2.r_Tx_Data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50583),
            .ce(N__51463),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i136_LC_19_26_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i136_LC_19_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i136_LC_19_26_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i136_LC_19_26_5  (
            .in0(N__51346),
            .in1(N__50634),
            .in2(_gnd_net_),
            .in3(N__51272),
            .lcout(data_out_frame2_16_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50594),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
