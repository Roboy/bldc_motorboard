-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Sep 16 2019 18:45:03

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    PIN_9 : in std_logic;
    PIN_8 : in std_logic;
    PIN_7 : in std_logic;
    PIN_6 : inout std_logic;
    PIN_5 : inout std_logic;
    PIN_4 : inout std_logic;
    PIN_3 : out std_logic;
    PIN_24 : out std_logic;
    PIN_23 : out std_logic;
    PIN_22 : out std_logic;
    PIN_21 : in std_logic;
    PIN_20 : in std_logic;
    PIN_2 : out std_logic;
    PIN_19 : in std_logic;
    PIN_18 : in std_logic;
    PIN_17 : in std_logic;
    PIN_16 : in std_logic;
    PIN_15 : in std_logic;
    PIN_14 : in std_logic;
    PIN_13 : in std_logic;
    PIN_12 : in std_logic;
    PIN_11 : inout std_logic;
    PIN_10 : inout std_logic;
    PIN_1 : out std_logic;
    LED : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__73031\ : std_logic;
signal \N__73030\ : std_logic;
signal \N__73029\ : std_logic;
signal \N__73022\ : std_logic;
signal \N__73021\ : std_logic;
signal \N__73020\ : std_logic;
signal \N__73013\ : std_logic;
signal \N__73012\ : std_logic;
signal \N__73011\ : std_logic;
signal \N__73004\ : std_logic;
signal \N__73003\ : std_logic;
signal \N__73002\ : std_logic;
signal \N__72995\ : std_logic;
signal \N__72994\ : std_logic;
signal \N__72993\ : std_logic;
signal \N__72986\ : std_logic;
signal \N__72985\ : std_logic;
signal \N__72984\ : std_logic;
signal \N__72977\ : std_logic;
signal \N__72976\ : std_logic;
signal \N__72975\ : std_logic;
signal \N__72968\ : std_logic;
signal \N__72967\ : std_logic;
signal \N__72966\ : std_logic;
signal \N__72959\ : std_logic;
signal \N__72958\ : std_logic;
signal \N__72957\ : std_logic;
signal \N__72950\ : std_logic;
signal \N__72949\ : std_logic;
signal \N__72948\ : std_logic;
signal \N__72941\ : std_logic;
signal \N__72940\ : std_logic;
signal \N__72939\ : std_logic;
signal \N__72932\ : std_logic;
signal \N__72931\ : std_logic;
signal \N__72930\ : std_logic;
signal \N__72923\ : std_logic;
signal \N__72922\ : std_logic;
signal \N__72921\ : std_logic;
signal \N__72914\ : std_logic;
signal \N__72913\ : std_logic;
signal \N__72912\ : std_logic;
signal \N__72905\ : std_logic;
signal \N__72904\ : std_logic;
signal \N__72903\ : std_logic;
signal \N__72896\ : std_logic;
signal \N__72895\ : std_logic;
signal \N__72894\ : std_logic;
signal \N__72887\ : std_logic;
signal \N__72886\ : std_logic;
signal \N__72885\ : std_logic;
signal \N__72878\ : std_logic;
signal \N__72877\ : std_logic;
signal \N__72876\ : std_logic;
signal \N__72859\ : std_logic;
signal \N__72858\ : std_logic;
signal \N__72855\ : std_logic;
signal \N__72852\ : std_logic;
signal \N__72851\ : std_logic;
signal \N__72848\ : std_logic;
signal \N__72845\ : std_logic;
signal \N__72844\ : std_logic;
signal \N__72841\ : std_logic;
signal \N__72838\ : std_logic;
signal \N__72835\ : std_logic;
signal \N__72834\ : std_logic;
signal \N__72833\ : std_logic;
signal \N__72832\ : std_logic;
signal \N__72831\ : std_logic;
signal \N__72828\ : std_logic;
signal \N__72827\ : std_logic;
signal \N__72824\ : std_logic;
signal \N__72819\ : std_logic;
signal \N__72812\ : std_logic;
signal \N__72809\ : std_logic;
signal \N__72806\ : std_logic;
signal \N__72803\ : std_logic;
signal \N__72800\ : std_logic;
signal \N__72795\ : std_logic;
signal \N__72790\ : std_logic;
signal \N__72781\ : std_logic;
signal \N__72778\ : std_logic;
signal \N__72775\ : std_logic;
signal \N__72774\ : std_logic;
signal \N__72771\ : std_logic;
signal \N__72768\ : std_logic;
signal \N__72767\ : std_logic;
signal \N__72766\ : std_logic;
signal \N__72761\ : std_logic;
signal \N__72756\ : std_logic;
signal \N__72755\ : std_logic;
signal \N__72754\ : std_logic;
signal \N__72749\ : std_logic;
signal \N__72748\ : std_logic;
signal \N__72745\ : std_logic;
signal \N__72744\ : std_logic;
signal \N__72741\ : std_logic;
signal \N__72740\ : std_logic;
signal \N__72739\ : std_logic;
signal \N__72738\ : std_logic;
signal \N__72737\ : std_logic;
signal \N__72734\ : std_logic;
signal \N__72733\ : std_logic;
signal \N__72730\ : std_logic;
signal \N__72729\ : std_logic;
signal \N__72726\ : std_logic;
signal \N__72723\ : std_logic;
signal \N__72720\ : std_logic;
signal \N__72717\ : std_logic;
signal \N__72712\ : std_logic;
signal \N__72711\ : std_logic;
signal \N__72710\ : std_logic;
signal \N__72707\ : std_logic;
signal \N__72704\ : std_logic;
signal \N__72701\ : std_logic;
signal \N__72700\ : std_logic;
signal \N__72699\ : std_logic;
signal \N__72698\ : std_logic;
signal \N__72697\ : std_logic;
signal \N__72694\ : std_logic;
signal \N__72691\ : std_logic;
signal \N__72686\ : std_logic;
signal \N__72681\ : std_logic;
signal \N__72678\ : std_logic;
signal \N__72677\ : std_logic;
signal \N__72674\ : std_logic;
signal \N__72673\ : std_logic;
signal \N__72672\ : std_logic;
signal \N__72669\ : std_logic;
signal \N__72666\ : std_logic;
signal \N__72661\ : std_logic;
signal \N__72660\ : std_logic;
signal \N__72659\ : std_logic;
signal \N__72656\ : std_logic;
signal \N__72653\ : std_logic;
signal \N__72650\ : std_logic;
signal \N__72649\ : std_logic;
signal \N__72646\ : std_logic;
signal \N__72641\ : std_logic;
signal \N__72636\ : std_logic;
signal \N__72633\ : std_logic;
signal \N__72630\ : std_logic;
signal \N__72627\ : std_logic;
signal \N__72622\ : std_logic;
signal \N__72615\ : std_logic;
signal \N__72614\ : std_logic;
signal \N__72613\ : std_logic;
signal \N__72612\ : std_logic;
signal \N__72611\ : std_logic;
signal \N__72610\ : std_logic;
signal \N__72607\ : std_logic;
signal \N__72604\ : std_logic;
signal \N__72601\ : std_logic;
signal \N__72598\ : std_logic;
signal \N__72595\ : std_logic;
signal \N__72592\ : std_logic;
signal \N__72589\ : std_logic;
signal \N__72584\ : std_logic;
signal \N__72575\ : std_logic;
signal \N__72572\ : std_logic;
signal \N__72569\ : std_logic;
signal \N__72566\ : std_logic;
signal \N__72563\ : std_logic;
signal \N__72558\ : std_logic;
signal \N__72549\ : std_logic;
signal \N__72546\ : std_logic;
signal \N__72541\ : std_logic;
signal \N__72538\ : std_logic;
signal \N__72535\ : std_logic;
signal \N__72532\ : std_logic;
signal \N__72531\ : std_logic;
signal \N__72528\ : std_logic;
signal \N__72525\ : std_logic;
signal \N__72522\ : std_logic;
signal \N__72517\ : std_logic;
signal \N__72510\ : std_logic;
signal \N__72505\ : std_logic;
signal \N__72502\ : std_logic;
signal \N__72499\ : std_logic;
signal \N__72496\ : std_logic;
signal \N__72491\ : std_logic;
signal \N__72486\ : std_logic;
signal \N__72475\ : std_logic;
signal \N__72474\ : std_logic;
signal \N__72473\ : std_logic;
signal \N__72468\ : std_logic;
signal \N__72467\ : std_logic;
signal \N__72466\ : std_logic;
signal \N__72463\ : std_logic;
signal \N__72460\ : std_logic;
signal \N__72455\ : std_logic;
signal \N__72452\ : std_logic;
signal \N__72449\ : std_logic;
signal \N__72446\ : std_logic;
signal \N__72439\ : std_logic;
signal \N__72438\ : std_logic;
signal \N__72437\ : std_logic;
signal \N__72434\ : std_logic;
signal \N__72429\ : std_logic;
signal \N__72426\ : std_logic;
signal \N__72425\ : std_logic;
signal \N__72424\ : std_logic;
signal \N__72421\ : std_logic;
signal \N__72418\ : std_logic;
signal \N__72415\ : std_logic;
signal \N__72412\ : std_logic;
signal \N__72409\ : std_logic;
signal \N__72404\ : std_logic;
signal \N__72397\ : std_logic;
signal \N__72394\ : std_logic;
signal \N__72393\ : std_logic;
signal \N__72392\ : std_logic;
signal \N__72389\ : std_logic;
signal \N__72386\ : std_logic;
signal \N__72385\ : std_logic;
signal \N__72382\ : std_logic;
signal \N__72379\ : std_logic;
signal \N__72376\ : std_logic;
signal \N__72373\ : std_logic;
signal \N__72370\ : std_logic;
signal \N__72369\ : std_logic;
signal \N__72366\ : std_logic;
signal \N__72359\ : std_logic;
signal \N__72356\ : std_logic;
signal \N__72349\ : std_logic;
signal \N__72346\ : std_logic;
signal \N__72343\ : std_logic;
signal \N__72342\ : std_logic;
signal \N__72339\ : std_logic;
signal \N__72338\ : std_logic;
signal \N__72337\ : std_logic;
signal \N__72336\ : std_logic;
signal \N__72335\ : std_logic;
signal \N__72332\ : std_logic;
signal \N__72329\ : std_logic;
signal \N__72324\ : std_logic;
signal \N__72319\ : std_logic;
signal \N__72316\ : std_logic;
signal \N__72309\ : std_logic;
signal \N__72304\ : std_logic;
signal \N__72301\ : std_logic;
signal \N__72298\ : std_logic;
signal \N__72295\ : std_logic;
signal \N__72294\ : std_logic;
signal \N__72293\ : std_logic;
signal \N__72292\ : std_logic;
signal \N__72291\ : std_logic;
signal \N__72288\ : std_logic;
signal \N__72287\ : std_logic;
signal \N__72286\ : std_logic;
signal \N__72285\ : std_logic;
signal \N__72284\ : std_logic;
signal \N__72283\ : std_logic;
signal \N__72280\ : std_logic;
signal \N__72277\ : std_logic;
signal \N__72274\ : std_logic;
signal \N__72271\ : std_logic;
signal \N__72270\ : std_logic;
signal \N__72267\ : std_logic;
signal \N__72262\ : std_logic;
signal \N__72261\ : std_logic;
signal \N__72260\ : std_logic;
signal \N__72257\ : std_logic;
signal \N__72256\ : std_logic;
signal \N__72255\ : std_logic;
signal \N__72254\ : std_logic;
signal \N__72251\ : std_logic;
signal \N__72248\ : std_logic;
signal \N__72243\ : std_logic;
signal \N__72242\ : std_logic;
signal \N__72241\ : std_logic;
signal \N__72238\ : std_logic;
signal \N__72235\ : std_logic;
signal \N__72232\ : std_logic;
signal \N__72231\ : std_logic;
signal \N__72228\ : std_logic;
signal \N__72225\ : std_logic;
signal \N__72222\ : std_logic;
signal \N__72221\ : std_logic;
signal \N__72218\ : std_logic;
signal \N__72217\ : std_logic;
signal \N__72214\ : std_logic;
signal \N__72211\ : std_logic;
signal \N__72208\ : std_logic;
signal \N__72207\ : std_logic;
signal \N__72206\ : std_logic;
signal \N__72205\ : std_logic;
signal \N__72202\ : std_logic;
signal \N__72201\ : std_logic;
signal \N__72200\ : std_logic;
signal \N__72199\ : std_logic;
signal \N__72196\ : std_logic;
signal \N__72193\ : std_logic;
signal \N__72190\ : std_logic;
signal \N__72187\ : std_logic;
signal \N__72184\ : std_logic;
signal \N__72181\ : std_logic;
signal \N__72178\ : std_logic;
signal \N__72175\ : std_logic;
signal \N__72172\ : std_logic;
signal \N__72165\ : std_logic;
signal \N__72162\ : std_logic;
signal \N__72159\ : std_logic;
signal \N__72156\ : std_logic;
signal \N__72153\ : std_logic;
signal \N__72150\ : std_logic;
signal \N__72149\ : std_logic;
signal \N__72146\ : std_logic;
signal \N__72145\ : std_logic;
signal \N__72144\ : std_logic;
signal \N__72141\ : std_logic;
signal \N__72136\ : std_logic;
signal \N__72133\ : std_logic;
signal \N__72132\ : std_logic;
signal \N__72129\ : std_logic;
signal \N__72128\ : std_logic;
signal \N__72125\ : std_logic;
signal \N__72122\ : std_logic;
signal \N__72117\ : std_logic;
signal \N__72114\ : std_logic;
signal \N__72105\ : std_logic;
signal \N__72100\ : std_logic;
signal \N__72097\ : std_logic;
signal \N__72092\ : std_logic;
signal \N__72085\ : std_logic;
signal \N__72082\ : std_logic;
signal \N__72079\ : std_logic;
signal \N__72074\ : std_logic;
signal \N__72071\ : std_logic;
signal \N__72066\ : std_logic;
signal \N__72059\ : std_logic;
signal \N__72054\ : std_logic;
signal \N__72051\ : std_logic;
signal \N__72046\ : std_logic;
signal \N__72043\ : std_logic;
signal \N__72036\ : std_logic;
signal \N__72031\ : std_logic;
signal \N__72024\ : std_logic;
signal \N__72019\ : std_logic;
signal \N__72014\ : std_logic;
signal \N__72009\ : std_logic;
signal \N__71998\ : std_logic;
signal \N__71995\ : std_logic;
signal \N__71994\ : std_logic;
signal \N__71993\ : std_logic;
signal \N__71992\ : std_logic;
signal \N__71989\ : std_logic;
signal \N__71982\ : std_logic;
signal \N__71977\ : std_logic;
signal \N__71974\ : std_logic;
signal \N__71973\ : std_logic;
signal \N__71972\ : std_logic;
signal \N__71971\ : std_logic;
signal \N__71970\ : std_logic;
signal \N__71969\ : std_logic;
signal \N__71966\ : std_logic;
signal \N__71965\ : std_logic;
signal \N__71964\ : std_logic;
signal \N__71963\ : std_logic;
signal \N__71962\ : std_logic;
signal \N__71961\ : std_logic;
signal \N__71960\ : std_logic;
signal \N__71959\ : std_logic;
signal \N__71958\ : std_logic;
signal \N__71955\ : std_logic;
signal \N__71952\ : std_logic;
signal \N__71949\ : std_logic;
signal \N__71948\ : std_logic;
signal \N__71947\ : std_logic;
signal \N__71942\ : std_logic;
signal \N__71941\ : std_logic;
signal \N__71938\ : std_logic;
signal \N__71935\ : std_logic;
signal \N__71934\ : std_logic;
signal \N__71933\ : std_logic;
signal \N__71932\ : std_logic;
signal \N__71929\ : std_logic;
signal \N__71922\ : std_logic;
signal \N__71917\ : std_logic;
signal \N__71912\ : std_logic;
signal \N__71907\ : std_logic;
signal \N__71902\ : std_logic;
signal \N__71899\ : std_logic;
signal \N__71898\ : std_logic;
signal \N__71895\ : std_logic;
signal \N__71890\ : std_logic;
signal \N__71883\ : std_logic;
signal \N__71876\ : std_logic;
signal \N__71871\ : std_logic;
signal \N__71870\ : std_logic;
signal \N__71869\ : std_logic;
signal \N__71868\ : std_logic;
signal \N__71863\ : std_logic;
signal \N__71860\ : std_logic;
signal \N__71857\ : std_logic;
signal \N__71854\ : std_logic;
signal \N__71851\ : std_logic;
signal \N__71846\ : std_logic;
signal \N__71839\ : std_logic;
signal \N__71836\ : std_logic;
signal \N__71833\ : std_logic;
signal \N__71830\ : std_logic;
signal \N__71825\ : std_logic;
signal \N__71822\ : std_logic;
signal \N__71817\ : std_logic;
signal \N__71806\ : std_logic;
signal \N__71803\ : std_logic;
signal \N__71802\ : std_logic;
signal \N__71801\ : std_logic;
signal \N__71800\ : std_logic;
signal \N__71797\ : std_logic;
signal \N__71794\ : std_logic;
signal \N__71793\ : std_logic;
signal \N__71792\ : std_logic;
signal \N__71791\ : std_logic;
signal \N__71788\ : std_logic;
signal \N__71787\ : std_logic;
signal \N__71786\ : std_logic;
signal \N__71783\ : std_logic;
signal \N__71782\ : std_logic;
signal \N__71781\ : std_logic;
signal \N__71780\ : std_logic;
signal \N__71779\ : std_logic;
signal \N__71778\ : std_logic;
signal \N__71777\ : std_logic;
signal \N__71776\ : std_logic;
signal \N__71775\ : std_logic;
signal \N__71770\ : std_logic;
signal \N__71767\ : std_logic;
signal \N__71766\ : std_logic;
signal \N__71763\ : std_logic;
signal \N__71762\ : std_logic;
signal \N__71759\ : std_logic;
signal \N__71756\ : std_logic;
signal \N__71755\ : std_logic;
signal \N__71754\ : std_logic;
signal \N__71749\ : std_logic;
signal \N__71746\ : std_logic;
signal \N__71745\ : std_logic;
signal \N__71744\ : std_logic;
signal \N__71741\ : std_logic;
signal \N__71740\ : std_logic;
signal \N__71739\ : std_logic;
signal \N__71738\ : std_logic;
signal \N__71735\ : std_logic;
signal \N__71734\ : std_logic;
signal \N__71729\ : std_logic;
signal \N__71726\ : std_logic;
signal \N__71723\ : std_logic;
signal \N__71718\ : std_logic;
signal \N__71713\ : std_logic;
signal \N__71710\ : std_logic;
signal \N__71707\ : std_logic;
signal \N__71704\ : std_logic;
signal \N__71701\ : std_logic;
signal \N__71698\ : std_logic;
signal \N__71693\ : std_logic;
signal \N__71688\ : std_logic;
signal \N__71681\ : std_logic;
signal \N__71678\ : std_logic;
signal \N__71671\ : std_logic;
signal \N__71668\ : std_logic;
signal \N__71665\ : std_logic;
signal \N__71662\ : std_logic;
signal \N__71659\ : std_logic;
signal \N__71656\ : std_logic;
signal \N__71653\ : std_logic;
signal \N__71650\ : std_logic;
signal \N__71647\ : std_logic;
signal \N__71644\ : std_logic;
signal \N__71641\ : std_logic;
signal \N__71636\ : std_logic;
signal \N__71633\ : std_logic;
signal \N__71630\ : std_logic;
signal \N__71625\ : std_logic;
signal \N__71624\ : std_logic;
signal \N__71623\ : std_logic;
signal \N__71620\ : std_logic;
signal \N__71615\ : std_logic;
signal \N__71612\ : std_logic;
signal \N__71607\ : std_logic;
signal \N__71604\ : std_logic;
signal \N__71601\ : std_logic;
signal \N__71594\ : std_logic;
signal \N__71591\ : std_logic;
signal \N__71586\ : std_logic;
signal \N__71583\ : std_logic;
signal \N__71580\ : std_logic;
signal \N__71573\ : std_logic;
signal \N__71570\ : std_logic;
signal \N__71563\ : std_logic;
signal \N__71548\ : std_logic;
signal \N__71547\ : std_logic;
signal \N__71544\ : std_logic;
signal \N__71543\ : std_logic;
signal \N__71540\ : std_logic;
signal \N__71537\ : std_logic;
signal \N__71536\ : std_logic;
signal \N__71535\ : std_logic;
signal \N__71534\ : std_logic;
signal \N__71531\ : std_logic;
signal \N__71528\ : std_logic;
signal \N__71527\ : std_logic;
signal \N__71526\ : std_logic;
signal \N__71525\ : std_logic;
signal \N__71524\ : std_logic;
signal \N__71521\ : std_logic;
signal \N__71518\ : std_logic;
signal \N__71513\ : std_logic;
signal \N__71510\ : std_logic;
signal \N__71507\ : std_logic;
signal \N__71506\ : std_logic;
signal \N__71505\ : std_logic;
signal \N__71504\ : std_logic;
signal \N__71503\ : std_logic;
signal \N__71500\ : std_logic;
signal \N__71497\ : std_logic;
signal \N__71496\ : std_logic;
signal \N__71493\ : std_logic;
signal \N__71492\ : std_logic;
signal \N__71489\ : std_logic;
signal \N__71488\ : std_logic;
signal \N__71487\ : std_logic;
signal \N__71486\ : std_logic;
signal \N__71485\ : std_logic;
signal \N__71480\ : std_logic;
signal \N__71473\ : std_logic;
signal \N__71470\ : std_logic;
signal \N__71467\ : std_logic;
signal \N__71466\ : std_logic;
signal \N__71465\ : std_logic;
signal \N__71464\ : std_logic;
signal \N__71459\ : std_logic;
signal \N__71456\ : std_logic;
signal \N__71453\ : std_logic;
signal \N__71450\ : std_logic;
signal \N__71445\ : std_logic;
signal \N__71442\ : std_logic;
signal \N__71437\ : std_logic;
signal \N__71436\ : std_logic;
signal \N__71433\ : std_logic;
signal \N__71430\ : std_logic;
signal \N__71427\ : std_logic;
signal \N__71420\ : std_logic;
signal \N__71419\ : std_logic;
signal \N__71412\ : std_logic;
signal \N__71409\ : std_logic;
signal \N__71404\ : std_logic;
signal \N__71399\ : std_logic;
signal \N__71394\ : std_logic;
signal \N__71393\ : std_logic;
signal \N__71390\ : std_logic;
signal \N__71385\ : std_logic;
signal \N__71380\ : std_logic;
signal \N__71377\ : std_logic;
signal \N__71376\ : std_logic;
signal \N__71375\ : std_logic;
signal \N__71374\ : std_logic;
signal \N__71369\ : std_logic;
signal \N__71362\ : std_logic;
signal \N__71359\ : std_logic;
signal \N__71356\ : std_logic;
signal \N__71353\ : std_logic;
signal \N__71350\ : std_logic;
signal \N__71349\ : std_logic;
signal \N__71348\ : std_logic;
signal \N__71347\ : std_logic;
signal \N__71344\ : std_logic;
signal \N__71341\ : std_logic;
signal \N__71336\ : std_logic;
signal \N__71333\ : std_logic;
signal \N__71330\ : std_logic;
signal \N__71323\ : std_logic;
signal \N__71320\ : std_logic;
signal \N__71315\ : std_logic;
signal \N__71312\ : std_logic;
signal \N__71307\ : std_logic;
signal \N__71302\ : std_logic;
signal \N__71295\ : std_logic;
signal \N__71284\ : std_logic;
signal \N__71283\ : std_logic;
signal \N__71280\ : std_logic;
signal \N__71277\ : std_logic;
signal \N__71274\ : std_logic;
signal \N__71273\ : std_logic;
signal \N__71270\ : std_logic;
signal \N__71267\ : std_logic;
signal \N__71266\ : std_logic;
signal \N__71265\ : std_logic;
signal \N__71262\ : std_logic;
signal \N__71259\ : std_logic;
signal \N__71256\ : std_logic;
signal \N__71251\ : std_logic;
signal \N__71248\ : std_logic;
signal \N__71245\ : std_logic;
signal \N__71240\ : std_logic;
signal \N__71233\ : std_logic;
signal \N__71232\ : std_logic;
signal \N__71231\ : std_logic;
signal \N__71230\ : std_logic;
signal \N__71229\ : std_logic;
signal \N__71228\ : std_logic;
signal \N__71227\ : std_logic;
signal \N__71226\ : std_logic;
signal \N__71225\ : std_logic;
signal \N__71224\ : std_logic;
signal \N__71223\ : std_logic;
signal \N__71222\ : std_logic;
signal \N__71221\ : std_logic;
signal \N__71220\ : std_logic;
signal \N__71219\ : std_logic;
signal \N__71218\ : std_logic;
signal \N__71217\ : std_logic;
signal \N__71216\ : std_logic;
signal \N__71215\ : std_logic;
signal \N__71214\ : std_logic;
signal \N__71213\ : std_logic;
signal \N__71212\ : std_logic;
signal \N__71211\ : std_logic;
signal \N__71210\ : std_logic;
signal \N__71209\ : std_logic;
signal \N__71208\ : std_logic;
signal \N__71207\ : std_logic;
signal \N__71206\ : std_logic;
signal \N__71205\ : std_logic;
signal \N__71204\ : std_logic;
signal \N__71203\ : std_logic;
signal \N__71202\ : std_logic;
signal \N__71201\ : std_logic;
signal \N__71200\ : std_logic;
signal \N__71199\ : std_logic;
signal \N__71198\ : std_logic;
signal \N__71197\ : std_logic;
signal \N__71196\ : std_logic;
signal \N__71195\ : std_logic;
signal \N__71194\ : std_logic;
signal \N__71193\ : std_logic;
signal \N__71192\ : std_logic;
signal \N__71191\ : std_logic;
signal \N__71190\ : std_logic;
signal \N__71189\ : std_logic;
signal \N__71188\ : std_logic;
signal \N__71187\ : std_logic;
signal \N__71186\ : std_logic;
signal \N__71185\ : std_logic;
signal \N__71184\ : std_logic;
signal \N__71183\ : std_logic;
signal \N__71182\ : std_logic;
signal \N__71181\ : std_logic;
signal \N__71180\ : std_logic;
signal \N__71179\ : std_logic;
signal \N__71178\ : std_logic;
signal \N__71177\ : std_logic;
signal \N__71176\ : std_logic;
signal \N__71175\ : std_logic;
signal \N__71174\ : std_logic;
signal \N__71173\ : std_logic;
signal \N__71172\ : std_logic;
signal \N__71171\ : std_logic;
signal \N__71170\ : std_logic;
signal \N__71169\ : std_logic;
signal \N__71168\ : std_logic;
signal \N__71167\ : std_logic;
signal \N__71166\ : std_logic;
signal \N__71165\ : std_logic;
signal \N__71164\ : std_logic;
signal \N__71163\ : std_logic;
signal \N__71162\ : std_logic;
signal \N__71161\ : std_logic;
signal \N__71160\ : std_logic;
signal \N__71159\ : std_logic;
signal \N__71158\ : std_logic;
signal \N__71157\ : std_logic;
signal \N__71156\ : std_logic;
signal \N__71155\ : std_logic;
signal \N__71154\ : std_logic;
signal \N__71153\ : std_logic;
signal \N__71152\ : std_logic;
signal \N__71151\ : std_logic;
signal \N__71150\ : std_logic;
signal \N__71149\ : std_logic;
signal \N__71148\ : std_logic;
signal \N__71147\ : std_logic;
signal \N__71146\ : std_logic;
signal \N__71145\ : std_logic;
signal \N__71144\ : std_logic;
signal \N__71143\ : std_logic;
signal \N__71142\ : std_logic;
signal \N__71141\ : std_logic;
signal \N__71140\ : std_logic;
signal \N__71139\ : std_logic;
signal \N__71138\ : std_logic;
signal \N__71137\ : std_logic;
signal \N__71136\ : std_logic;
signal \N__71135\ : std_logic;
signal \N__71134\ : std_logic;
signal \N__71133\ : std_logic;
signal \N__71132\ : std_logic;
signal \N__71131\ : std_logic;
signal \N__71130\ : std_logic;
signal \N__71129\ : std_logic;
signal \N__71128\ : std_logic;
signal \N__71127\ : std_logic;
signal \N__71126\ : std_logic;
signal \N__71125\ : std_logic;
signal \N__71124\ : std_logic;
signal \N__71123\ : std_logic;
signal \N__71122\ : std_logic;
signal \N__71121\ : std_logic;
signal \N__71120\ : std_logic;
signal \N__71119\ : std_logic;
signal \N__71118\ : std_logic;
signal \N__71117\ : std_logic;
signal \N__71116\ : std_logic;
signal \N__71115\ : std_logic;
signal \N__71114\ : std_logic;
signal \N__71113\ : std_logic;
signal \N__71112\ : std_logic;
signal \N__71111\ : std_logic;
signal \N__71110\ : std_logic;
signal \N__71109\ : std_logic;
signal \N__71108\ : std_logic;
signal \N__71107\ : std_logic;
signal \N__71106\ : std_logic;
signal \N__71105\ : std_logic;
signal \N__71104\ : std_logic;
signal \N__71103\ : std_logic;
signal \N__71102\ : std_logic;
signal \N__71101\ : std_logic;
signal \N__71100\ : std_logic;
signal \N__71099\ : std_logic;
signal \N__71098\ : std_logic;
signal \N__71097\ : std_logic;
signal \N__71096\ : std_logic;
signal \N__71095\ : std_logic;
signal \N__71094\ : std_logic;
signal \N__71093\ : std_logic;
signal \N__71092\ : std_logic;
signal \N__71091\ : std_logic;
signal \N__71090\ : std_logic;
signal \N__71089\ : std_logic;
signal \N__71088\ : std_logic;
signal \N__71087\ : std_logic;
signal \N__71086\ : std_logic;
signal \N__71085\ : std_logic;
signal \N__71084\ : std_logic;
signal \N__71083\ : std_logic;
signal \N__71082\ : std_logic;
signal \N__71081\ : std_logic;
signal \N__71080\ : std_logic;
signal \N__71079\ : std_logic;
signal \N__71078\ : std_logic;
signal \N__71077\ : std_logic;
signal \N__71076\ : std_logic;
signal \N__71075\ : std_logic;
signal \N__71074\ : std_logic;
signal \N__71073\ : std_logic;
signal \N__71072\ : std_logic;
signal \N__71071\ : std_logic;
signal \N__71070\ : std_logic;
signal \N__71069\ : std_logic;
signal \N__71068\ : std_logic;
signal \N__71067\ : std_logic;
signal \N__71066\ : std_logic;
signal \N__71065\ : std_logic;
signal \N__71064\ : std_logic;
signal \N__71063\ : std_logic;
signal \N__71062\ : std_logic;
signal \N__71061\ : std_logic;
signal \N__71060\ : std_logic;
signal \N__71059\ : std_logic;
signal \N__71058\ : std_logic;
signal \N__71057\ : std_logic;
signal \N__71056\ : std_logic;
signal \N__71055\ : std_logic;
signal \N__71054\ : std_logic;
signal \N__71053\ : std_logic;
signal \N__71052\ : std_logic;
signal \N__71051\ : std_logic;
signal \N__71050\ : std_logic;
signal \N__71049\ : std_logic;
signal \N__71048\ : std_logic;
signal \N__71047\ : std_logic;
signal \N__71046\ : std_logic;
signal \N__71045\ : std_logic;
signal \N__71044\ : std_logic;
signal \N__71043\ : std_logic;
signal \N__71042\ : std_logic;
signal \N__71041\ : std_logic;
signal \N__71040\ : std_logic;
signal \N__71039\ : std_logic;
signal \N__71038\ : std_logic;
signal \N__71037\ : std_logic;
signal \N__71036\ : std_logic;
signal \N__71035\ : std_logic;
signal \N__71034\ : std_logic;
signal \N__71033\ : std_logic;
signal \N__71032\ : std_logic;
signal \N__71031\ : std_logic;
signal \N__71030\ : std_logic;
signal \N__71029\ : std_logic;
signal \N__71028\ : std_logic;
signal \N__71027\ : std_logic;
signal \N__71026\ : std_logic;
signal \N__71025\ : std_logic;
signal \N__71024\ : std_logic;
signal \N__71023\ : std_logic;
signal \N__71022\ : std_logic;
signal \N__71021\ : std_logic;
signal \N__71020\ : std_logic;
signal \N__71019\ : std_logic;
signal \N__71018\ : std_logic;
signal \N__71017\ : std_logic;
signal \N__71016\ : std_logic;
signal \N__71015\ : std_logic;
signal \N__71014\ : std_logic;
signal \N__71013\ : std_logic;
signal \N__71012\ : std_logic;
signal \N__71011\ : std_logic;
signal \N__71010\ : std_logic;
signal \N__71009\ : std_logic;
signal \N__71008\ : std_logic;
signal \N__71007\ : std_logic;
signal \N__71006\ : std_logic;
signal \N__71005\ : std_logic;
signal \N__71004\ : std_logic;
signal \N__71003\ : std_logic;
signal \N__71002\ : std_logic;
signal \N__71001\ : std_logic;
signal \N__71000\ : std_logic;
signal \N__70999\ : std_logic;
signal \N__70998\ : std_logic;
signal \N__70997\ : std_logic;
signal \N__70996\ : std_logic;
signal \N__70995\ : std_logic;
signal \N__70994\ : std_logic;
signal \N__70993\ : std_logic;
signal \N__70992\ : std_logic;
signal \N__70991\ : std_logic;
signal \N__70504\ : std_logic;
signal \N__70501\ : std_logic;
signal \N__70498\ : std_logic;
signal \N__70495\ : std_logic;
signal \N__70494\ : std_logic;
signal \N__70491\ : std_logic;
signal \N__70488\ : std_logic;
signal \N__70485\ : std_logic;
signal \N__70482\ : std_logic;
signal \N__70481\ : std_logic;
signal \N__70478\ : std_logic;
signal \N__70475\ : std_logic;
signal \N__70472\ : std_logic;
signal \N__70465\ : std_logic;
signal \N__70464\ : std_logic;
signal \N__70461\ : std_logic;
signal \N__70460\ : std_logic;
signal \N__70457\ : std_logic;
signal \N__70456\ : std_logic;
signal \N__70451\ : std_logic;
signal \N__70448\ : std_logic;
signal \N__70445\ : std_logic;
signal \N__70442\ : std_logic;
signal \N__70439\ : std_logic;
signal \N__70438\ : std_logic;
signal \N__70435\ : std_logic;
signal \N__70432\ : std_logic;
signal \N__70429\ : std_logic;
signal \N__70428\ : std_logic;
signal \N__70425\ : std_logic;
signal \N__70420\ : std_logic;
signal \N__70417\ : std_logic;
signal \N__70414\ : std_logic;
signal \N__70405\ : std_logic;
signal \N__70402\ : std_logic;
signal \N__70399\ : std_logic;
signal \N__70396\ : std_logic;
signal \N__70393\ : std_logic;
signal \N__70390\ : std_logic;
signal \N__70389\ : std_logic;
signal \N__70386\ : std_logic;
signal \N__70383\ : std_logic;
signal \N__70382\ : std_logic;
signal \N__70379\ : std_logic;
signal \N__70376\ : std_logic;
signal \N__70375\ : std_logic;
signal \N__70374\ : std_logic;
signal \N__70371\ : std_logic;
signal \N__70368\ : std_logic;
signal \N__70365\ : std_logic;
signal \N__70362\ : std_logic;
signal \N__70359\ : std_logic;
signal \N__70354\ : std_logic;
signal \N__70351\ : std_logic;
signal \N__70348\ : std_logic;
signal \N__70339\ : std_logic;
signal \N__70338\ : std_logic;
signal \N__70337\ : std_logic;
signal \N__70334\ : std_logic;
signal \N__70331\ : std_logic;
signal \N__70328\ : std_logic;
signal \N__70325\ : std_logic;
signal \N__70324\ : std_logic;
signal \N__70321\ : std_logic;
signal \N__70318\ : std_logic;
signal \N__70315\ : std_logic;
signal \N__70314\ : std_logic;
signal \N__70311\ : std_logic;
signal \N__70308\ : std_logic;
signal \N__70303\ : std_logic;
signal \N__70300\ : std_logic;
signal \N__70291\ : std_logic;
signal \N__70288\ : std_logic;
signal \N__70285\ : std_logic;
signal \N__70282\ : std_logic;
signal \N__70279\ : std_logic;
signal \N__70276\ : std_logic;
signal \N__70273\ : std_logic;
signal \N__70270\ : std_logic;
signal \N__70267\ : std_logic;
signal \N__70264\ : std_logic;
signal \N__70261\ : std_logic;
signal \N__70258\ : std_logic;
signal \N__70257\ : std_logic;
signal \N__70254\ : std_logic;
signal \N__70251\ : std_logic;
signal \N__70248\ : std_logic;
signal \N__70243\ : std_logic;
signal \N__70242\ : std_logic;
signal \N__70239\ : std_logic;
signal \N__70236\ : std_logic;
signal \N__70233\ : std_logic;
signal \N__70230\ : std_logic;
signal \N__70225\ : std_logic;
signal \N__70224\ : std_logic;
signal \N__70221\ : std_logic;
signal \N__70218\ : std_logic;
signal \N__70213\ : std_logic;
signal \N__70210\ : std_logic;
signal \N__70209\ : std_logic;
signal \N__70208\ : std_logic;
signal \N__70205\ : std_logic;
signal \N__70202\ : std_logic;
signal \N__70199\ : std_logic;
signal \N__70196\ : std_logic;
signal \N__70189\ : std_logic;
signal \N__70188\ : std_logic;
signal \N__70183\ : std_logic;
signal \N__70180\ : std_logic;
signal \N__70177\ : std_logic;
signal \N__70174\ : std_logic;
signal \N__70171\ : std_logic;
signal \N__70168\ : std_logic;
signal \N__70165\ : std_logic;
signal \N__70162\ : std_logic;
signal \N__70161\ : std_logic;
signal \N__70158\ : std_logic;
signal \N__70155\ : std_logic;
signal \N__70154\ : std_logic;
signal \N__70151\ : std_logic;
signal \N__70148\ : std_logic;
signal \N__70147\ : std_logic;
signal \N__70144\ : std_logic;
signal \N__70139\ : std_logic;
signal \N__70134\ : std_logic;
signal \N__70131\ : std_logic;
signal \N__70126\ : std_logic;
signal \N__70125\ : std_logic;
signal \N__70124\ : std_logic;
signal \N__70123\ : std_logic;
signal \N__70120\ : std_logic;
signal \N__70117\ : std_logic;
signal \N__70114\ : std_logic;
signal \N__70111\ : std_logic;
signal \N__70108\ : std_logic;
signal \N__70105\ : std_logic;
signal \N__70102\ : std_logic;
signal \N__70099\ : std_logic;
signal \N__70096\ : std_logic;
signal \N__70091\ : std_logic;
signal \N__70084\ : std_logic;
signal \N__70083\ : std_logic;
signal \N__70080\ : std_logic;
signal \N__70077\ : std_logic;
signal \N__70074\ : std_logic;
signal \N__70069\ : std_logic;
signal \N__70066\ : std_logic;
signal \N__70063\ : std_logic;
signal \N__70060\ : std_logic;
signal \N__70057\ : std_logic;
signal \N__70056\ : std_logic;
signal \N__70053\ : std_logic;
signal \N__70050\ : std_logic;
signal \N__70045\ : std_logic;
signal \N__70044\ : std_logic;
signal \N__70041\ : std_logic;
signal \N__70038\ : std_logic;
signal \N__70037\ : std_logic;
signal \N__70032\ : std_logic;
signal \N__70029\ : std_logic;
signal \N__70026\ : std_logic;
signal \N__70021\ : std_logic;
signal \N__70018\ : std_logic;
signal \N__70017\ : std_logic;
signal \N__70016\ : std_logic;
signal \N__70013\ : std_logic;
signal \N__70010\ : std_logic;
signal \N__70007\ : std_logic;
signal \N__70004\ : std_logic;
signal \N__70001\ : std_logic;
signal \N__69998\ : std_logic;
signal \N__69991\ : std_logic;
signal \N__69988\ : std_logic;
signal \N__69987\ : std_logic;
signal \N__69986\ : std_logic;
signal \N__69983\ : std_logic;
signal \N__69980\ : std_logic;
signal \N__69977\ : std_logic;
signal \N__69974\ : std_logic;
signal \N__69971\ : std_logic;
signal \N__69968\ : std_logic;
signal \N__69967\ : std_logic;
signal \N__69966\ : std_logic;
signal \N__69965\ : std_logic;
signal \N__69964\ : std_logic;
signal \N__69961\ : std_logic;
signal \N__69958\ : std_logic;
signal \N__69955\ : std_logic;
signal \N__69946\ : std_logic;
signal \N__69937\ : std_logic;
signal \N__69934\ : std_logic;
signal \N__69933\ : std_logic;
signal \N__69930\ : std_logic;
signal \N__69927\ : std_logic;
signal \N__69922\ : std_logic;
signal \N__69919\ : std_logic;
signal \N__69918\ : std_logic;
signal \N__69913\ : std_logic;
signal \N__69910\ : std_logic;
signal \N__69907\ : std_logic;
signal \N__69904\ : std_logic;
signal \N__69903\ : std_logic;
signal \N__69900\ : std_logic;
signal \N__69897\ : std_logic;
signal \N__69896\ : std_logic;
signal \N__69893\ : std_logic;
signal \N__69890\ : std_logic;
signal \N__69889\ : std_logic;
signal \N__69886\ : std_logic;
signal \N__69883\ : std_logic;
signal \N__69880\ : std_logic;
signal \N__69879\ : std_logic;
signal \N__69876\ : std_logic;
signal \N__69873\ : std_logic;
signal \N__69870\ : std_logic;
signal \N__69867\ : std_logic;
signal \N__69862\ : std_logic;
signal \N__69853\ : std_logic;
signal \N__69850\ : std_logic;
signal \N__69849\ : std_logic;
signal \N__69848\ : std_logic;
signal \N__69845\ : std_logic;
signal \N__69840\ : std_logic;
signal \N__69835\ : std_logic;
signal \N__69834\ : std_logic;
signal \N__69831\ : std_logic;
signal \N__69828\ : std_logic;
signal \N__69827\ : std_logic;
signal \N__69826\ : std_logic;
signal \N__69825\ : std_logic;
signal \N__69822\ : std_logic;
signal \N__69819\ : std_logic;
signal \N__69818\ : std_logic;
signal \N__69817\ : std_logic;
signal \N__69812\ : std_logic;
signal \N__69809\ : std_logic;
signal \N__69804\ : std_logic;
signal \N__69801\ : std_logic;
signal \N__69798\ : std_logic;
signal \N__69787\ : std_logic;
signal \N__69784\ : std_logic;
signal \N__69781\ : std_logic;
signal \N__69778\ : std_logic;
signal \N__69777\ : std_logic;
signal \N__69774\ : std_logic;
signal \N__69773\ : std_logic;
signal \N__69772\ : std_logic;
signal \N__69769\ : std_logic;
signal \N__69766\ : std_logic;
signal \N__69761\ : std_logic;
signal \N__69758\ : std_logic;
signal \N__69753\ : std_logic;
signal \N__69748\ : std_logic;
signal \N__69747\ : std_logic;
signal \N__69746\ : std_logic;
signal \N__69745\ : std_logic;
signal \N__69744\ : std_logic;
signal \N__69739\ : std_logic;
signal \N__69734\ : std_logic;
signal \N__69731\ : std_logic;
signal \N__69726\ : std_logic;
signal \N__69723\ : std_logic;
signal \N__69718\ : std_logic;
signal \N__69715\ : std_logic;
signal \N__69714\ : std_logic;
signal \N__69711\ : std_logic;
signal \N__69708\ : std_logic;
signal \N__69707\ : std_logic;
signal \N__69704\ : std_logic;
signal \N__69701\ : std_logic;
signal \N__69698\ : std_logic;
signal \N__69695\ : std_logic;
signal \N__69688\ : std_logic;
signal \N__69685\ : std_logic;
signal \N__69684\ : std_logic;
signal \N__69683\ : std_logic;
signal \N__69682\ : std_logic;
signal \N__69679\ : std_logic;
signal \N__69676\ : std_logic;
signal \N__69673\ : std_logic;
signal \N__69670\ : std_logic;
signal \N__69661\ : std_logic;
signal \N__69658\ : std_logic;
signal \N__69657\ : std_logic;
signal \N__69656\ : std_logic;
signal \N__69653\ : std_logic;
signal \N__69652\ : std_logic;
signal \N__69649\ : std_logic;
signal \N__69648\ : std_logic;
signal \N__69645\ : std_logic;
signal \N__69642\ : std_logic;
signal \N__69637\ : std_logic;
signal \N__69636\ : std_logic;
signal \N__69633\ : std_logic;
signal \N__69630\ : std_logic;
signal \N__69625\ : std_logic;
signal \N__69622\ : std_logic;
signal \N__69619\ : std_logic;
signal \N__69614\ : std_logic;
signal \N__69607\ : std_logic;
signal \N__69606\ : std_logic;
signal \N__69603\ : std_logic;
signal \N__69602\ : std_logic;
signal \N__69599\ : std_logic;
signal \N__69596\ : std_logic;
signal \N__69595\ : std_logic;
signal \N__69592\ : std_logic;
signal \N__69589\ : std_logic;
signal \N__69586\ : std_logic;
signal \N__69583\ : std_logic;
signal \N__69580\ : std_logic;
signal \N__69577\ : std_logic;
signal \N__69572\ : std_logic;
signal \N__69565\ : std_logic;
signal \N__69564\ : std_logic;
signal \N__69561\ : std_logic;
signal \N__69558\ : std_logic;
signal \N__69557\ : std_logic;
signal \N__69556\ : std_logic;
signal \N__69555\ : std_logic;
signal \N__69552\ : std_logic;
signal \N__69547\ : std_logic;
signal \N__69544\ : std_logic;
signal \N__69543\ : std_logic;
signal \N__69540\ : std_logic;
signal \N__69537\ : std_logic;
signal \N__69534\ : std_logic;
signal \N__69529\ : std_logic;
signal \N__69526\ : std_logic;
signal \N__69517\ : std_logic;
signal \N__69514\ : std_logic;
signal \N__69511\ : std_logic;
signal \N__69510\ : std_logic;
signal \N__69509\ : std_logic;
signal \N__69506\ : std_logic;
signal \N__69501\ : std_logic;
signal \N__69496\ : std_logic;
signal \N__69493\ : std_logic;
signal \N__69492\ : std_logic;
signal \N__69489\ : std_logic;
signal \N__69486\ : std_logic;
signal \N__69483\ : std_logic;
signal \N__69480\ : std_logic;
signal \N__69475\ : std_logic;
signal \N__69472\ : std_logic;
signal \N__69469\ : std_logic;
signal \N__69466\ : std_logic;
signal \N__69465\ : std_logic;
signal \N__69462\ : std_logic;
signal \N__69459\ : std_logic;
signal \N__69458\ : std_logic;
signal \N__69455\ : std_logic;
signal \N__69450\ : std_logic;
signal \N__69445\ : std_logic;
signal \N__69444\ : std_logic;
signal \N__69443\ : std_logic;
signal \N__69442\ : std_logic;
signal \N__69439\ : std_logic;
signal \N__69438\ : std_logic;
signal \N__69437\ : std_logic;
signal \N__69436\ : std_logic;
signal \N__69435\ : std_logic;
signal \N__69432\ : std_logic;
signal \N__69429\ : std_logic;
signal \N__69426\ : std_logic;
signal \N__69425\ : std_logic;
signal \N__69424\ : std_logic;
signal \N__69423\ : std_logic;
signal \N__69422\ : std_logic;
signal \N__69421\ : std_logic;
signal \N__69418\ : std_logic;
signal \N__69415\ : std_logic;
signal \N__69414\ : std_logic;
signal \N__69411\ : std_logic;
signal \N__69410\ : std_logic;
signal \N__69409\ : std_logic;
signal \N__69408\ : std_logic;
signal \N__69405\ : std_logic;
signal \N__69402\ : std_logic;
signal \N__69399\ : std_logic;
signal \N__69396\ : std_logic;
signal \N__69393\ : std_logic;
signal \N__69390\ : std_logic;
signal \N__69385\ : std_logic;
signal \N__69382\ : std_logic;
signal \N__69381\ : std_logic;
signal \N__69380\ : std_logic;
signal \N__69377\ : std_logic;
signal \N__69376\ : std_logic;
signal \N__69371\ : std_logic;
signal \N__69364\ : std_logic;
signal \N__69363\ : std_logic;
signal \N__69360\ : std_logic;
signal \N__69357\ : std_logic;
signal \N__69352\ : std_logic;
signal \N__69349\ : std_logic;
signal \N__69342\ : std_logic;
signal \N__69339\ : std_logic;
signal \N__69336\ : std_logic;
signal \N__69331\ : std_logic;
signal \N__69328\ : std_logic;
signal \N__69325\ : std_logic;
signal \N__69320\ : std_logic;
signal \N__69317\ : std_logic;
signal \N__69316\ : std_logic;
signal \N__69315\ : std_logic;
signal \N__69314\ : std_logic;
signal \N__69311\ : std_logic;
signal \N__69308\ : std_logic;
signal \N__69301\ : std_logic;
signal \N__69298\ : std_logic;
signal \N__69293\ : std_logic;
signal \N__69288\ : std_logic;
signal \N__69287\ : std_logic;
signal \N__69284\ : std_logic;
signal \N__69279\ : std_logic;
signal \N__69278\ : std_logic;
signal \N__69277\ : std_logic;
signal \N__69274\ : std_logic;
signal \N__69271\ : std_logic;
signal \N__69264\ : std_logic;
signal \N__69261\ : std_logic;
signal \N__69256\ : std_logic;
signal \N__69253\ : std_logic;
signal \N__69248\ : std_logic;
signal \N__69247\ : std_logic;
signal \N__69242\ : std_logic;
signal \N__69239\ : std_logic;
signal \N__69236\ : std_logic;
signal \N__69233\ : std_logic;
signal \N__69228\ : std_logic;
signal \N__69225\ : std_logic;
signal \N__69222\ : std_logic;
signal \N__69219\ : std_logic;
signal \N__69218\ : std_logic;
signal \N__69217\ : std_logic;
signal \N__69216\ : std_logic;
signal \N__69215\ : std_logic;
signal \N__69212\ : std_logic;
signal \N__69207\ : std_logic;
signal \N__69204\ : std_logic;
signal \N__69201\ : std_logic;
signal \N__69194\ : std_logic;
signal \N__69189\ : std_logic;
signal \N__69184\ : std_logic;
signal \N__69169\ : std_logic;
signal \N__69168\ : std_logic;
signal \N__69167\ : std_logic;
signal \N__69164\ : std_logic;
signal \N__69161\ : std_logic;
signal \N__69158\ : std_logic;
signal \N__69155\ : std_logic;
signal \N__69152\ : std_logic;
signal \N__69151\ : std_logic;
signal \N__69150\ : std_logic;
signal \N__69147\ : std_logic;
signal \N__69146\ : std_logic;
signal \N__69143\ : std_logic;
signal \N__69140\ : std_logic;
signal \N__69139\ : std_logic;
signal \N__69138\ : std_logic;
signal \N__69133\ : std_logic;
signal \N__69130\ : std_logic;
signal \N__69127\ : std_logic;
signal \N__69124\ : std_logic;
signal \N__69121\ : std_logic;
signal \N__69116\ : std_logic;
signal \N__69111\ : std_logic;
signal \N__69108\ : std_logic;
signal \N__69105\ : std_logic;
signal \N__69102\ : std_logic;
signal \N__69097\ : std_logic;
signal \N__69092\ : std_logic;
signal \N__69089\ : std_logic;
signal \N__69082\ : std_logic;
signal \N__69081\ : std_logic;
signal \N__69080\ : std_logic;
signal \N__69079\ : std_logic;
signal \N__69078\ : std_logic;
signal \N__69071\ : std_logic;
signal \N__69066\ : std_logic;
signal \N__69063\ : std_logic;
signal \N__69060\ : std_logic;
signal \N__69057\ : std_logic;
signal \N__69056\ : std_logic;
signal \N__69055\ : std_logic;
signal \N__69050\ : std_logic;
signal \N__69045\ : std_logic;
signal \N__69040\ : std_logic;
signal \N__69037\ : std_logic;
signal \N__69036\ : std_logic;
signal \N__69035\ : std_logic;
signal \N__69032\ : std_logic;
signal \N__69031\ : std_logic;
signal \N__69026\ : std_logic;
signal \N__69025\ : std_logic;
signal \N__69024\ : std_logic;
signal \N__69023\ : std_logic;
signal \N__69022\ : std_logic;
signal \N__69019\ : std_logic;
signal \N__69016\ : std_logic;
signal \N__69015\ : std_logic;
signal \N__69014\ : std_logic;
signal \N__69013\ : std_logic;
signal \N__69012\ : std_logic;
signal \N__69011\ : std_logic;
signal \N__69008\ : std_logic;
signal \N__69007\ : std_logic;
signal \N__69006\ : std_logic;
signal \N__69003\ : std_logic;
signal \N__69002\ : std_logic;
signal \N__69001\ : std_logic;
signal \N__68998\ : std_logic;
signal \N__68995\ : std_logic;
signal \N__68994\ : std_logic;
signal \N__68991\ : std_logic;
signal \N__68986\ : std_logic;
signal \N__68981\ : std_logic;
signal \N__68980\ : std_logic;
signal \N__68977\ : std_logic;
signal \N__68974\ : std_logic;
signal \N__68973\ : std_logic;
signal \N__68970\ : std_logic;
signal \N__68967\ : std_logic;
signal \N__68964\ : std_logic;
signal \N__68961\ : std_logic;
signal \N__68956\ : std_logic;
signal \N__68953\ : std_logic;
signal \N__68950\ : std_logic;
signal \N__68945\ : std_logic;
signal \N__68938\ : std_logic;
signal \N__68935\ : std_logic;
signal \N__68932\ : std_logic;
signal \N__68929\ : std_logic;
signal \N__68928\ : std_logic;
signal \N__68927\ : std_logic;
signal \N__68924\ : std_logic;
signal \N__68923\ : std_logic;
signal \N__68920\ : std_logic;
signal \N__68917\ : std_logic;
signal \N__68912\ : std_logic;
signal \N__68909\ : std_logic;
signal \N__68904\ : std_logic;
signal \N__68903\ : std_logic;
signal \N__68898\ : std_logic;
signal \N__68895\ : std_logic;
signal \N__68890\ : std_logic;
signal \N__68887\ : std_logic;
signal \N__68882\ : std_logic;
signal \N__68879\ : std_logic;
signal \N__68872\ : std_logic;
signal \N__68867\ : std_logic;
signal \N__68866\ : std_logic;
signal \N__68863\ : std_logic;
signal \N__68860\ : std_logic;
signal \N__68855\ : std_logic;
signal \N__68854\ : std_logic;
signal \N__68853\ : std_logic;
signal \N__68850\ : std_logic;
signal \N__68845\ : std_logic;
signal \N__68844\ : std_logic;
signal \N__68843\ : std_logic;
signal \N__68840\ : std_logic;
signal \N__68837\ : std_logic;
signal \N__68834\ : std_logic;
signal \N__68827\ : std_logic;
signal \N__68826\ : std_logic;
signal \N__68825\ : std_logic;
signal \N__68824\ : std_logic;
signal \N__68821\ : std_logic;
signal \N__68818\ : std_logic;
signal \N__68813\ : std_logic;
signal \N__68808\ : std_logic;
signal \N__68803\ : std_logic;
signal \N__68800\ : std_logic;
signal \N__68797\ : std_logic;
signal \N__68794\ : std_logic;
signal \N__68789\ : std_logic;
signal \N__68786\ : std_logic;
signal \N__68781\ : std_logic;
signal \N__68776\ : std_logic;
signal \N__68771\ : std_logic;
signal \N__68758\ : std_logic;
signal \N__68755\ : std_logic;
signal \N__68752\ : std_logic;
signal \N__68751\ : std_logic;
signal \N__68750\ : std_logic;
signal \N__68747\ : std_logic;
signal \N__68746\ : std_logic;
signal \N__68745\ : std_logic;
signal \N__68744\ : std_logic;
signal \N__68741\ : std_logic;
signal \N__68740\ : std_logic;
signal \N__68737\ : std_logic;
signal \N__68734\ : std_logic;
signal \N__68731\ : std_logic;
signal \N__68728\ : std_logic;
signal \N__68727\ : std_logic;
signal \N__68726\ : std_logic;
signal \N__68725\ : std_logic;
signal \N__68724\ : std_logic;
signal \N__68723\ : std_logic;
signal \N__68722\ : std_logic;
signal \N__68719\ : std_logic;
signal \N__68716\ : std_logic;
signal \N__68713\ : std_logic;
signal \N__68712\ : std_logic;
signal \N__68711\ : std_logic;
signal \N__68708\ : std_logic;
signal \N__68701\ : std_logic;
signal \N__68698\ : std_logic;
signal \N__68695\ : std_logic;
signal \N__68692\ : std_logic;
signal \N__68691\ : std_logic;
signal \N__68688\ : std_logic;
signal \N__68683\ : std_logic;
signal \N__68682\ : std_logic;
signal \N__68675\ : std_logic;
signal \N__68674\ : std_logic;
signal \N__68671\ : std_logic;
signal \N__68668\ : std_logic;
signal \N__68657\ : std_logic;
signal \N__68656\ : std_logic;
signal \N__68655\ : std_logic;
signal \N__68652\ : std_logic;
signal \N__68649\ : std_logic;
signal \N__68648\ : std_logic;
signal \N__68647\ : std_logic;
signal \N__68646\ : std_logic;
signal \N__68645\ : std_logic;
signal \N__68644\ : std_logic;
signal \N__68641\ : std_logic;
signal \N__68638\ : std_logic;
signal \N__68635\ : std_logic;
signal \N__68632\ : std_logic;
signal \N__68629\ : std_logic;
signal \N__68626\ : std_logic;
signal \N__68623\ : std_logic;
signal \N__68622\ : std_logic;
signal \N__68619\ : std_logic;
signal \N__68616\ : std_logic;
signal \N__68613\ : std_logic;
signal \N__68612\ : std_logic;
signal \N__68609\ : std_logic;
signal \N__68604\ : std_logic;
signal \N__68601\ : std_logic;
signal \N__68598\ : std_logic;
signal \N__68595\ : std_logic;
signal \N__68594\ : std_logic;
signal \N__68593\ : std_logic;
signal \N__68590\ : std_logic;
signal \N__68587\ : std_logic;
signal \N__68584\ : std_logic;
signal \N__68581\ : std_logic;
signal \N__68576\ : std_logic;
signal \N__68573\ : std_logic;
signal \N__68570\ : std_logic;
signal \N__68565\ : std_logic;
signal \N__68562\ : std_logic;
signal \N__68559\ : std_logic;
signal \N__68554\ : std_logic;
signal \N__68553\ : std_logic;
signal \N__68546\ : std_logic;
signal \N__68543\ : std_logic;
signal \N__68540\ : std_logic;
signal \N__68535\ : std_logic;
signal \N__68532\ : std_logic;
signal \N__68529\ : std_logic;
signal \N__68526\ : std_logic;
signal \N__68523\ : std_logic;
signal \N__68522\ : std_logic;
signal \N__68521\ : std_logic;
signal \N__68518\ : std_logic;
signal \N__68515\ : std_logic;
signal \N__68512\ : std_logic;
signal \N__68509\ : std_logic;
signal \N__68506\ : std_logic;
signal \N__68503\ : std_logic;
signal \N__68500\ : std_logic;
signal \N__68495\ : std_logic;
signal \N__68492\ : std_logic;
signal \N__68489\ : std_logic;
signal \N__68484\ : std_logic;
signal \N__68481\ : std_logic;
signal \N__68476\ : std_logic;
signal \N__68473\ : std_logic;
signal \N__68470\ : std_logic;
signal \N__68463\ : std_logic;
signal \N__68456\ : std_logic;
signal \N__68447\ : std_logic;
signal \N__68434\ : std_logic;
signal \N__68431\ : std_logic;
signal \N__68430\ : std_logic;
signal \N__68429\ : std_logic;
signal \N__68428\ : std_logic;
signal \N__68425\ : std_logic;
signal \N__68422\ : std_logic;
signal \N__68419\ : std_logic;
signal \N__68416\ : std_logic;
signal \N__68413\ : std_logic;
signal \N__68410\ : std_logic;
signal \N__68405\ : std_logic;
signal \N__68398\ : std_logic;
signal \N__68395\ : std_logic;
signal \N__68392\ : std_logic;
signal \N__68391\ : std_logic;
signal \N__68388\ : std_logic;
signal \N__68385\ : std_logic;
signal \N__68384\ : std_logic;
signal \N__68383\ : std_logic;
signal \N__68378\ : std_logic;
signal \N__68375\ : std_logic;
signal \N__68374\ : std_logic;
signal \N__68371\ : std_logic;
signal \N__68368\ : std_logic;
signal \N__68365\ : std_logic;
signal \N__68364\ : std_logic;
signal \N__68361\ : std_logic;
signal \N__68356\ : std_logic;
signal \N__68355\ : std_logic;
signal \N__68352\ : std_logic;
signal \N__68349\ : std_logic;
signal \N__68348\ : std_logic;
signal \N__68345\ : std_logic;
signal \N__68342\ : std_logic;
signal \N__68339\ : std_logic;
signal \N__68336\ : std_logic;
signal \N__68333\ : std_logic;
signal \N__68330\ : std_logic;
signal \N__68327\ : std_logic;
signal \N__68324\ : std_logic;
signal \N__68317\ : std_logic;
signal \N__68308\ : std_logic;
signal \N__68307\ : std_logic;
signal \N__68304\ : std_logic;
signal \N__68301\ : std_logic;
signal \N__68300\ : std_logic;
signal \N__68299\ : std_logic;
signal \N__68296\ : std_logic;
signal \N__68293\ : std_logic;
signal \N__68290\ : std_logic;
signal \N__68289\ : std_logic;
signal \N__68286\ : std_logic;
signal \N__68283\ : std_logic;
signal \N__68278\ : std_logic;
signal \N__68275\ : std_logic;
signal \N__68274\ : std_logic;
signal \N__68271\ : std_logic;
signal \N__68266\ : std_logic;
signal \N__68263\ : std_logic;
signal \N__68260\ : std_logic;
signal \N__68257\ : std_logic;
signal \N__68252\ : std_logic;
signal \N__68245\ : std_logic;
signal \N__68242\ : std_logic;
signal \N__68239\ : std_logic;
signal \N__68236\ : std_logic;
signal \N__68235\ : std_logic;
signal \N__68234\ : std_logic;
signal \N__68229\ : std_logic;
signal \N__68228\ : std_logic;
signal \N__68227\ : std_logic;
signal \N__68224\ : std_logic;
signal \N__68221\ : std_logic;
signal \N__68218\ : std_logic;
signal \N__68217\ : std_logic;
signal \N__68214\ : std_logic;
signal \N__68213\ : std_logic;
signal \N__68208\ : std_logic;
signal \N__68203\ : std_logic;
signal \N__68200\ : std_logic;
signal \N__68197\ : std_logic;
signal \N__68196\ : std_logic;
signal \N__68195\ : std_logic;
signal \N__68192\ : std_logic;
signal \N__68185\ : std_logic;
signal \N__68180\ : std_logic;
signal \N__68173\ : std_logic;
signal \N__68170\ : std_logic;
signal \N__68169\ : std_logic;
signal \N__68166\ : std_logic;
signal \N__68165\ : std_logic;
signal \N__68162\ : std_logic;
signal \N__68159\ : std_logic;
signal \N__68158\ : std_logic;
signal \N__68157\ : std_logic;
signal \N__68154\ : std_logic;
signal \N__68151\ : std_logic;
signal \N__68148\ : std_logic;
signal \N__68143\ : std_logic;
signal \N__68140\ : std_logic;
signal \N__68133\ : std_logic;
signal \N__68130\ : std_logic;
signal \N__68125\ : std_logic;
signal \N__68124\ : std_logic;
signal \N__68121\ : std_logic;
signal \N__68120\ : std_logic;
signal \N__68119\ : std_logic;
signal \N__68114\ : std_logic;
signal \N__68113\ : std_logic;
signal \N__68112\ : std_logic;
signal \N__68109\ : std_logic;
signal \N__68106\ : std_logic;
signal \N__68105\ : std_logic;
signal \N__68104\ : std_logic;
signal \N__68101\ : std_logic;
signal \N__68096\ : std_logic;
signal \N__68093\ : std_logic;
signal \N__68090\ : std_logic;
signal \N__68085\ : std_logic;
signal \N__68084\ : std_logic;
signal \N__68081\ : std_logic;
signal \N__68076\ : std_logic;
signal \N__68071\ : std_logic;
signal \N__68070\ : std_logic;
signal \N__68067\ : std_logic;
signal \N__68064\ : std_logic;
signal \N__68059\ : std_logic;
signal \N__68056\ : std_logic;
signal \N__68047\ : std_logic;
signal \N__68044\ : std_logic;
signal \N__68043\ : std_logic;
signal \N__68040\ : std_logic;
signal \N__68037\ : std_logic;
signal \N__68034\ : std_logic;
signal \N__68031\ : std_logic;
signal \N__68026\ : std_logic;
signal \N__68023\ : std_logic;
signal \N__68022\ : std_logic;
signal \N__68019\ : std_logic;
signal \N__68018\ : std_logic;
signal \N__68017\ : std_logic;
signal \N__68014\ : std_logic;
signal \N__68011\ : std_logic;
signal \N__68008\ : std_logic;
signal \N__68005\ : std_logic;
signal \N__68002\ : std_logic;
signal \N__67993\ : std_logic;
signal \N__67990\ : std_logic;
signal \N__67987\ : std_logic;
signal \N__67984\ : std_logic;
signal \N__67983\ : std_logic;
signal \N__67982\ : std_logic;
signal \N__67981\ : std_logic;
signal \N__67980\ : std_logic;
signal \N__67979\ : std_logic;
signal \N__67976\ : std_logic;
signal \N__67973\ : std_logic;
signal \N__67972\ : std_logic;
signal \N__67971\ : std_logic;
signal \N__67968\ : std_logic;
signal \N__67965\ : std_logic;
signal \N__67964\ : std_logic;
signal \N__67961\ : std_logic;
signal \N__67958\ : std_logic;
signal \N__67953\ : std_logic;
signal \N__67952\ : std_logic;
signal \N__67951\ : std_logic;
signal \N__67950\ : std_logic;
signal \N__67949\ : std_logic;
signal \N__67948\ : std_logic;
signal \N__67947\ : std_logic;
signal \N__67946\ : std_logic;
signal \N__67945\ : std_logic;
signal \N__67944\ : std_logic;
signal \N__67941\ : std_logic;
signal \N__67940\ : std_logic;
signal \N__67939\ : std_logic;
signal \N__67936\ : std_logic;
signal \N__67933\ : std_logic;
signal \N__67932\ : std_logic;
signal \N__67929\ : std_logic;
signal \N__67926\ : std_logic;
signal \N__67923\ : std_logic;
signal \N__67922\ : std_logic;
signal \N__67921\ : std_logic;
signal \N__67920\ : std_logic;
signal \N__67919\ : std_logic;
signal \N__67916\ : std_logic;
signal \N__67913\ : std_logic;
signal \N__67912\ : std_logic;
signal \N__67911\ : std_logic;
signal \N__67908\ : std_logic;
signal \N__67905\ : std_logic;
signal \N__67900\ : std_logic;
signal \N__67897\ : std_logic;
signal \N__67890\ : std_logic;
signal \N__67889\ : std_logic;
signal \N__67886\ : std_logic;
signal \N__67883\ : std_logic;
signal \N__67880\ : std_logic;
signal \N__67877\ : std_logic;
signal \N__67872\ : std_logic;
signal \N__67869\ : std_logic;
signal \N__67866\ : std_logic;
signal \N__67861\ : std_logic;
signal \N__67858\ : std_logic;
signal \N__67855\ : std_logic;
signal \N__67854\ : std_logic;
signal \N__67849\ : std_logic;
signal \N__67846\ : std_logic;
signal \N__67843\ : std_logic;
signal \N__67840\ : std_logic;
signal \N__67837\ : std_logic;
signal \N__67826\ : std_logic;
signal \N__67821\ : std_logic;
signal \N__67818\ : std_logic;
signal \N__67813\ : std_logic;
signal \N__67808\ : std_logic;
signal \N__67803\ : std_logic;
signal \N__67802\ : std_logic;
signal \N__67799\ : std_logic;
signal \N__67796\ : std_logic;
signal \N__67793\ : std_logic;
signal \N__67790\ : std_logic;
signal \N__67785\ : std_logic;
signal \N__67778\ : std_logic;
signal \N__67777\ : std_logic;
signal \N__67776\ : std_logic;
signal \N__67773\ : std_logic;
signal \N__67770\ : std_logic;
signal \N__67763\ : std_logic;
signal \N__67760\ : std_logic;
signal \N__67757\ : std_logic;
signal \N__67750\ : std_logic;
signal \N__67747\ : std_logic;
signal \N__67744\ : std_logic;
signal \N__67741\ : std_logic;
signal \N__67738\ : std_logic;
signal \N__67733\ : std_logic;
signal \N__67730\ : std_logic;
signal \N__67723\ : std_logic;
signal \N__67718\ : std_logic;
signal \N__67705\ : std_logic;
signal \N__67704\ : std_logic;
signal \N__67701\ : std_logic;
signal \N__67698\ : std_logic;
signal \N__67697\ : std_logic;
signal \N__67696\ : std_logic;
signal \N__67693\ : std_logic;
signal \N__67690\ : std_logic;
signal \N__67685\ : std_logic;
signal \N__67682\ : std_logic;
signal \N__67675\ : std_logic;
signal \N__67674\ : std_logic;
signal \N__67673\ : std_logic;
signal \N__67670\ : std_logic;
signal \N__67667\ : std_logic;
signal \N__67666\ : std_logic;
signal \N__67663\ : std_logic;
signal \N__67658\ : std_logic;
signal \N__67657\ : std_logic;
signal \N__67654\ : std_logic;
signal \N__67649\ : std_logic;
signal \N__67646\ : std_logic;
signal \N__67639\ : std_logic;
signal \N__67636\ : std_logic;
signal \N__67633\ : std_logic;
signal \N__67630\ : std_logic;
signal \N__67629\ : std_logic;
signal \N__67626\ : std_logic;
signal \N__67623\ : std_logic;
signal \N__67618\ : std_logic;
signal \N__67615\ : std_logic;
signal \N__67614\ : std_logic;
signal \N__67613\ : std_logic;
signal \N__67610\ : std_logic;
signal \N__67607\ : std_logic;
signal \N__67604\ : std_logic;
signal \N__67601\ : std_logic;
signal \N__67598\ : std_logic;
signal \N__67595\ : std_logic;
signal \N__67590\ : std_logic;
signal \N__67587\ : std_logic;
signal \N__67582\ : std_logic;
signal \N__67579\ : std_logic;
signal \N__67576\ : std_logic;
signal \N__67573\ : std_logic;
signal \N__67570\ : std_logic;
signal \N__67567\ : std_logic;
signal \N__67566\ : std_logic;
signal \N__67563\ : std_logic;
signal \N__67562\ : std_logic;
signal \N__67559\ : std_logic;
signal \N__67556\ : std_logic;
signal \N__67553\ : std_logic;
signal \N__67550\ : std_logic;
signal \N__67547\ : std_logic;
signal \N__67544\ : std_logic;
signal \N__67541\ : std_logic;
signal \N__67538\ : std_logic;
signal \N__67531\ : std_logic;
signal \N__67530\ : std_logic;
signal \N__67529\ : std_logic;
signal \N__67528\ : std_logic;
signal \N__67527\ : std_logic;
signal \N__67526\ : std_logic;
signal \N__67523\ : std_logic;
signal \N__67522\ : std_logic;
signal \N__67519\ : std_logic;
signal \N__67516\ : std_logic;
signal \N__67511\ : std_logic;
signal \N__67508\ : std_logic;
signal \N__67505\ : std_logic;
signal \N__67504\ : std_logic;
signal \N__67501\ : std_logic;
signal \N__67498\ : std_logic;
signal \N__67495\ : std_logic;
signal \N__67492\ : std_logic;
signal \N__67489\ : std_logic;
signal \N__67486\ : std_logic;
signal \N__67483\ : std_logic;
signal \N__67478\ : std_logic;
signal \N__67475\ : std_logic;
signal \N__67472\ : std_logic;
signal \N__67467\ : std_logic;
signal \N__67462\ : std_logic;
signal \N__67459\ : std_logic;
signal \N__67456\ : std_logic;
signal \N__67453\ : std_logic;
signal \N__67450\ : std_logic;
signal \N__67447\ : std_logic;
signal \N__67438\ : std_logic;
signal \N__67435\ : std_logic;
signal \N__67434\ : std_logic;
signal \N__67431\ : std_logic;
signal \N__67428\ : std_logic;
signal \N__67427\ : std_logic;
signal \N__67424\ : std_logic;
signal \N__67421\ : std_logic;
signal \N__67418\ : std_logic;
signal \N__67413\ : std_logic;
signal \N__67408\ : std_logic;
signal \N__67405\ : std_logic;
signal \N__67404\ : std_logic;
signal \N__67401\ : std_logic;
signal \N__67398\ : std_logic;
signal \N__67393\ : std_logic;
signal \N__67390\ : std_logic;
signal \N__67387\ : std_logic;
signal \N__67386\ : std_logic;
signal \N__67383\ : std_logic;
signal \N__67380\ : std_logic;
signal \N__67379\ : std_logic;
signal \N__67378\ : std_logic;
signal \N__67373\ : std_logic;
signal \N__67368\ : std_logic;
signal \N__67365\ : std_logic;
signal \N__67360\ : std_logic;
signal \N__67357\ : std_logic;
signal \N__67354\ : std_logic;
signal \N__67351\ : std_logic;
signal \N__67348\ : std_logic;
signal \N__67345\ : std_logic;
signal \N__67342\ : std_logic;
signal \N__67339\ : std_logic;
signal \N__67336\ : std_logic;
signal \N__67333\ : std_logic;
signal \N__67330\ : std_logic;
signal \N__67327\ : std_logic;
signal \N__67324\ : std_logic;
signal \N__67321\ : std_logic;
signal \N__67318\ : std_logic;
signal \N__67315\ : std_logic;
signal \N__67312\ : std_logic;
signal \N__67309\ : std_logic;
signal \N__67306\ : std_logic;
signal \N__67303\ : std_logic;
signal \N__67302\ : std_logic;
signal \N__67299\ : std_logic;
signal \N__67296\ : std_logic;
signal \N__67293\ : std_logic;
signal \N__67290\ : std_logic;
signal \N__67289\ : std_logic;
signal \N__67288\ : std_logic;
signal \N__67285\ : std_logic;
signal \N__67282\ : std_logic;
signal \N__67277\ : std_logic;
signal \N__67270\ : std_logic;
signal \N__67267\ : std_logic;
signal \N__67266\ : std_logic;
signal \N__67265\ : std_logic;
signal \N__67264\ : std_logic;
signal \N__67263\ : std_logic;
signal \N__67260\ : std_logic;
signal \N__67255\ : std_logic;
signal \N__67250\ : std_logic;
signal \N__67243\ : std_logic;
signal \N__67242\ : std_logic;
signal \N__67241\ : std_logic;
signal \N__67234\ : std_logic;
signal \N__67231\ : std_logic;
signal \N__67228\ : std_logic;
signal \N__67227\ : std_logic;
signal \N__67226\ : std_logic;
signal \N__67225\ : std_logic;
signal \N__67224\ : std_logic;
signal \N__67223\ : std_logic;
signal \N__67222\ : std_logic;
signal \N__67221\ : std_logic;
signal \N__67220\ : std_logic;
signal \N__67219\ : std_logic;
signal \N__67218\ : std_logic;
signal \N__67213\ : std_logic;
signal \N__67204\ : std_logic;
signal \N__67201\ : std_logic;
signal \N__67200\ : std_logic;
signal \N__67199\ : std_logic;
signal \N__67198\ : std_logic;
signal \N__67197\ : std_logic;
signal \N__67196\ : std_logic;
signal \N__67191\ : std_logic;
signal \N__67188\ : std_logic;
signal \N__67187\ : std_logic;
signal \N__67184\ : std_logic;
signal \N__67179\ : std_logic;
signal \N__67178\ : std_logic;
signal \N__67173\ : std_logic;
signal \N__67170\ : std_logic;
signal \N__67167\ : std_logic;
signal \N__67166\ : std_logic;
signal \N__67163\ : std_logic;
signal \N__67160\ : std_logic;
signal \N__67157\ : std_logic;
signal \N__67154\ : std_logic;
signal \N__67151\ : std_logic;
signal \N__67148\ : std_logic;
signal \N__67145\ : std_logic;
signal \N__67144\ : std_logic;
signal \N__67141\ : std_logic;
signal \N__67138\ : std_logic;
signal \N__67135\ : std_logic;
signal \N__67132\ : std_logic;
signal \N__67131\ : std_logic;
signal \N__67130\ : std_logic;
signal \N__67127\ : std_logic;
signal \N__67122\ : std_logic;
signal \N__67119\ : std_logic;
signal \N__67118\ : std_logic;
signal \N__67113\ : std_logic;
signal \N__67108\ : std_logic;
signal \N__67105\ : std_logic;
signal \N__67102\ : std_logic;
signal \N__67095\ : std_logic;
signal \N__67092\ : std_logic;
signal \N__67089\ : std_logic;
signal \N__67086\ : std_logic;
signal \N__67081\ : std_logic;
signal \N__67078\ : std_logic;
signal \N__67075\ : std_logic;
signal \N__67072\ : std_logic;
signal \N__67065\ : std_logic;
signal \N__67062\ : std_logic;
signal \N__67057\ : std_logic;
signal \N__67054\ : std_logic;
signal \N__67051\ : std_logic;
signal \N__67044\ : std_logic;
signal \N__67041\ : std_logic;
signal \N__67038\ : std_logic;
signal \N__67035\ : std_logic;
signal \N__67030\ : std_logic;
signal \N__67021\ : std_logic;
signal \N__67020\ : std_logic;
signal \N__67017\ : std_logic;
signal \N__67014\ : std_logic;
signal \N__67011\ : std_logic;
signal \N__67008\ : std_logic;
signal \N__67005\ : std_logic;
signal \N__67002\ : std_logic;
signal \N__66999\ : std_logic;
signal \N__66994\ : std_logic;
signal \N__66991\ : std_logic;
signal \N__66988\ : std_logic;
signal \N__66987\ : std_logic;
signal \N__66984\ : std_logic;
signal \N__66981\ : std_logic;
signal \N__66980\ : std_logic;
signal \N__66979\ : std_logic;
signal \N__66978\ : std_logic;
signal \N__66977\ : std_logic;
signal \N__66976\ : std_logic;
signal \N__66975\ : std_logic;
signal \N__66974\ : std_logic;
signal \N__66973\ : std_logic;
signal \N__66972\ : std_logic;
signal \N__66963\ : std_logic;
signal \N__66962\ : std_logic;
signal \N__66959\ : std_logic;
signal \N__66958\ : std_logic;
signal \N__66957\ : std_logic;
signal \N__66956\ : std_logic;
signal \N__66955\ : std_logic;
signal \N__66954\ : std_logic;
signal \N__66953\ : std_logic;
signal \N__66952\ : std_logic;
signal \N__66949\ : std_logic;
signal \N__66948\ : std_logic;
signal \N__66947\ : std_logic;
signal \N__66944\ : std_logic;
signal \N__66943\ : std_logic;
signal \N__66942\ : std_logic;
signal \N__66941\ : std_logic;
signal \N__66938\ : std_logic;
signal \N__66935\ : std_logic;
signal \N__66934\ : std_logic;
signal \N__66933\ : std_logic;
signal \N__66928\ : std_logic;
signal \N__66925\ : std_logic;
signal \N__66924\ : std_logic;
signal \N__66923\ : std_logic;
signal \N__66918\ : std_logic;
signal \N__66917\ : std_logic;
signal \N__66916\ : std_logic;
signal \N__66913\ : std_logic;
signal \N__66912\ : std_logic;
signal \N__66909\ : std_logic;
signal \N__66900\ : std_logic;
signal \N__66899\ : std_logic;
signal \N__66898\ : std_logic;
signal \N__66897\ : std_logic;
signal \N__66896\ : std_logic;
signal \N__66889\ : std_logic;
signal \N__66882\ : std_logic;
signal \N__66881\ : std_logic;
signal \N__66880\ : std_logic;
signal \N__66879\ : std_logic;
signal \N__66868\ : std_logic;
signal \N__66865\ : std_logic;
signal \N__66860\ : std_logic;
signal \N__66857\ : std_logic;
signal \N__66854\ : std_logic;
signal \N__66851\ : std_logic;
signal \N__66850\ : std_logic;
signal \N__66849\ : std_logic;
signal \N__66846\ : std_logic;
signal \N__66841\ : std_logic;
signal \N__66838\ : std_logic;
signal \N__66835\ : std_logic;
signal \N__66832\ : std_logic;
signal \N__66829\ : std_logic;
signal \N__66826\ : std_logic;
signal \N__66821\ : std_logic;
signal \N__66816\ : std_logic;
signal \N__66809\ : std_logic;
signal \N__66806\ : std_logic;
signal \N__66799\ : std_logic;
signal \N__66794\ : std_logic;
signal \N__66791\ : std_logic;
signal \N__66788\ : std_logic;
signal \N__66785\ : std_logic;
signal \N__66782\ : std_logic;
signal \N__66777\ : std_logic;
signal \N__66774\ : std_logic;
signal \N__66771\ : std_logic;
signal \N__66768\ : std_logic;
signal \N__66761\ : std_logic;
signal \N__66758\ : std_logic;
signal \N__66755\ : std_logic;
signal \N__66754\ : std_logic;
signal \N__66751\ : std_logic;
signal \N__66748\ : std_logic;
signal \N__66739\ : std_logic;
signal \N__66732\ : std_logic;
signal \N__66729\ : std_logic;
signal \N__66724\ : std_logic;
signal \N__66721\ : std_logic;
signal \N__66718\ : std_logic;
signal \N__66711\ : std_logic;
signal \N__66708\ : std_logic;
signal \N__66705\ : std_logic;
signal \N__66694\ : std_logic;
signal \N__66691\ : std_logic;
signal \N__66690\ : std_logic;
signal \N__66687\ : std_logic;
signal \N__66684\ : std_logic;
signal \N__66681\ : std_logic;
signal \N__66676\ : std_logic;
signal \N__66673\ : std_logic;
signal \N__66670\ : std_logic;
signal \N__66667\ : std_logic;
signal \N__66664\ : std_logic;
signal \N__66661\ : std_logic;
signal \N__66658\ : std_logic;
signal \N__66655\ : std_logic;
signal \N__66652\ : std_logic;
signal \N__66649\ : std_logic;
signal \N__66648\ : std_logic;
signal \N__66647\ : std_logic;
signal \N__66644\ : std_logic;
signal \N__66641\ : std_logic;
signal \N__66636\ : std_logic;
signal \N__66633\ : std_logic;
signal \N__66632\ : std_logic;
signal \N__66631\ : std_logic;
signal \N__66628\ : std_logic;
signal \N__66625\ : std_logic;
signal \N__66622\ : std_logic;
signal \N__66619\ : std_logic;
signal \N__66616\ : std_logic;
signal \N__66613\ : std_logic;
signal \N__66604\ : std_logic;
signal \N__66601\ : std_logic;
signal \N__66598\ : std_logic;
signal \N__66595\ : std_logic;
signal \N__66592\ : std_logic;
signal \N__66589\ : std_logic;
signal \N__66586\ : std_logic;
signal \N__66583\ : std_logic;
signal \N__66582\ : std_logic;
signal \N__66579\ : std_logic;
signal \N__66576\ : std_logic;
signal \N__66571\ : std_logic;
signal \N__66570\ : std_logic;
signal \N__66567\ : std_logic;
signal \N__66564\ : std_logic;
signal \N__66559\ : std_logic;
signal \N__66556\ : std_logic;
signal \N__66553\ : std_logic;
signal \N__66550\ : std_logic;
signal \N__66547\ : std_logic;
signal \N__66546\ : std_logic;
signal \N__66545\ : std_logic;
signal \N__66542\ : std_logic;
signal \N__66537\ : std_logic;
signal \N__66532\ : std_logic;
signal \N__66529\ : std_logic;
signal \N__66526\ : std_logic;
signal \N__66523\ : std_logic;
signal \N__66520\ : std_logic;
signal \N__66517\ : std_logic;
signal \N__66514\ : std_logic;
signal \N__66511\ : std_logic;
signal \N__66510\ : std_logic;
signal \N__66507\ : std_logic;
signal \N__66504\ : std_logic;
signal \N__66501\ : std_logic;
signal \N__66500\ : std_logic;
signal \N__66497\ : std_logic;
signal \N__66496\ : std_logic;
signal \N__66493\ : std_logic;
signal \N__66490\ : std_logic;
signal \N__66487\ : std_logic;
signal \N__66484\ : std_logic;
signal \N__66481\ : std_logic;
signal \N__66476\ : std_logic;
signal \N__66469\ : std_logic;
signal \N__66466\ : std_logic;
signal \N__66465\ : std_logic;
signal \N__66464\ : std_logic;
signal \N__66461\ : std_logic;
signal \N__66458\ : std_logic;
signal \N__66455\ : std_logic;
signal \N__66454\ : std_logic;
signal \N__66453\ : std_logic;
signal \N__66448\ : std_logic;
signal \N__66445\ : std_logic;
signal \N__66440\ : std_logic;
signal \N__66437\ : std_logic;
signal \N__66434\ : std_logic;
signal \N__66427\ : std_logic;
signal \N__66424\ : std_logic;
signal \N__66421\ : std_logic;
signal \N__66418\ : std_logic;
signal \N__66417\ : std_logic;
signal \N__66416\ : std_logic;
signal \N__66411\ : std_logic;
signal \N__66408\ : std_logic;
signal \N__66405\ : std_logic;
signal \N__66402\ : std_logic;
signal \N__66397\ : std_logic;
signal \N__66396\ : std_logic;
signal \N__66395\ : std_logic;
signal \N__66392\ : std_logic;
signal \N__66387\ : std_logic;
signal \N__66382\ : std_logic;
signal \N__66381\ : std_logic;
signal \N__66378\ : std_logic;
signal \N__66375\ : std_logic;
signal \N__66370\ : std_logic;
signal \N__66367\ : std_logic;
signal \N__66364\ : std_logic;
signal \N__66361\ : std_logic;
signal \N__66358\ : std_logic;
signal \N__66355\ : std_logic;
signal \N__66354\ : std_logic;
signal \N__66351\ : std_logic;
signal \N__66348\ : std_logic;
signal \N__66345\ : std_logic;
signal \N__66342\ : std_logic;
signal \N__66337\ : std_logic;
signal \N__66336\ : std_logic;
signal \N__66333\ : std_logic;
signal \N__66330\ : std_logic;
signal \N__66327\ : std_logic;
signal \N__66326\ : std_logic;
signal \N__66323\ : std_logic;
signal \N__66320\ : std_logic;
signal \N__66317\ : std_logic;
signal \N__66310\ : std_logic;
signal \N__66307\ : std_logic;
signal \N__66304\ : std_logic;
signal \N__66301\ : std_logic;
signal \N__66298\ : std_logic;
signal \N__66295\ : std_logic;
signal \N__66294\ : std_logic;
signal \N__66291\ : std_logic;
signal \N__66288\ : std_logic;
signal \N__66287\ : std_logic;
signal \N__66286\ : std_logic;
signal \N__66281\ : std_logic;
signal \N__66278\ : std_logic;
signal \N__66275\ : std_logic;
signal \N__66272\ : std_logic;
signal \N__66269\ : std_logic;
signal \N__66266\ : std_logic;
signal \N__66261\ : std_logic;
signal \N__66256\ : std_logic;
signal \N__66253\ : std_logic;
signal \N__66250\ : std_logic;
signal \N__66247\ : std_logic;
signal \N__66244\ : std_logic;
signal \N__66243\ : std_logic;
signal \N__66240\ : std_logic;
signal \N__66239\ : std_logic;
signal \N__66236\ : std_logic;
signal \N__66233\ : std_logic;
signal \N__66230\ : std_logic;
signal \N__66227\ : std_logic;
signal \N__66224\ : std_logic;
signal \N__66221\ : std_logic;
signal \N__66216\ : std_logic;
signal \N__66211\ : std_logic;
signal \N__66210\ : std_logic;
signal \N__66209\ : std_logic;
signal \N__66206\ : std_logic;
signal \N__66205\ : std_logic;
signal \N__66204\ : std_logic;
signal \N__66203\ : std_logic;
signal \N__66198\ : std_logic;
signal \N__66195\ : std_logic;
signal \N__66194\ : std_logic;
signal \N__66193\ : std_logic;
signal \N__66190\ : std_logic;
signal \N__66189\ : std_logic;
signal \N__66188\ : std_logic;
signal \N__66187\ : std_logic;
signal \N__66186\ : std_logic;
signal \N__66185\ : std_logic;
signal \N__66184\ : std_logic;
signal \N__66181\ : std_logic;
signal \N__66178\ : std_logic;
signal \N__66177\ : std_logic;
signal \N__66172\ : std_logic;
signal \N__66169\ : std_logic;
signal \N__66166\ : std_logic;
signal \N__66163\ : std_logic;
signal \N__66162\ : std_logic;
signal \N__66159\ : std_logic;
signal \N__66158\ : std_logic;
signal \N__66157\ : std_logic;
signal \N__66156\ : std_logic;
signal \N__66155\ : std_logic;
signal \N__66154\ : std_logic;
signal \N__66153\ : std_logic;
signal \N__66150\ : std_logic;
signal \N__66147\ : std_logic;
signal \N__66146\ : std_logic;
signal \N__66145\ : std_logic;
signal \N__66144\ : std_logic;
signal \N__66141\ : std_logic;
signal \N__66140\ : std_logic;
signal \N__66139\ : std_logic;
signal \N__66136\ : std_logic;
signal \N__66133\ : std_logic;
signal \N__66126\ : std_logic;
signal \N__66125\ : std_logic;
signal \N__66122\ : std_logic;
signal \N__66121\ : std_logic;
signal \N__66120\ : std_logic;
signal \N__66117\ : std_logic;
signal \N__66114\ : std_logic;
signal \N__66111\ : std_logic;
signal \N__66102\ : std_logic;
signal \N__66099\ : std_logic;
signal \N__66096\ : std_logic;
signal \N__66093\ : std_logic;
signal \N__66084\ : std_logic;
signal \N__66081\ : std_logic;
signal \N__66078\ : std_logic;
signal \N__66071\ : std_logic;
signal \N__66068\ : std_logic;
signal \N__66067\ : std_logic;
signal \N__66066\ : std_logic;
signal \N__66061\ : std_logic;
signal \N__66060\ : std_logic;
signal \N__66057\ : std_logic;
signal \N__66054\ : std_logic;
signal \N__66051\ : std_logic;
signal \N__66050\ : std_logic;
signal \N__66047\ : std_logic;
signal \N__66046\ : std_logic;
signal \N__66045\ : std_logic;
signal \N__66040\ : std_logic;
signal \N__66039\ : std_logic;
signal \N__66038\ : std_logic;
signal \N__66033\ : std_logic;
signal \N__66026\ : std_logic;
signal \N__66023\ : std_logic;
signal \N__66020\ : std_logic;
signal \N__66013\ : std_logic;
signal \N__66012\ : std_logic;
signal \N__66011\ : std_logic;
signal \N__66008\ : std_logic;
signal \N__66007\ : std_logic;
signal \N__66004\ : std_logic;
signal \N__66001\ : std_logic;
signal \N__65998\ : std_logic;
signal \N__65995\ : std_logic;
signal \N__65992\ : std_logic;
signal \N__65989\ : std_logic;
signal \N__65986\ : std_logic;
signal \N__65979\ : std_logic;
signal \N__65976\ : std_logic;
signal \N__65971\ : std_logic;
signal \N__65968\ : std_logic;
signal \N__65965\ : std_logic;
signal \N__65958\ : std_logic;
signal \N__65955\ : std_logic;
signal \N__65952\ : std_logic;
signal \N__65949\ : std_logic;
signal \N__65944\ : std_logic;
signal \N__65941\ : std_logic;
signal \N__65936\ : std_logic;
signal \N__65933\ : std_logic;
signal \N__65930\ : std_logic;
signal \N__65921\ : std_logic;
signal \N__65918\ : std_logic;
signal \N__65913\ : std_logic;
signal \N__65904\ : std_logic;
signal \N__65901\ : std_logic;
signal \N__65894\ : std_logic;
signal \N__65891\ : std_logic;
signal \N__65888\ : std_logic;
signal \N__65885\ : std_logic;
signal \N__65878\ : std_logic;
signal \N__65869\ : std_logic;
signal \N__65868\ : std_logic;
signal \N__65865\ : std_logic;
signal \N__65864\ : std_logic;
signal \N__65863\ : std_logic;
signal \N__65860\ : std_logic;
signal \N__65857\ : std_logic;
signal \N__65854\ : std_logic;
signal \N__65853\ : std_logic;
signal \N__65850\ : std_logic;
signal \N__65849\ : std_logic;
signal \N__65846\ : std_logic;
signal \N__65843\ : std_logic;
signal \N__65840\ : std_logic;
signal \N__65837\ : std_logic;
signal \N__65834\ : std_logic;
signal \N__65831\ : std_logic;
signal \N__65828\ : std_logic;
signal \N__65823\ : std_logic;
signal \N__65818\ : std_logic;
signal \N__65815\ : std_logic;
signal \N__65812\ : std_logic;
signal \N__65809\ : std_logic;
signal \N__65806\ : std_logic;
signal \N__65797\ : std_logic;
signal \N__65796\ : std_logic;
signal \N__65795\ : std_logic;
signal \N__65792\ : std_logic;
signal \N__65789\ : std_logic;
signal \N__65786\ : std_logic;
signal \N__65783\ : std_logic;
signal \N__65782\ : std_logic;
signal \N__65781\ : std_logic;
signal \N__65780\ : std_logic;
signal \N__65775\ : std_logic;
signal \N__65772\ : std_logic;
signal \N__65769\ : std_logic;
signal \N__65766\ : std_logic;
signal \N__65763\ : std_logic;
signal \N__65762\ : std_logic;
signal \N__65759\ : std_logic;
signal \N__65752\ : std_logic;
signal \N__65749\ : std_logic;
signal \N__65746\ : std_logic;
signal \N__65743\ : std_logic;
signal \N__65738\ : std_logic;
signal \N__65735\ : std_logic;
signal \N__65732\ : std_logic;
signal \N__65729\ : std_logic;
signal \N__65722\ : std_logic;
signal \N__65719\ : std_logic;
signal \N__65716\ : std_logic;
signal \N__65715\ : std_logic;
signal \N__65712\ : std_logic;
signal \N__65711\ : std_logic;
signal \N__65708\ : std_logic;
signal \N__65705\ : std_logic;
signal \N__65702\ : std_logic;
signal \N__65695\ : std_logic;
signal \N__65694\ : std_logic;
signal \N__65693\ : std_logic;
signal \N__65690\ : std_logic;
signal \N__65687\ : std_logic;
signal \N__65684\ : std_logic;
signal \N__65681\ : std_logic;
signal \N__65680\ : std_logic;
signal \N__65675\ : std_logic;
signal \N__65674\ : std_logic;
signal \N__65671\ : std_logic;
signal \N__65668\ : std_logic;
signal \N__65665\ : std_logic;
signal \N__65662\ : std_logic;
signal \N__65661\ : std_logic;
signal \N__65658\ : std_logic;
signal \N__65655\ : std_logic;
signal \N__65652\ : std_logic;
signal \N__65649\ : std_logic;
signal \N__65646\ : std_logic;
signal \N__65643\ : std_logic;
signal \N__65638\ : std_logic;
signal \N__65635\ : std_logic;
signal \N__65626\ : std_logic;
signal \N__65623\ : std_logic;
signal \N__65620\ : std_logic;
signal \N__65619\ : std_logic;
signal \N__65618\ : std_logic;
signal \N__65615\ : std_logic;
signal \N__65610\ : std_logic;
signal \N__65605\ : std_logic;
signal \N__65602\ : std_logic;
signal \N__65599\ : std_logic;
signal \N__65598\ : std_logic;
signal \N__65597\ : std_logic;
signal \N__65596\ : std_logic;
signal \N__65595\ : std_logic;
signal \N__65594\ : std_logic;
signal \N__65591\ : std_logic;
signal \N__65590\ : std_logic;
signal \N__65587\ : std_logic;
signal \N__65584\ : std_logic;
signal \N__65581\ : std_logic;
signal \N__65580\ : std_logic;
signal \N__65575\ : std_logic;
signal \N__65572\ : std_logic;
signal \N__65569\ : std_logic;
signal \N__65566\ : std_logic;
signal \N__65563\ : std_logic;
signal \N__65560\ : std_logic;
signal \N__65557\ : std_logic;
signal \N__65554\ : std_logic;
signal \N__65551\ : std_logic;
signal \N__65544\ : std_logic;
signal \N__65541\ : std_logic;
signal \N__65532\ : std_logic;
signal \N__65527\ : std_logic;
signal \N__65526\ : std_logic;
signal \N__65525\ : std_logic;
signal \N__65522\ : std_logic;
signal \N__65521\ : std_logic;
signal \N__65520\ : std_logic;
signal \N__65519\ : std_logic;
signal \N__65516\ : std_logic;
signal \N__65515\ : std_logic;
signal \N__65512\ : std_logic;
signal \N__65509\ : std_logic;
signal \N__65504\ : std_logic;
signal \N__65499\ : std_logic;
signal \N__65496\ : std_logic;
signal \N__65495\ : std_logic;
signal \N__65494\ : std_logic;
signal \N__65493\ : std_logic;
signal \N__65490\ : std_logic;
signal \N__65485\ : std_logic;
signal \N__65482\ : std_logic;
signal \N__65479\ : std_logic;
signal \N__65474\ : std_logic;
signal \N__65471\ : std_logic;
signal \N__65466\ : std_logic;
signal \N__65459\ : std_logic;
signal \N__65452\ : std_logic;
signal \N__65449\ : std_logic;
signal \N__65448\ : std_logic;
signal \N__65445\ : std_logic;
signal \N__65442\ : std_logic;
signal \N__65439\ : std_logic;
signal \N__65434\ : std_logic;
signal \N__65433\ : std_logic;
signal \N__65430\ : std_logic;
signal \N__65429\ : std_logic;
signal \N__65426\ : std_logic;
signal \N__65423\ : std_logic;
signal \N__65420\ : std_logic;
signal \N__65417\ : std_logic;
signal \N__65412\ : std_logic;
signal \N__65407\ : std_logic;
signal \N__65406\ : std_logic;
signal \N__65403\ : std_logic;
signal \N__65400\ : std_logic;
signal \N__65399\ : std_logic;
signal \N__65398\ : std_logic;
signal \N__65397\ : std_logic;
signal \N__65394\ : std_logic;
signal \N__65391\ : std_logic;
signal \N__65388\ : std_logic;
signal \N__65385\ : std_logic;
signal \N__65382\ : std_logic;
signal \N__65379\ : std_logic;
signal \N__65374\ : std_logic;
signal \N__65371\ : std_logic;
signal \N__65368\ : std_logic;
signal \N__65365\ : std_logic;
signal \N__65362\ : std_logic;
signal \N__65359\ : std_logic;
signal \N__65350\ : std_logic;
signal \N__65347\ : std_logic;
signal \N__65344\ : std_logic;
signal \N__65343\ : std_logic;
signal \N__65340\ : std_logic;
signal \N__65337\ : std_logic;
signal \N__65334\ : std_logic;
signal \N__65331\ : std_logic;
signal \N__65326\ : std_logic;
signal \N__65325\ : std_logic;
signal \N__65322\ : std_logic;
signal \N__65321\ : std_logic;
signal \N__65320\ : std_logic;
signal \N__65317\ : std_logic;
signal \N__65314\ : std_logic;
signal \N__65309\ : std_logic;
signal \N__65306\ : std_logic;
signal \N__65299\ : std_logic;
signal \N__65298\ : std_logic;
signal \N__65293\ : std_logic;
signal \N__65292\ : std_logic;
signal \N__65289\ : std_logic;
signal \N__65286\ : std_logic;
signal \N__65281\ : std_logic;
signal \N__65278\ : std_logic;
signal \N__65275\ : std_logic;
signal \N__65272\ : std_logic;
signal \N__65269\ : std_logic;
signal \N__65266\ : std_logic;
signal \N__65263\ : std_logic;
signal \N__65262\ : std_logic;
signal \N__65261\ : std_logic;
signal \N__65260\ : std_logic;
signal \N__65259\ : std_logic;
signal \N__65258\ : std_logic;
signal \N__65253\ : std_logic;
signal \N__65250\ : std_logic;
signal \N__65249\ : std_logic;
signal \N__65248\ : std_logic;
signal \N__65247\ : std_logic;
signal \N__65246\ : std_logic;
signal \N__65243\ : std_logic;
signal \N__65242\ : std_logic;
signal \N__65241\ : std_logic;
signal \N__65240\ : std_logic;
signal \N__65239\ : std_logic;
signal \N__65238\ : std_logic;
signal \N__65235\ : std_logic;
signal \N__65234\ : std_logic;
signal \N__65231\ : std_logic;
signal \N__65230\ : std_logic;
signal \N__65227\ : std_logic;
signal \N__65226\ : std_logic;
signal \N__65223\ : std_logic;
signal \N__65218\ : std_logic;
signal \N__65217\ : std_logic;
signal \N__65212\ : std_logic;
signal \N__65209\ : std_logic;
signal \N__65206\ : std_logic;
signal \N__65203\ : std_logic;
signal \N__65202\ : std_logic;
signal \N__65199\ : std_logic;
signal \N__65198\ : std_logic;
signal \N__65195\ : std_logic;
signal \N__65192\ : std_logic;
signal \N__65191\ : std_logic;
signal \N__65190\ : std_logic;
signal \N__65189\ : std_logic;
signal \N__65186\ : std_logic;
signal \N__65179\ : std_logic;
signal \N__65176\ : std_logic;
signal \N__65173\ : std_logic;
signal \N__65172\ : std_logic;
signal \N__65169\ : std_logic;
signal \N__65166\ : std_logic;
signal \N__65163\ : std_logic;
signal \N__65160\ : std_logic;
signal \N__65155\ : std_logic;
signal \N__65152\ : std_logic;
signal \N__65149\ : std_logic;
signal \N__65148\ : std_logic;
signal \N__65147\ : std_logic;
signal \N__65144\ : std_logic;
signal \N__65141\ : std_logic;
signal \N__65136\ : std_logic;
signal \N__65129\ : std_logic;
signal \N__65124\ : std_logic;
signal \N__65119\ : std_logic;
signal \N__65118\ : std_logic;
signal \N__65117\ : std_logic;
signal \N__65114\ : std_logic;
signal \N__65109\ : std_logic;
signal \N__65104\ : std_logic;
signal \N__65101\ : std_logic;
signal \N__65098\ : std_logic;
signal \N__65095\ : std_logic;
signal \N__65094\ : std_logic;
signal \N__65091\ : std_logic;
signal \N__65088\ : std_logic;
signal \N__65085\ : std_logic;
signal \N__65082\ : std_logic;
signal \N__65079\ : std_logic;
signal \N__65074\ : std_logic;
signal \N__65071\ : std_logic;
signal \N__65070\ : std_logic;
signal \N__65069\ : std_logic;
signal \N__65064\ : std_logic;
signal \N__65057\ : std_logic;
signal \N__65052\ : std_logic;
signal \N__65049\ : std_logic;
signal \N__65046\ : std_logic;
signal \N__65037\ : std_logic;
signal \N__65034\ : std_logic;
signal \N__65031\ : std_logic;
signal \N__65028\ : std_logic;
signal \N__65025\ : std_logic;
signal \N__65022\ : std_logic;
signal \N__65019\ : std_logic;
signal \N__65014\ : std_logic;
signal \N__65011\ : std_logic;
signal \N__65000\ : std_logic;
signal \N__64991\ : std_logic;
signal \N__64984\ : std_logic;
signal \N__64983\ : std_logic;
signal \N__64980\ : std_logic;
signal \N__64979\ : std_logic;
signal \N__64976\ : std_logic;
signal \N__64973\ : std_logic;
signal \N__64972\ : std_logic;
signal \N__64969\ : std_logic;
signal \N__64966\ : std_logic;
signal \N__64963\ : std_logic;
signal \N__64960\ : std_logic;
signal \N__64951\ : std_logic;
signal \N__64950\ : std_logic;
signal \N__64949\ : std_logic;
signal \N__64946\ : std_logic;
signal \N__64943\ : std_logic;
signal \N__64942\ : std_logic;
signal \N__64939\ : std_logic;
signal \N__64936\ : std_logic;
signal \N__64933\ : std_logic;
signal \N__64930\ : std_logic;
signal \N__64927\ : std_logic;
signal \N__64924\ : std_logic;
signal \N__64921\ : std_logic;
signal \N__64920\ : std_logic;
signal \N__64917\ : std_logic;
signal \N__64910\ : std_logic;
signal \N__64907\ : std_logic;
signal \N__64900\ : std_logic;
signal \N__64899\ : std_logic;
signal \N__64896\ : std_logic;
signal \N__64893\ : std_logic;
signal \N__64892\ : std_logic;
signal \N__64889\ : std_logic;
signal \N__64888\ : std_logic;
signal \N__64887\ : std_logic;
signal \N__64886\ : std_logic;
signal \N__64883\ : std_logic;
signal \N__64880\ : std_logic;
signal \N__64877\ : std_logic;
signal \N__64874\ : std_logic;
signal \N__64871\ : std_logic;
signal \N__64868\ : std_logic;
signal \N__64865\ : std_logic;
signal \N__64860\ : std_logic;
signal \N__64857\ : std_logic;
signal \N__64854\ : std_logic;
signal \N__64849\ : std_logic;
signal \N__64846\ : std_logic;
signal \N__64843\ : std_logic;
signal \N__64834\ : std_logic;
signal \N__64833\ : std_logic;
signal \N__64832\ : std_logic;
signal \N__64831\ : std_logic;
signal \N__64830\ : std_logic;
signal \N__64827\ : std_logic;
signal \N__64822\ : std_logic;
signal \N__64821\ : std_logic;
signal \N__64818\ : std_logic;
signal \N__64815\ : std_logic;
signal \N__64812\ : std_logic;
signal \N__64809\ : std_logic;
signal \N__64806\ : std_logic;
signal \N__64803\ : std_logic;
signal \N__64800\ : std_logic;
signal \N__64795\ : std_logic;
signal \N__64792\ : std_logic;
signal \N__64789\ : std_logic;
signal \N__64786\ : std_logic;
signal \N__64781\ : std_logic;
signal \N__64776\ : std_logic;
signal \N__64771\ : std_logic;
signal \N__64770\ : std_logic;
signal \N__64769\ : std_logic;
signal \N__64764\ : std_logic;
signal \N__64761\ : std_logic;
signal \N__64760\ : std_logic;
signal \N__64757\ : std_logic;
signal \N__64754\ : std_logic;
signal \N__64751\ : std_logic;
signal \N__64748\ : std_logic;
signal \N__64745\ : std_logic;
signal \N__64742\ : std_logic;
signal \N__64739\ : std_logic;
signal \N__64736\ : std_logic;
signal \N__64731\ : std_logic;
signal \N__64728\ : std_logic;
signal \N__64723\ : std_logic;
signal \N__64720\ : std_logic;
signal \N__64717\ : std_logic;
signal \N__64714\ : std_logic;
signal \N__64711\ : std_logic;
signal \N__64708\ : std_logic;
signal \N__64707\ : std_logic;
signal \N__64704\ : std_logic;
signal \N__64703\ : std_logic;
signal \N__64700\ : std_logic;
signal \N__64699\ : std_logic;
signal \N__64696\ : std_logic;
signal \N__64693\ : std_logic;
signal \N__64690\ : std_logic;
signal \N__64687\ : std_logic;
signal \N__64684\ : std_logic;
signal \N__64683\ : std_logic;
signal \N__64680\ : std_logic;
signal \N__64675\ : std_logic;
signal \N__64672\ : std_logic;
signal \N__64669\ : std_logic;
signal \N__64666\ : std_logic;
signal \N__64661\ : std_logic;
signal \N__64658\ : std_logic;
signal \N__64655\ : std_logic;
signal \N__64652\ : std_logic;
signal \N__64645\ : std_logic;
signal \N__64642\ : std_logic;
signal \N__64639\ : std_logic;
signal \N__64636\ : std_logic;
signal \N__64633\ : std_logic;
signal \N__64632\ : std_logic;
signal \N__64629\ : std_logic;
signal \N__64628\ : std_logic;
signal \N__64625\ : std_logic;
signal \N__64624\ : std_logic;
signal \N__64623\ : std_logic;
signal \N__64620\ : std_logic;
signal \N__64617\ : std_logic;
signal \N__64614\ : std_logic;
signal \N__64609\ : std_logic;
signal \N__64608\ : std_logic;
signal \N__64603\ : std_logic;
signal \N__64598\ : std_logic;
signal \N__64595\ : std_logic;
signal \N__64590\ : std_logic;
signal \N__64585\ : std_logic;
signal \N__64584\ : std_logic;
signal \N__64583\ : std_logic;
signal \N__64582\ : std_logic;
signal \N__64579\ : std_logic;
signal \N__64578\ : std_logic;
signal \N__64577\ : std_logic;
signal \N__64574\ : std_logic;
signal \N__64569\ : std_logic;
signal \N__64566\ : std_logic;
signal \N__64565\ : std_logic;
signal \N__64564\ : std_logic;
signal \N__64561\ : std_logic;
signal \N__64558\ : std_logic;
signal \N__64555\ : std_logic;
signal \N__64552\ : std_logic;
signal \N__64551\ : std_logic;
signal \N__64550\ : std_logic;
signal \N__64549\ : std_logic;
signal \N__64548\ : std_logic;
signal \N__64547\ : std_logic;
signal \N__64546\ : std_logic;
signal \N__64543\ : std_logic;
signal \N__64542\ : std_logic;
signal \N__64535\ : std_logic;
signal \N__64530\ : std_logic;
signal \N__64527\ : std_logic;
signal \N__64524\ : std_logic;
signal \N__64519\ : std_logic;
signal \N__64512\ : std_logic;
signal \N__64509\ : std_logic;
signal \N__64506\ : std_logic;
signal \N__64503\ : std_logic;
signal \N__64502\ : std_logic;
signal \N__64499\ : std_logic;
signal \N__64496\ : std_logic;
signal \N__64493\ : std_logic;
signal \N__64486\ : std_logic;
signal \N__64481\ : std_logic;
signal \N__64478\ : std_logic;
signal \N__64475\ : std_logic;
signal \N__64472\ : std_logic;
signal \N__64467\ : std_logic;
signal \N__64464\ : std_logic;
signal \N__64453\ : std_logic;
signal \N__64450\ : std_logic;
signal \N__64449\ : std_logic;
signal \N__64446\ : std_logic;
signal \N__64443\ : std_logic;
signal \N__64442\ : std_logic;
signal \N__64439\ : std_logic;
signal \N__64438\ : std_logic;
signal \N__64435\ : std_logic;
signal \N__64432\ : std_logic;
signal \N__64429\ : std_logic;
signal \N__64426\ : std_logic;
signal \N__64423\ : std_logic;
signal \N__64414\ : std_logic;
signal \N__64413\ : std_logic;
signal \N__64412\ : std_logic;
signal \N__64411\ : std_logic;
signal \N__64410\ : std_logic;
signal \N__64409\ : std_logic;
signal \N__64406\ : std_logic;
signal \N__64401\ : std_logic;
signal \N__64398\ : std_logic;
signal \N__64397\ : std_logic;
signal \N__64394\ : std_logic;
signal \N__64393\ : std_logic;
signal \N__64390\ : std_logic;
signal \N__64389\ : std_logic;
signal \N__64388\ : std_logic;
signal \N__64387\ : std_logic;
signal \N__64386\ : std_logic;
signal \N__64379\ : std_logic;
signal \N__64376\ : std_logic;
signal \N__64373\ : std_logic;
signal \N__64370\ : std_logic;
signal \N__64367\ : std_logic;
signal \N__64366\ : std_logic;
signal \N__64363\ : std_logic;
signal \N__64362\ : std_logic;
signal \N__64355\ : std_logic;
signal \N__64352\ : std_logic;
signal \N__64349\ : std_logic;
signal \N__64346\ : std_logic;
signal \N__64345\ : std_logic;
signal \N__64344\ : std_logic;
signal \N__64341\ : std_logic;
signal \N__64340\ : std_logic;
signal \N__64337\ : std_logic;
signal \N__64330\ : std_logic;
signal \N__64327\ : std_logic;
signal \N__64322\ : std_logic;
signal \N__64319\ : std_logic;
signal \N__64314\ : std_logic;
signal \N__64311\ : std_logic;
signal \N__64308\ : std_logic;
signal \N__64305\ : std_logic;
signal \N__64302\ : std_logic;
signal \N__64299\ : std_logic;
signal \N__64296\ : std_logic;
signal \N__64293\ : std_logic;
signal \N__64290\ : std_logic;
signal \N__64287\ : std_logic;
signal \N__64284\ : std_logic;
signal \N__64279\ : std_logic;
signal \N__64272\ : std_logic;
signal \N__64267\ : std_logic;
signal \N__64264\ : std_logic;
signal \N__64255\ : std_logic;
signal \N__64254\ : std_logic;
signal \N__64253\ : std_logic;
signal \N__64252\ : std_logic;
signal \N__64251\ : std_logic;
signal \N__64250\ : std_logic;
signal \N__64249\ : std_logic;
signal \N__64248\ : std_logic;
signal \N__64247\ : std_logic;
signal \N__64246\ : std_logic;
signal \N__64245\ : std_logic;
signal \N__64244\ : std_logic;
signal \N__64243\ : std_logic;
signal \N__64242\ : std_logic;
signal \N__64239\ : std_logic;
signal \N__64238\ : std_logic;
signal \N__64237\ : std_logic;
signal \N__64228\ : std_logic;
signal \N__64225\ : std_logic;
signal \N__64222\ : std_logic;
signal \N__64221\ : std_logic;
signal \N__64220\ : std_logic;
signal \N__64217\ : std_logic;
signal \N__64210\ : std_logic;
signal \N__64203\ : std_logic;
signal \N__64200\ : std_logic;
signal \N__64199\ : std_logic;
signal \N__64198\ : std_logic;
signal \N__64193\ : std_logic;
signal \N__64188\ : std_logic;
signal \N__64185\ : std_logic;
signal \N__64184\ : std_logic;
signal \N__64183\ : std_logic;
signal \N__64180\ : std_logic;
signal \N__64177\ : std_logic;
signal \N__64174\ : std_logic;
signal \N__64167\ : std_logic;
signal \N__64164\ : std_logic;
signal \N__64161\ : std_logic;
signal \N__64158\ : std_logic;
signal \N__64153\ : std_logic;
signal \N__64148\ : std_logic;
signal \N__64145\ : std_logic;
signal \N__64140\ : std_logic;
signal \N__64137\ : std_logic;
signal \N__64136\ : std_logic;
signal \N__64133\ : std_logic;
signal \N__64130\ : std_logic;
signal \N__64127\ : std_logic;
signal \N__64124\ : std_logic;
signal \N__64121\ : std_logic;
signal \N__64114\ : std_logic;
signal \N__64113\ : std_logic;
signal \N__64110\ : std_logic;
signal \N__64107\ : std_logic;
signal \N__64104\ : std_logic;
signal \N__64101\ : std_logic;
signal \N__64096\ : std_logic;
signal \N__64093\ : std_logic;
signal \N__64090\ : std_logic;
signal \N__64087\ : std_logic;
signal \N__64084\ : std_logic;
signal \N__64081\ : std_logic;
signal \N__64078\ : std_logic;
signal \N__64075\ : std_logic;
signal \N__64072\ : std_logic;
signal \N__64057\ : std_logic;
signal \N__64056\ : std_logic;
signal \N__64053\ : std_logic;
signal \N__64050\ : std_logic;
signal \N__64049\ : std_logic;
signal \N__64046\ : std_logic;
signal \N__64043\ : std_logic;
signal \N__64040\ : std_logic;
signal \N__64039\ : std_logic;
signal \N__64036\ : std_logic;
signal \N__64033\ : std_logic;
signal \N__64028\ : std_logic;
signal \N__64021\ : std_logic;
signal \N__64018\ : std_logic;
signal \N__64015\ : std_logic;
signal \N__64014\ : std_logic;
signal \N__64013\ : std_logic;
signal \N__64010\ : std_logic;
signal \N__64007\ : std_logic;
signal \N__64004\ : std_logic;
signal \N__64003\ : std_logic;
signal \N__64002\ : std_logic;
signal \N__63999\ : std_logic;
signal \N__63996\ : std_logic;
signal \N__63995\ : std_logic;
signal \N__63994\ : std_logic;
signal \N__63991\ : std_logic;
signal \N__63988\ : std_logic;
signal \N__63985\ : std_logic;
signal \N__63982\ : std_logic;
signal \N__63979\ : std_logic;
signal \N__63974\ : std_logic;
signal \N__63971\ : std_logic;
signal \N__63968\ : std_logic;
signal \N__63955\ : std_logic;
signal \N__63952\ : std_logic;
signal \N__63949\ : std_logic;
signal \N__63948\ : std_logic;
signal \N__63945\ : std_logic;
signal \N__63944\ : std_logic;
signal \N__63943\ : std_logic;
signal \N__63940\ : std_logic;
signal \N__63939\ : std_logic;
signal \N__63938\ : std_logic;
signal \N__63937\ : std_logic;
signal \N__63934\ : std_logic;
signal \N__63931\ : std_logic;
signal \N__63928\ : std_logic;
signal \N__63925\ : std_logic;
signal \N__63922\ : std_logic;
signal \N__63919\ : std_logic;
signal \N__63916\ : std_logic;
signal \N__63915\ : std_logic;
signal \N__63910\ : std_logic;
signal \N__63907\ : std_logic;
signal \N__63900\ : std_logic;
signal \N__63897\ : std_logic;
signal \N__63894\ : std_logic;
signal \N__63891\ : std_logic;
signal \N__63888\ : std_logic;
signal \N__63885\ : std_logic;
signal \N__63880\ : std_logic;
signal \N__63871\ : std_logic;
signal \N__63870\ : std_logic;
signal \N__63865\ : std_logic;
signal \N__63862\ : std_logic;
signal \N__63861\ : std_logic;
signal \N__63858\ : std_logic;
signal \N__63855\ : std_logic;
signal \N__63854\ : std_logic;
signal \N__63853\ : std_logic;
signal \N__63850\ : std_logic;
signal \N__63847\ : std_logic;
signal \N__63844\ : std_logic;
signal \N__63843\ : std_logic;
signal \N__63840\ : std_logic;
signal \N__63837\ : std_logic;
signal \N__63834\ : std_logic;
signal \N__63831\ : std_logic;
signal \N__63828\ : std_logic;
signal \N__63825\ : std_logic;
signal \N__63822\ : std_logic;
signal \N__63819\ : std_logic;
signal \N__63814\ : std_logic;
signal \N__63805\ : std_logic;
signal \N__63802\ : std_logic;
signal \N__63799\ : std_logic;
signal \N__63796\ : std_logic;
signal \N__63795\ : std_logic;
signal \N__63794\ : std_logic;
signal \N__63791\ : std_logic;
signal \N__63786\ : std_logic;
signal \N__63781\ : std_logic;
signal \N__63778\ : std_logic;
signal \N__63777\ : std_logic;
signal \N__63776\ : std_logic;
signal \N__63775\ : std_logic;
signal \N__63774\ : std_logic;
signal \N__63771\ : std_logic;
signal \N__63768\ : std_logic;
signal \N__63767\ : std_logic;
signal \N__63766\ : std_logic;
signal \N__63765\ : std_logic;
signal \N__63762\ : std_logic;
signal \N__63759\ : std_logic;
signal \N__63756\ : std_logic;
signal \N__63753\ : std_logic;
signal \N__63748\ : std_logic;
signal \N__63743\ : std_logic;
signal \N__63742\ : std_logic;
signal \N__63741\ : std_logic;
signal \N__63736\ : std_logic;
signal \N__63733\ : std_logic;
signal \N__63728\ : std_logic;
signal \N__63725\ : std_logic;
signal \N__63720\ : std_logic;
signal \N__63715\ : std_logic;
signal \N__63712\ : std_logic;
signal \N__63709\ : std_logic;
signal \N__63700\ : std_logic;
signal \N__63697\ : std_logic;
signal \N__63694\ : std_logic;
signal \N__63691\ : std_logic;
signal \N__63688\ : std_logic;
signal \N__63687\ : std_logic;
signal \N__63684\ : std_logic;
signal \N__63683\ : std_logic;
signal \N__63680\ : std_logic;
signal \N__63679\ : std_logic;
signal \N__63678\ : std_logic;
signal \N__63673\ : std_logic;
signal \N__63670\ : std_logic;
signal \N__63665\ : std_logic;
signal \N__63658\ : std_logic;
signal \N__63655\ : std_logic;
signal \N__63652\ : std_logic;
signal \N__63651\ : std_logic;
signal \N__63648\ : std_logic;
signal \N__63647\ : std_logic;
signal \N__63646\ : std_logic;
signal \N__63643\ : std_logic;
signal \N__63640\ : std_logic;
signal \N__63637\ : std_logic;
signal \N__63634\ : std_logic;
signal \N__63631\ : std_logic;
signal \N__63630\ : std_logic;
signal \N__63629\ : std_logic;
signal \N__63628\ : std_logic;
signal \N__63627\ : std_logic;
signal \N__63622\ : std_logic;
signal \N__63619\ : std_logic;
signal \N__63616\ : std_logic;
signal \N__63611\ : std_logic;
signal \N__63608\ : std_logic;
signal \N__63605\ : std_logic;
signal \N__63602\ : std_logic;
signal \N__63597\ : std_logic;
signal \N__63590\ : std_logic;
signal \N__63583\ : std_logic;
signal \N__63580\ : std_logic;
signal \N__63577\ : std_logic;
signal \N__63576\ : std_logic;
signal \N__63575\ : std_logic;
signal \N__63574\ : std_logic;
signal \N__63573\ : std_logic;
signal \N__63570\ : std_logic;
signal \N__63567\ : std_logic;
signal \N__63564\ : std_logic;
signal \N__63561\ : std_logic;
signal \N__63560\ : std_logic;
signal \N__63557\ : std_logic;
signal \N__63552\ : std_logic;
signal \N__63549\ : std_logic;
signal \N__63546\ : std_logic;
signal \N__63543\ : std_logic;
signal \N__63540\ : std_logic;
signal \N__63535\ : std_logic;
signal \N__63534\ : std_logic;
signal \N__63529\ : std_logic;
signal \N__63526\ : std_logic;
signal \N__63523\ : std_logic;
signal \N__63520\ : std_logic;
signal \N__63517\ : std_logic;
signal \N__63512\ : std_logic;
signal \N__63509\ : std_logic;
signal \N__63506\ : std_logic;
signal \N__63503\ : std_logic;
signal \N__63496\ : std_logic;
signal \N__63495\ : std_logic;
signal \N__63494\ : std_logic;
signal \N__63489\ : std_logic;
signal \N__63486\ : std_logic;
signal \N__63485\ : std_logic;
signal \N__63482\ : std_logic;
signal \N__63479\ : std_logic;
signal \N__63476\ : std_logic;
signal \N__63473\ : std_logic;
signal \N__63468\ : std_logic;
signal \N__63465\ : std_logic;
signal \N__63462\ : std_logic;
signal \N__63457\ : std_logic;
signal \N__63456\ : std_logic;
signal \N__63455\ : std_logic;
signal \N__63452\ : std_logic;
signal \N__63449\ : std_logic;
signal \N__63446\ : std_logic;
signal \N__63441\ : std_logic;
signal \N__63438\ : std_logic;
signal \N__63435\ : std_logic;
signal \N__63432\ : std_logic;
signal \N__63429\ : std_logic;
signal \N__63426\ : std_logic;
signal \N__63423\ : std_logic;
signal \N__63418\ : std_logic;
signal \N__63417\ : std_logic;
signal \N__63416\ : std_logic;
signal \N__63415\ : std_logic;
signal \N__63414\ : std_logic;
signal \N__63413\ : std_logic;
signal \N__63412\ : std_logic;
signal \N__63409\ : std_logic;
signal \N__63404\ : std_logic;
signal \N__63399\ : std_logic;
signal \N__63396\ : std_logic;
signal \N__63395\ : std_logic;
signal \N__63394\ : std_logic;
signal \N__63391\ : std_logic;
signal \N__63390\ : std_logic;
signal \N__63389\ : std_logic;
signal \N__63386\ : std_logic;
signal \N__63381\ : std_logic;
signal \N__63380\ : std_logic;
signal \N__63379\ : std_logic;
signal \N__63378\ : std_logic;
signal \N__63377\ : std_logic;
signal \N__63374\ : std_logic;
signal \N__63371\ : std_logic;
signal \N__63368\ : std_logic;
signal \N__63365\ : std_logic;
signal \N__63362\ : std_logic;
signal \N__63359\ : std_logic;
signal \N__63358\ : std_logic;
signal \N__63357\ : std_logic;
signal \N__63356\ : std_logic;
signal \N__63355\ : std_logic;
signal \N__63354\ : std_logic;
signal \N__63353\ : std_logic;
signal \N__63348\ : std_logic;
signal \N__63343\ : std_logic;
signal \N__63340\ : std_logic;
signal \N__63337\ : std_logic;
signal \N__63334\ : std_logic;
signal \N__63331\ : std_logic;
signal \N__63328\ : std_logic;
signal \N__63325\ : std_logic;
signal \N__63318\ : std_logic;
signal \N__63315\ : std_logic;
signal \N__63312\ : std_logic;
signal \N__63305\ : std_logic;
signal \N__63300\ : std_logic;
signal \N__63295\ : std_logic;
signal \N__63292\ : std_logic;
signal \N__63287\ : std_logic;
signal \N__63282\ : std_logic;
signal \N__63281\ : std_logic;
signal \N__63280\ : std_logic;
signal \N__63273\ : std_logic;
signal \N__63270\ : std_logic;
signal \N__63265\ : std_logic;
signal \N__63260\ : std_logic;
signal \N__63257\ : std_logic;
signal \N__63254\ : std_logic;
signal \N__63251\ : std_logic;
signal \N__63246\ : std_logic;
signal \N__63243\ : std_logic;
signal \N__63232\ : std_logic;
signal \N__63231\ : std_logic;
signal \N__63228\ : std_logic;
signal \N__63225\ : std_logic;
signal \N__63224\ : std_logic;
signal \N__63219\ : std_logic;
signal \N__63218\ : std_logic;
signal \N__63215\ : std_logic;
signal \N__63212\ : std_logic;
signal \N__63209\ : std_logic;
signal \N__63202\ : std_logic;
signal \N__63201\ : std_logic;
signal \N__63198\ : std_logic;
signal \N__63197\ : std_logic;
signal \N__63194\ : std_logic;
signal \N__63191\ : std_logic;
signal \N__63188\ : std_logic;
signal \N__63181\ : std_logic;
signal \N__63180\ : std_logic;
signal \N__63175\ : std_logic;
signal \N__63172\ : std_logic;
signal \N__63169\ : std_logic;
signal \N__63166\ : std_logic;
signal \N__63163\ : std_logic;
signal \N__63162\ : std_logic;
signal \N__63159\ : std_logic;
signal \N__63156\ : std_logic;
signal \N__63155\ : std_logic;
signal \N__63150\ : std_logic;
signal \N__63149\ : std_logic;
signal \N__63148\ : std_logic;
signal \N__63145\ : std_logic;
signal \N__63142\ : std_logic;
signal \N__63139\ : std_logic;
signal \N__63136\ : std_logic;
signal \N__63135\ : std_logic;
signal \N__63132\ : std_logic;
signal \N__63129\ : std_logic;
signal \N__63124\ : std_logic;
signal \N__63121\ : std_logic;
signal \N__63118\ : std_logic;
signal \N__63109\ : std_logic;
signal \N__63106\ : std_logic;
signal \N__63105\ : std_logic;
signal \N__63104\ : std_logic;
signal \N__63101\ : std_logic;
signal \N__63100\ : std_logic;
signal \N__63099\ : std_logic;
signal \N__63096\ : std_logic;
signal \N__63093\ : std_logic;
signal \N__63090\ : std_logic;
signal \N__63087\ : std_logic;
signal \N__63084\ : std_logic;
signal \N__63081\ : std_logic;
signal \N__63070\ : std_logic;
signal \N__63067\ : std_logic;
signal \N__63066\ : std_logic;
signal \N__63065\ : std_logic;
signal \N__63062\ : std_logic;
signal \N__63057\ : std_logic;
signal \N__63054\ : std_logic;
signal \N__63049\ : std_logic;
signal \N__63048\ : std_logic;
signal \N__63045\ : std_logic;
signal \N__63044\ : std_logic;
signal \N__63041\ : std_logic;
signal \N__63038\ : std_logic;
signal \N__63035\ : std_logic;
signal \N__63034\ : std_logic;
signal \N__63031\ : std_logic;
signal \N__63028\ : std_logic;
signal \N__63025\ : std_logic;
signal \N__63022\ : std_logic;
signal \N__63013\ : std_logic;
signal \N__63010\ : std_logic;
signal \N__63007\ : std_logic;
signal \N__63004\ : std_logic;
signal \N__63001\ : std_logic;
signal \N__62998\ : std_logic;
signal \N__62995\ : std_logic;
signal \N__62992\ : std_logic;
signal \N__62989\ : std_logic;
signal \N__62988\ : std_logic;
signal \N__62985\ : std_logic;
signal \N__62982\ : std_logic;
signal \N__62981\ : std_logic;
signal \N__62976\ : std_logic;
signal \N__62973\ : std_logic;
signal \N__62970\ : std_logic;
signal \N__62969\ : std_logic;
signal \N__62968\ : std_logic;
signal \N__62965\ : std_logic;
signal \N__62962\ : std_logic;
signal \N__62957\ : std_logic;
signal \N__62950\ : std_logic;
signal \N__62947\ : std_logic;
signal \N__62944\ : std_logic;
signal \N__62941\ : std_logic;
signal \N__62938\ : std_logic;
signal \N__62935\ : std_logic;
signal \N__62934\ : std_logic;
signal \N__62931\ : std_logic;
signal \N__62928\ : std_logic;
signal \N__62927\ : std_logic;
signal \N__62926\ : std_logic;
signal \N__62923\ : std_logic;
signal \N__62916\ : std_logic;
signal \N__62911\ : std_logic;
signal \N__62908\ : std_logic;
signal \N__62905\ : std_logic;
signal \N__62904\ : std_logic;
signal \N__62901\ : std_logic;
signal \N__62898\ : std_logic;
signal \N__62895\ : std_logic;
signal \N__62890\ : std_logic;
signal \N__62889\ : std_logic;
signal \N__62886\ : std_logic;
signal \N__62885\ : std_logic;
signal \N__62882\ : std_logic;
signal \N__62879\ : std_logic;
signal \N__62878\ : std_logic;
signal \N__62875\ : std_logic;
signal \N__62872\ : std_logic;
signal \N__62869\ : std_logic;
signal \N__62866\ : std_logic;
signal \N__62863\ : std_logic;
signal \N__62858\ : std_logic;
signal \N__62855\ : std_logic;
signal \N__62848\ : std_logic;
signal \N__62847\ : std_logic;
signal \N__62846\ : std_logic;
signal \N__62845\ : std_logic;
signal \N__62844\ : std_logic;
signal \N__62839\ : std_logic;
signal \N__62838\ : std_logic;
signal \N__62837\ : std_logic;
signal \N__62834\ : std_logic;
signal \N__62831\ : std_logic;
signal \N__62830\ : std_logic;
signal \N__62827\ : std_logic;
signal \N__62824\ : std_logic;
signal \N__62819\ : std_logic;
signal \N__62816\ : std_logic;
signal \N__62813\ : std_logic;
signal \N__62812\ : std_logic;
signal \N__62811\ : std_logic;
signal \N__62810\ : std_logic;
signal \N__62807\ : std_logic;
signal \N__62804\ : std_logic;
signal \N__62803\ : std_logic;
signal \N__62802\ : std_logic;
signal \N__62801\ : std_logic;
signal \N__62798\ : std_logic;
signal \N__62795\ : std_logic;
signal \N__62794\ : std_logic;
signal \N__62793\ : std_logic;
signal \N__62788\ : std_logic;
signal \N__62785\ : std_logic;
signal \N__62782\ : std_logic;
signal \N__62779\ : std_logic;
signal \N__62774\ : std_logic;
signal \N__62771\ : std_logic;
signal \N__62766\ : std_logic;
signal \N__62763\ : std_logic;
signal \N__62760\ : std_logic;
signal \N__62755\ : std_logic;
signal \N__62752\ : std_logic;
signal \N__62743\ : std_logic;
signal \N__62734\ : std_logic;
signal \N__62725\ : std_logic;
signal \N__62724\ : std_logic;
signal \N__62721\ : std_logic;
signal \N__62720\ : std_logic;
signal \N__62717\ : std_logic;
signal \N__62716\ : std_logic;
signal \N__62713\ : std_logic;
signal \N__62710\ : std_logic;
signal \N__62705\ : std_logic;
signal \N__62698\ : std_logic;
signal \N__62695\ : std_logic;
signal \N__62692\ : std_logic;
signal \N__62689\ : std_logic;
signal \N__62686\ : std_logic;
signal \N__62683\ : std_logic;
signal \N__62682\ : std_logic;
signal \N__62681\ : std_logic;
signal \N__62680\ : std_logic;
signal \N__62679\ : std_logic;
signal \N__62676\ : std_logic;
signal \N__62673\ : std_logic;
signal \N__62670\ : std_logic;
signal \N__62667\ : std_logic;
signal \N__62664\ : std_logic;
signal \N__62659\ : std_logic;
signal \N__62658\ : std_logic;
signal \N__62655\ : std_logic;
signal \N__62650\ : std_logic;
signal \N__62647\ : std_logic;
signal \N__62644\ : std_logic;
signal \N__62635\ : std_logic;
signal \N__62632\ : std_logic;
signal \N__62629\ : std_logic;
signal \N__62626\ : std_logic;
signal \N__62625\ : std_logic;
signal \N__62624\ : std_logic;
signal \N__62621\ : std_logic;
signal \N__62620\ : std_logic;
signal \N__62619\ : std_logic;
signal \N__62618\ : std_logic;
signal \N__62615\ : std_logic;
signal \N__62612\ : std_logic;
signal \N__62609\ : std_logic;
signal \N__62606\ : std_logic;
signal \N__62601\ : std_logic;
signal \N__62596\ : std_logic;
signal \N__62587\ : std_logic;
signal \N__62584\ : std_logic;
signal \N__62583\ : std_logic;
signal \N__62582\ : std_logic;
signal \N__62579\ : std_logic;
signal \N__62576\ : std_logic;
signal \N__62573\ : std_logic;
signal \N__62570\ : std_logic;
signal \N__62567\ : std_logic;
signal \N__62564\ : std_logic;
signal \N__62561\ : std_logic;
signal \N__62556\ : std_logic;
signal \N__62551\ : std_logic;
signal \N__62548\ : std_logic;
signal \N__62545\ : std_logic;
signal \N__62544\ : std_logic;
signal \N__62541\ : std_logic;
signal \N__62538\ : std_logic;
signal \N__62535\ : std_logic;
signal \N__62532\ : std_logic;
signal \N__62527\ : std_logic;
signal \N__62524\ : std_logic;
signal \N__62523\ : std_logic;
signal \N__62522\ : std_logic;
signal \N__62519\ : std_logic;
signal \N__62516\ : std_logic;
signal \N__62513\ : std_logic;
signal \N__62512\ : std_logic;
signal \N__62507\ : std_logic;
signal \N__62502\ : std_logic;
signal \N__62497\ : std_logic;
signal \N__62496\ : std_logic;
signal \N__62495\ : std_logic;
signal \N__62492\ : std_logic;
signal \N__62489\ : std_logic;
signal \N__62486\ : std_logic;
signal \N__62483\ : std_logic;
signal \N__62480\ : std_logic;
signal \N__62477\ : std_logic;
signal \N__62474\ : std_logic;
signal \N__62467\ : std_logic;
signal \N__62466\ : std_logic;
signal \N__62465\ : std_logic;
signal \N__62464\ : std_logic;
signal \N__62461\ : std_logic;
signal \N__62456\ : std_logic;
signal \N__62453\ : std_logic;
signal \N__62448\ : std_logic;
signal \N__62447\ : std_logic;
signal \N__62444\ : std_logic;
signal \N__62441\ : std_logic;
signal \N__62440\ : std_logic;
signal \N__62437\ : std_logic;
signal \N__62434\ : std_logic;
signal \N__62431\ : std_logic;
signal \N__62428\ : std_logic;
signal \N__62419\ : std_logic;
signal \N__62418\ : std_logic;
signal \N__62415\ : std_logic;
signal \N__62412\ : std_logic;
signal \N__62411\ : std_logic;
signal \N__62410\ : std_logic;
signal \N__62409\ : std_logic;
signal \N__62406\ : std_logic;
signal \N__62403\ : std_logic;
signal \N__62400\ : std_logic;
signal \N__62399\ : std_logic;
signal \N__62396\ : std_logic;
signal \N__62393\ : std_logic;
signal \N__62386\ : std_logic;
signal \N__62383\ : std_logic;
signal \N__62382\ : std_logic;
signal \N__62379\ : std_logic;
signal \N__62374\ : std_logic;
signal \N__62371\ : std_logic;
signal \N__62368\ : std_logic;
signal \N__62359\ : std_logic;
signal \N__62356\ : std_logic;
signal \N__62355\ : std_logic;
signal \N__62354\ : std_logic;
signal \N__62353\ : std_logic;
signal \N__62350\ : std_logic;
signal \N__62347\ : std_logic;
signal \N__62344\ : std_logic;
signal \N__62343\ : std_logic;
signal \N__62340\ : std_logic;
signal \N__62335\ : std_logic;
signal \N__62332\ : std_logic;
signal \N__62329\ : std_logic;
signal \N__62320\ : std_logic;
signal \N__62317\ : std_logic;
signal \N__62314\ : std_logic;
signal \N__62313\ : std_logic;
signal \N__62310\ : std_logic;
signal \N__62309\ : std_logic;
signal \N__62308\ : std_logic;
signal \N__62307\ : std_logic;
signal \N__62304\ : std_logic;
signal \N__62301\ : std_logic;
signal \N__62298\ : std_logic;
signal \N__62293\ : std_logic;
signal \N__62290\ : std_logic;
signal \N__62287\ : std_logic;
signal \N__62284\ : std_logic;
signal \N__62281\ : std_logic;
signal \N__62278\ : std_logic;
signal \N__62275\ : std_logic;
signal \N__62270\ : std_logic;
signal \N__62267\ : std_logic;
signal \N__62264\ : std_logic;
signal \N__62257\ : std_logic;
signal \N__62256\ : std_logic;
signal \N__62255\ : std_logic;
signal \N__62254\ : std_logic;
signal \N__62251\ : std_logic;
signal \N__62250\ : std_logic;
signal \N__62247\ : std_logic;
signal \N__62244\ : std_logic;
signal \N__62241\ : std_logic;
signal \N__62238\ : std_logic;
signal \N__62235\ : std_logic;
signal \N__62232\ : std_logic;
signal \N__62229\ : std_logic;
signal \N__62226\ : std_logic;
signal \N__62223\ : std_logic;
signal \N__62218\ : std_logic;
signal \N__62215\ : std_logic;
signal \N__62206\ : std_logic;
signal \N__62203\ : std_logic;
signal \N__62200\ : std_logic;
signal \N__62199\ : std_logic;
signal \N__62198\ : std_logic;
signal \N__62197\ : std_logic;
signal \N__62194\ : std_logic;
signal \N__62187\ : std_logic;
signal \N__62182\ : std_logic;
signal \N__62181\ : std_logic;
signal \N__62180\ : std_logic;
signal \N__62177\ : std_logic;
signal \N__62176\ : std_logic;
signal \N__62173\ : std_logic;
signal \N__62172\ : std_logic;
signal \N__62169\ : std_logic;
signal \N__62166\ : std_logic;
signal \N__62165\ : std_logic;
signal \N__62164\ : std_logic;
signal \N__62163\ : std_logic;
signal \N__62160\ : std_logic;
signal \N__62157\ : std_logic;
signal \N__62156\ : std_logic;
signal \N__62153\ : std_logic;
signal \N__62148\ : std_logic;
signal \N__62145\ : std_logic;
signal \N__62140\ : std_logic;
signal \N__62135\ : std_logic;
signal \N__62132\ : std_logic;
signal \N__62131\ : std_logic;
signal \N__62130\ : std_logic;
signal \N__62129\ : std_logic;
signal \N__62128\ : std_logic;
signal \N__62127\ : std_logic;
signal \N__62126\ : std_logic;
signal \N__62123\ : std_logic;
signal \N__62118\ : std_logic;
signal \N__62111\ : std_logic;
signal \N__62108\ : std_logic;
signal \N__62105\ : std_logic;
signal \N__62100\ : std_logic;
signal \N__62095\ : std_logic;
signal \N__62080\ : std_logic;
signal \N__62077\ : std_logic;
signal \N__62076\ : std_logic;
signal \N__62073\ : std_logic;
signal \N__62070\ : std_logic;
signal \N__62067\ : std_logic;
signal \N__62062\ : std_logic;
signal \N__62059\ : std_logic;
signal \N__62058\ : std_logic;
signal \N__62053\ : std_logic;
signal \N__62050\ : std_logic;
signal \N__62049\ : std_logic;
signal \N__62048\ : std_logic;
signal \N__62045\ : std_logic;
signal \N__62042\ : std_logic;
signal \N__62041\ : std_logic;
signal \N__62040\ : std_logic;
signal \N__62039\ : std_logic;
signal \N__62036\ : std_logic;
signal \N__62035\ : std_logic;
signal \N__62034\ : std_logic;
signal \N__62031\ : std_logic;
signal \N__62030\ : std_logic;
signal \N__62027\ : std_logic;
signal \N__62024\ : std_logic;
signal \N__62019\ : std_logic;
signal \N__62018\ : std_logic;
signal \N__62013\ : std_logic;
signal \N__62010\ : std_logic;
signal \N__62009\ : std_logic;
signal \N__62006\ : std_logic;
signal \N__62003\ : std_logic;
signal \N__62002\ : std_logic;
signal \N__61997\ : std_logic;
signal \N__61994\ : std_logic;
signal \N__61991\ : std_logic;
signal \N__61988\ : std_logic;
signal \N__61987\ : std_logic;
signal \N__61984\ : std_logic;
signal \N__61981\ : std_logic;
signal \N__61976\ : std_logic;
signal \N__61973\ : std_logic;
signal \N__61968\ : std_logic;
signal \N__61965\ : std_logic;
signal \N__61962\ : std_logic;
signal \N__61959\ : std_logic;
signal \N__61956\ : std_logic;
signal \N__61955\ : std_logic;
signal \N__61954\ : std_logic;
signal \N__61951\ : std_logic;
signal \N__61948\ : std_logic;
signal \N__61945\ : std_logic;
signal \N__61942\ : std_logic;
signal \N__61937\ : std_logic;
signal \N__61934\ : std_logic;
signal \N__61931\ : std_logic;
signal \N__61928\ : std_logic;
signal \N__61927\ : std_logic;
signal \N__61924\ : std_logic;
signal \N__61921\ : std_logic;
signal \N__61916\ : std_logic;
signal \N__61911\ : std_logic;
signal \N__61904\ : std_logic;
signal \N__61901\ : std_logic;
signal \N__61898\ : std_logic;
signal \N__61893\ : std_logic;
signal \N__61888\ : std_logic;
signal \N__61879\ : std_logic;
signal \N__61878\ : std_logic;
signal \N__61875\ : std_logic;
signal \N__61874\ : std_logic;
signal \N__61873\ : std_logic;
signal \N__61872\ : std_logic;
signal \N__61871\ : std_logic;
signal \N__61868\ : std_logic;
signal \N__61865\ : std_logic;
signal \N__61862\ : std_logic;
signal \N__61861\ : std_logic;
signal \N__61860\ : std_logic;
signal \N__61857\ : std_logic;
signal \N__61852\ : std_logic;
signal \N__61847\ : std_logic;
signal \N__61844\ : std_logic;
signal \N__61841\ : std_logic;
signal \N__61838\ : std_logic;
signal \N__61833\ : std_logic;
signal \N__61830\ : std_logic;
signal \N__61827\ : std_logic;
signal \N__61826\ : std_logic;
signal \N__61823\ : std_logic;
signal \N__61820\ : std_logic;
signal \N__61813\ : std_logic;
signal \N__61810\ : std_logic;
signal \N__61801\ : std_logic;
signal \N__61798\ : std_logic;
signal \N__61797\ : std_logic;
signal \N__61796\ : std_logic;
signal \N__61795\ : std_logic;
signal \N__61794\ : std_logic;
signal \N__61791\ : std_logic;
signal \N__61786\ : std_logic;
signal \N__61781\ : std_logic;
signal \N__61780\ : std_logic;
signal \N__61779\ : std_logic;
signal \N__61778\ : std_logic;
signal \N__61777\ : std_logic;
signal \N__61774\ : std_logic;
signal \N__61769\ : std_logic;
signal \N__61768\ : std_logic;
signal \N__61767\ : std_logic;
signal \N__61766\ : std_logic;
signal \N__61761\ : std_logic;
signal \N__61760\ : std_logic;
signal \N__61759\ : std_logic;
signal \N__61758\ : std_logic;
signal \N__61757\ : std_logic;
signal \N__61756\ : std_logic;
signal \N__61755\ : std_logic;
signal \N__61754\ : std_logic;
signal \N__61753\ : std_logic;
signal \N__61752\ : std_logic;
signal \N__61749\ : std_logic;
signal \N__61746\ : std_logic;
signal \N__61745\ : std_logic;
signal \N__61744\ : std_logic;
signal \N__61739\ : std_logic;
signal \N__61732\ : std_logic;
signal \N__61731\ : std_logic;
signal \N__61730\ : std_logic;
signal \N__61727\ : std_logic;
signal \N__61726\ : std_logic;
signal \N__61725\ : std_logic;
signal \N__61724\ : std_logic;
signal \N__61723\ : std_logic;
signal \N__61716\ : std_logic;
signal \N__61713\ : std_logic;
signal \N__61702\ : std_logic;
signal \N__61693\ : std_logic;
signal \N__61692\ : std_logic;
signal \N__61691\ : std_logic;
signal \N__61690\ : std_logic;
signal \N__61689\ : std_logic;
signal \N__61688\ : std_logic;
signal \N__61687\ : std_logic;
signal \N__61686\ : std_logic;
signal \N__61685\ : std_logic;
signal \N__61684\ : std_logic;
signal \N__61683\ : std_logic;
signal \N__61678\ : std_logic;
signal \N__61677\ : std_logic;
signal \N__61674\ : std_logic;
signal \N__61673\ : std_logic;
signal \N__61672\ : std_logic;
signal \N__61671\ : std_logic;
signal \N__61670\ : std_logic;
signal \N__61667\ : std_logic;
signal \N__61664\ : std_logic;
signal \N__61659\ : std_logic;
signal \N__61654\ : std_logic;
signal \N__61651\ : std_logic;
signal \N__61644\ : std_logic;
signal \N__61635\ : std_logic;
signal \N__61632\ : std_logic;
signal \N__61627\ : std_logic;
signal \N__61624\ : std_logic;
signal \N__61619\ : std_logic;
signal \N__61616\ : std_logic;
signal \N__61615\ : std_logic;
signal \N__61612\ : std_logic;
signal \N__61609\ : std_logic;
signal \N__61600\ : std_logic;
signal \N__61599\ : std_logic;
signal \N__61598\ : std_logic;
signal \N__61597\ : std_logic;
signal \N__61596\ : std_logic;
signal \N__61595\ : std_logic;
signal \N__61594\ : std_logic;
signal \N__61593\ : std_logic;
signal \N__61584\ : std_logic;
signal \N__61577\ : std_logic;
signal \N__61572\ : std_logic;
signal \N__61567\ : std_logic;
signal \N__61564\ : std_logic;
signal \N__61561\ : std_logic;
signal \N__61560\ : std_logic;
signal \N__61553\ : std_logic;
signal \N__61552\ : std_logic;
signal \N__61551\ : std_logic;
signal \N__61550\ : std_logic;
signal \N__61549\ : std_logic;
signal \N__61546\ : std_logic;
signal \N__61543\ : std_logic;
signal \N__61538\ : std_logic;
signal \N__61531\ : std_logic;
signal \N__61522\ : std_logic;
signal \N__61519\ : std_logic;
signal \N__61516\ : std_logic;
signal \N__61513\ : std_logic;
signal \N__61510\ : std_logic;
signal \N__61501\ : std_logic;
signal \N__61498\ : std_logic;
signal \N__61485\ : std_logic;
signal \N__61478\ : std_logic;
signal \N__61475\ : std_logic;
signal \N__61472\ : std_logic;
signal \N__61469\ : std_logic;
signal \N__61466\ : std_logic;
signal \N__61461\ : std_logic;
signal \N__61456\ : std_logic;
signal \N__61455\ : std_logic;
signal \N__61454\ : std_logic;
signal \N__61453\ : std_logic;
signal \N__61450\ : std_logic;
signal \N__61449\ : std_logic;
signal \N__61448\ : std_logic;
signal \N__61443\ : std_logic;
signal \N__61440\ : std_logic;
signal \N__61437\ : std_logic;
signal \N__61434\ : std_logic;
signal \N__61431\ : std_logic;
signal \N__61430\ : std_logic;
signal \N__61425\ : std_logic;
signal \N__61424\ : std_logic;
signal \N__61421\ : std_logic;
signal \N__61418\ : std_logic;
signal \N__61415\ : std_logic;
signal \N__61412\ : std_logic;
signal \N__61409\ : std_logic;
signal \N__61408\ : std_logic;
signal \N__61407\ : std_logic;
signal \N__61404\ : std_logic;
signal \N__61401\ : std_logic;
signal \N__61398\ : std_logic;
signal \N__61395\ : std_logic;
signal \N__61392\ : std_logic;
signal \N__61389\ : std_logic;
signal \N__61384\ : std_logic;
signal \N__61381\ : std_logic;
signal \N__61378\ : std_logic;
signal \N__61373\ : std_logic;
signal \N__61368\ : std_logic;
signal \N__61361\ : std_logic;
signal \N__61354\ : std_logic;
signal \N__61351\ : std_logic;
signal \N__61348\ : std_logic;
signal \N__61347\ : std_logic;
signal \N__61346\ : std_logic;
signal \N__61345\ : std_logic;
signal \N__61342\ : std_logic;
signal \N__61337\ : std_logic;
signal \N__61334\ : std_logic;
signal \N__61331\ : std_logic;
signal \N__61328\ : std_logic;
signal \N__61327\ : std_logic;
signal \N__61326\ : std_logic;
signal \N__61323\ : std_logic;
signal \N__61318\ : std_logic;
signal \N__61313\ : std_logic;
signal \N__61306\ : std_logic;
signal \N__61303\ : std_logic;
signal \N__61300\ : std_logic;
signal \N__61297\ : std_logic;
signal \N__61294\ : std_logic;
signal \N__61291\ : std_logic;
signal \N__61288\ : std_logic;
signal \N__61285\ : std_logic;
signal \N__61284\ : std_logic;
signal \N__61281\ : std_logic;
signal \N__61278\ : std_logic;
signal \N__61275\ : std_logic;
signal \N__61272\ : std_logic;
signal \N__61269\ : std_logic;
signal \N__61266\ : std_logic;
signal \N__61261\ : std_logic;
signal \N__61258\ : std_logic;
signal \N__61255\ : std_logic;
signal \N__61254\ : std_logic;
signal \N__61251\ : std_logic;
signal \N__61248\ : std_logic;
signal \N__61247\ : std_logic;
signal \N__61246\ : std_logic;
signal \N__61241\ : std_logic;
signal \N__61236\ : std_logic;
signal \N__61231\ : std_logic;
signal \N__61228\ : std_logic;
signal \N__61227\ : std_logic;
signal \N__61226\ : std_logic;
signal \N__61225\ : std_logic;
signal \N__61222\ : std_logic;
signal \N__61219\ : std_logic;
signal \N__61216\ : std_logic;
signal \N__61213\ : std_logic;
signal \N__61212\ : std_logic;
signal \N__61209\ : std_logic;
signal \N__61206\ : std_logic;
signal \N__61205\ : std_logic;
signal \N__61202\ : std_logic;
signal \N__61199\ : std_logic;
signal \N__61198\ : std_logic;
signal \N__61197\ : std_logic;
signal \N__61196\ : std_logic;
signal \N__61195\ : std_logic;
signal \N__61194\ : std_logic;
signal \N__61193\ : std_logic;
signal \N__61190\ : std_logic;
signal \N__61187\ : std_logic;
signal \N__61184\ : std_logic;
signal \N__61181\ : std_logic;
signal \N__61176\ : std_logic;
signal \N__61173\ : std_logic;
signal \N__61170\ : std_logic;
signal \N__61163\ : std_logic;
signal \N__61160\ : std_logic;
signal \N__61141\ : std_logic;
signal \N__61138\ : std_logic;
signal \N__61135\ : std_logic;
signal \N__61132\ : std_logic;
signal \N__61131\ : std_logic;
signal \N__61128\ : std_logic;
signal \N__61127\ : std_logic;
signal \N__61126\ : std_logic;
signal \N__61123\ : std_logic;
signal \N__61122\ : std_logic;
signal \N__61119\ : std_logic;
signal \N__61118\ : std_logic;
signal \N__61117\ : std_logic;
signal \N__61112\ : std_logic;
signal \N__61109\ : std_logic;
signal \N__61106\ : std_logic;
signal \N__61103\ : std_logic;
signal \N__61100\ : std_logic;
signal \N__61099\ : std_logic;
signal \N__61096\ : std_logic;
signal \N__61093\ : std_logic;
signal \N__61092\ : std_logic;
signal \N__61087\ : std_logic;
signal \N__61082\ : std_logic;
signal \N__61081\ : std_logic;
signal \N__61080\ : std_logic;
signal \N__61079\ : std_logic;
signal \N__61078\ : std_logic;
signal \N__61077\ : std_logic;
signal \N__61074\ : std_logic;
signal \N__61073\ : std_logic;
signal \N__61070\ : std_logic;
signal \N__61067\ : std_logic;
signal \N__61064\ : std_logic;
signal \N__61061\ : std_logic;
signal \N__61058\ : std_logic;
signal \N__61055\ : std_logic;
signal \N__61048\ : std_logic;
signal \N__61045\ : std_logic;
signal \N__61040\ : std_logic;
signal \N__61033\ : std_logic;
signal \N__61018\ : std_logic;
signal \N__61015\ : std_logic;
signal \N__61012\ : std_logic;
signal \N__61011\ : std_logic;
signal \N__61008\ : std_logic;
signal \N__61005\ : std_logic;
signal \N__61002\ : std_logic;
signal \N__60999\ : std_logic;
signal \N__60994\ : std_logic;
signal \N__60991\ : std_logic;
signal \N__60988\ : std_logic;
signal \N__60987\ : std_logic;
signal \N__60984\ : std_logic;
signal \N__60983\ : std_logic;
signal \N__60980\ : std_logic;
signal \N__60977\ : std_logic;
signal \N__60976\ : std_logic;
signal \N__60973\ : std_logic;
signal \N__60970\ : std_logic;
signal \N__60967\ : std_logic;
signal \N__60964\ : std_logic;
signal \N__60961\ : std_logic;
signal \N__60958\ : std_logic;
signal \N__60957\ : std_logic;
signal \N__60956\ : std_logic;
signal \N__60953\ : std_logic;
signal \N__60950\ : std_logic;
signal \N__60945\ : std_logic;
signal \N__60940\ : std_logic;
signal \N__60931\ : std_logic;
signal \N__60928\ : std_logic;
signal \N__60927\ : std_logic;
signal \N__60926\ : std_logic;
signal \N__60923\ : std_logic;
signal \N__60922\ : std_logic;
signal \N__60917\ : std_logic;
signal \N__60916\ : std_logic;
signal \N__60913\ : std_logic;
signal \N__60910\ : std_logic;
signal \N__60909\ : std_logic;
signal \N__60908\ : std_logic;
signal \N__60907\ : std_logic;
signal \N__60906\ : std_logic;
signal \N__60905\ : std_logic;
signal \N__60902\ : std_logic;
signal \N__60901\ : std_logic;
signal \N__60900\ : std_logic;
signal \N__60899\ : std_logic;
signal \N__60896\ : std_logic;
signal \N__60893\ : std_logic;
signal \N__60890\ : std_logic;
signal \N__60887\ : std_logic;
signal \N__60884\ : std_logic;
signal \N__60881\ : std_logic;
signal \N__60876\ : std_logic;
signal \N__60873\ : std_logic;
signal \N__60868\ : std_logic;
signal \N__60865\ : std_logic;
signal \N__60844\ : std_logic;
signal \N__60843\ : std_logic;
signal \N__60842\ : std_logic;
signal \N__60839\ : std_logic;
signal \N__60836\ : std_logic;
signal \N__60833\ : std_logic;
signal \N__60830\ : std_logic;
signal \N__60829\ : std_logic;
signal \N__60826\ : std_logic;
signal \N__60823\ : std_logic;
signal \N__60820\ : std_logic;
signal \N__60817\ : std_logic;
signal \N__60814\ : std_logic;
signal \N__60811\ : std_logic;
signal \N__60808\ : std_logic;
signal \N__60805\ : std_logic;
signal \N__60802\ : std_logic;
signal \N__60793\ : std_logic;
signal \N__60792\ : std_logic;
signal \N__60791\ : std_logic;
signal \N__60788\ : std_logic;
signal \N__60785\ : std_logic;
signal \N__60782\ : std_logic;
signal \N__60779\ : std_logic;
signal \N__60778\ : std_logic;
signal \N__60775\ : std_logic;
signal \N__60772\ : std_logic;
signal \N__60771\ : std_logic;
signal \N__60768\ : std_logic;
signal \N__60765\ : std_logic;
signal \N__60762\ : std_logic;
signal \N__60759\ : std_logic;
signal \N__60756\ : std_logic;
signal \N__60745\ : std_logic;
signal \N__60742\ : std_logic;
signal \N__60739\ : std_logic;
signal \N__60736\ : std_logic;
signal \N__60733\ : std_logic;
signal \N__60730\ : std_logic;
signal \N__60729\ : std_logic;
signal \N__60726\ : std_logic;
signal \N__60723\ : std_logic;
signal \N__60718\ : std_logic;
signal \N__60717\ : std_logic;
signal \N__60714\ : std_logic;
signal \N__60711\ : std_logic;
signal \N__60710\ : std_logic;
signal \N__60709\ : std_logic;
signal \N__60704\ : std_logic;
signal \N__60699\ : std_logic;
signal \N__60696\ : std_logic;
signal \N__60695\ : std_logic;
signal \N__60694\ : std_logic;
signal \N__60693\ : std_logic;
signal \N__60692\ : std_logic;
signal \N__60691\ : std_logic;
signal \N__60690\ : std_logic;
signal \N__60689\ : std_logic;
signal \N__60688\ : std_logic;
signal \N__60687\ : std_logic;
signal \N__60686\ : std_logic;
signal \N__60683\ : std_logic;
signal \N__60680\ : std_logic;
signal \N__60677\ : std_logic;
signal \N__60668\ : std_logic;
signal \N__60663\ : std_logic;
signal \N__60660\ : std_logic;
signal \N__60655\ : std_logic;
signal \N__60654\ : std_logic;
signal \N__60653\ : std_logic;
signal \N__60652\ : std_logic;
signal \N__60651\ : std_logic;
signal \N__60650\ : std_logic;
signal \N__60647\ : std_logic;
signal \N__60644\ : std_logic;
signal \N__60641\ : std_logic;
signal \N__60636\ : std_logic;
signal \N__60635\ : std_logic;
signal \N__60634\ : std_logic;
signal \N__60633\ : std_logic;
signal \N__60632\ : std_logic;
signal \N__60629\ : std_logic;
signal \N__60626\ : std_logic;
signal \N__60621\ : std_logic;
signal \N__60620\ : std_logic;
signal \N__60619\ : std_logic;
signal \N__60618\ : std_logic;
signal \N__60617\ : std_logic;
signal \N__60612\ : std_logic;
signal \N__60609\ : std_logic;
signal \N__60606\ : std_logic;
signal \N__60603\ : std_logic;
signal \N__60600\ : std_logic;
signal \N__60597\ : std_logic;
signal \N__60592\ : std_logic;
signal \N__60589\ : std_logic;
signal \N__60586\ : std_logic;
signal \N__60585\ : std_logic;
signal \N__60584\ : std_logic;
signal \N__60583\ : std_logic;
signal \N__60576\ : std_logic;
signal \N__60567\ : std_logic;
signal \N__60560\ : std_logic;
signal \N__60555\ : std_logic;
signal \N__60552\ : std_logic;
signal \N__60549\ : std_logic;
signal \N__60546\ : std_logic;
signal \N__60543\ : std_logic;
signal \N__60538\ : std_logic;
signal \N__60535\ : std_logic;
signal \N__60528\ : std_logic;
signal \N__60511\ : std_logic;
signal \N__60508\ : std_logic;
signal \N__60505\ : std_logic;
signal \N__60502\ : std_logic;
signal \N__60499\ : std_logic;
signal \N__60496\ : std_logic;
signal \N__60493\ : std_logic;
signal \N__60492\ : std_logic;
signal \N__60489\ : std_logic;
signal \N__60488\ : std_logic;
signal \N__60487\ : std_logic;
signal \N__60482\ : std_logic;
signal \N__60479\ : std_logic;
signal \N__60478\ : std_logic;
signal \N__60475\ : std_logic;
signal \N__60472\ : std_logic;
signal \N__60469\ : std_logic;
signal \N__60466\ : std_logic;
signal \N__60461\ : std_logic;
signal \N__60458\ : std_logic;
signal \N__60451\ : std_logic;
signal \N__60450\ : std_logic;
signal \N__60449\ : std_logic;
signal \N__60448\ : std_logic;
signal \N__60445\ : std_logic;
signal \N__60442\ : std_logic;
signal \N__60439\ : std_logic;
signal \N__60436\ : std_logic;
signal \N__60433\ : std_logic;
signal \N__60430\ : std_logic;
signal \N__60427\ : std_logic;
signal \N__60422\ : std_logic;
signal \N__60419\ : std_logic;
signal \N__60412\ : std_logic;
signal \N__60411\ : std_logic;
signal \N__60408\ : std_logic;
signal \N__60405\ : std_logic;
signal \N__60402\ : std_logic;
signal \N__60399\ : std_logic;
signal \N__60398\ : std_logic;
signal \N__60395\ : std_logic;
signal \N__60392\ : std_logic;
signal \N__60391\ : std_logic;
signal \N__60390\ : std_logic;
signal \N__60389\ : std_logic;
signal \N__60388\ : std_logic;
signal \N__60385\ : std_logic;
signal \N__60382\ : std_logic;
signal \N__60379\ : std_logic;
signal \N__60372\ : std_logic;
signal \N__60369\ : std_logic;
signal \N__60358\ : std_logic;
signal \N__60355\ : std_logic;
signal \N__60354\ : std_logic;
signal \N__60353\ : std_logic;
signal \N__60352\ : std_logic;
signal \N__60347\ : std_logic;
signal \N__60346\ : std_logic;
signal \N__60343\ : std_logic;
signal \N__60340\ : std_logic;
signal \N__60337\ : std_logic;
signal \N__60336\ : std_logic;
signal \N__60333\ : std_logic;
signal \N__60330\ : std_logic;
signal \N__60329\ : std_logic;
signal \N__60326\ : std_logic;
signal \N__60323\ : std_logic;
signal \N__60320\ : std_logic;
signal \N__60319\ : std_logic;
signal \N__60316\ : std_logic;
signal \N__60313\ : std_logic;
signal \N__60310\ : std_logic;
signal \N__60309\ : std_logic;
signal \N__60302\ : std_logic;
signal \N__60299\ : std_logic;
signal \N__60296\ : std_logic;
signal \N__60293\ : std_logic;
signal \N__60288\ : std_logic;
signal \N__60281\ : std_logic;
signal \N__60274\ : std_logic;
signal \N__60273\ : std_logic;
signal \N__60272\ : std_logic;
signal \N__60269\ : std_logic;
signal \N__60268\ : std_logic;
signal \N__60265\ : std_logic;
signal \N__60264\ : std_logic;
signal \N__60263\ : std_logic;
signal \N__60260\ : std_logic;
signal \N__60257\ : std_logic;
signal \N__60256\ : std_logic;
signal \N__60253\ : std_logic;
signal \N__60252\ : std_logic;
signal \N__60249\ : std_logic;
signal \N__60246\ : std_logic;
signal \N__60243\ : std_logic;
signal \N__60242\ : std_logic;
signal \N__60239\ : std_logic;
signal \N__60236\ : std_logic;
signal \N__60235\ : std_logic;
signal \N__60232\ : std_logic;
signal \N__60229\ : std_logic;
signal \N__60226\ : std_logic;
signal \N__60223\ : std_logic;
signal \N__60220\ : std_logic;
signal \N__60215\ : std_logic;
signal \N__60212\ : std_logic;
signal \N__60209\ : std_logic;
signal \N__60208\ : std_logic;
signal \N__60205\ : std_logic;
signal \N__60204\ : std_logic;
signal \N__60201\ : std_logic;
signal \N__60198\ : std_logic;
signal \N__60195\ : std_logic;
signal \N__60192\ : std_logic;
signal \N__60189\ : std_logic;
signal \N__60186\ : std_logic;
signal \N__60183\ : std_logic;
signal \N__60180\ : std_logic;
signal \N__60177\ : std_logic;
signal \N__60174\ : std_logic;
signal \N__60171\ : std_logic;
signal \N__60168\ : std_logic;
signal \N__60163\ : std_logic;
signal \N__60154\ : std_logic;
signal \N__60151\ : std_logic;
signal \N__60148\ : std_logic;
signal \N__60133\ : std_logic;
signal \N__60132\ : std_logic;
signal \N__60129\ : std_logic;
signal \N__60128\ : std_logic;
signal \N__60125\ : std_logic;
signal \N__60122\ : std_logic;
signal \N__60121\ : std_logic;
signal \N__60118\ : std_logic;
signal \N__60117\ : std_logic;
signal \N__60116\ : std_logic;
signal \N__60115\ : std_logic;
signal \N__60112\ : std_logic;
signal \N__60109\ : std_logic;
signal \N__60108\ : std_logic;
signal \N__60105\ : std_logic;
signal \N__60104\ : std_logic;
signal \N__60101\ : std_logic;
signal \N__60098\ : std_logic;
signal \N__60095\ : std_logic;
signal \N__60092\ : std_logic;
signal \N__60089\ : std_logic;
signal \N__60086\ : std_logic;
signal \N__60083\ : std_logic;
signal \N__60080\ : std_logic;
signal \N__60077\ : std_logic;
signal \N__60072\ : std_logic;
signal \N__60069\ : std_logic;
signal \N__60064\ : std_logic;
signal \N__60061\ : std_logic;
signal \N__60058\ : std_logic;
signal \N__60053\ : std_logic;
signal \N__60050\ : std_logic;
signal \N__60049\ : std_logic;
signal \N__60048\ : std_logic;
signal \N__60047\ : std_logic;
signal \N__60042\ : std_logic;
signal \N__60041\ : std_logic;
signal \N__60038\ : std_logic;
signal \N__60035\ : std_logic;
signal \N__60032\ : std_logic;
signal \N__60029\ : std_logic;
signal \N__60022\ : std_logic;
signal \N__60019\ : std_logic;
signal \N__60016\ : std_logic;
signal \N__60001\ : std_logic;
signal \N__60000\ : std_logic;
signal \N__59997\ : std_logic;
signal \N__59996\ : std_logic;
signal \N__59993\ : std_logic;
signal \N__59992\ : std_logic;
signal \N__59989\ : std_logic;
signal \N__59986\ : std_logic;
signal \N__59985\ : std_logic;
signal \N__59982\ : std_logic;
signal \N__59979\ : std_logic;
signal \N__59978\ : std_logic;
signal \N__59977\ : std_logic;
signal \N__59972\ : std_logic;
signal \N__59969\ : std_logic;
signal \N__59966\ : std_logic;
signal \N__59965\ : std_logic;
signal \N__59962\ : std_logic;
signal \N__59959\ : std_logic;
signal \N__59956\ : std_logic;
signal \N__59951\ : std_logic;
signal \N__59948\ : std_logic;
signal \N__59945\ : std_logic;
signal \N__59944\ : std_logic;
signal \N__59939\ : std_logic;
signal \N__59934\ : std_logic;
signal \N__59931\ : std_logic;
signal \N__59928\ : std_logic;
signal \N__59927\ : std_logic;
signal \N__59924\ : std_logic;
signal \N__59923\ : std_logic;
signal \N__59922\ : std_logic;
signal \N__59921\ : std_logic;
signal \N__59914\ : std_logic;
signal \N__59911\ : std_logic;
signal \N__59908\ : std_logic;
signal \N__59899\ : std_logic;
signal \N__59896\ : std_logic;
signal \N__59893\ : std_logic;
signal \N__59884\ : std_logic;
signal \N__59883\ : std_logic;
signal \N__59880\ : std_logic;
signal \N__59877\ : std_logic;
signal \N__59876\ : std_logic;
signal \N__59875\ : std_logic;
signal \N__59870\ : std_logic;
signal \N__59869\ : std_logic;
signal \N__59868\ : std_logic;
signal \N__59867\ : std_logic;
signal \N__59866\ : std_logic;
signal \N__59861\ : std_logic;
signal \N__59858\ : std_logic;
signal \N__59855\ : std_logic;
signal \N__59848\ : std_logic;
signal \N__59845\ : std_logic;
signal \N__59842\ : std_logic;
signal \N__59833\ : std_logic;
signal \N__59832\ : std_logic;
signal \N__59829\ : std_logic;
signal \N__59828\ : std_logic;
signal \N__59825\ : std_logic;
signal \N__59822\ : std_logic;
signal \N__59819\ : std_logic;
signal \N__59812\ : std_logic;
signal \N__59809\ : std_logic;
signal \N__59806\ : std_logic;
signal \N__59803\ : std_logic;
signal \N__59800\ : std_logic;
signal \N__59797\ : std_logic;
signal \N__59794\ : std_logic;
signal \N__59791\ : std_logic;
signal \N__59788\ : std_logic;
signal \N__59785\ : std_logic;
signal \N__59784\ : std_logic;
signal \N__59783\ : std_logic;
signal \N__59780\ : std_logic;
signal \N__59779\ : std_logic;
signal \N__59776\ : std_logic;
signal \N__59775\ : std_logic;
signal \N__59772\ : std_logic;
signal \N__59769\ : std_logic;
signal \N__59766\ : std_logic;
signal \N__59763\ : std_logic;
signal \N__59760\ : std_logic;
signal \N__59757\ : std_logic;
signal \N__59748\ : std_logic;
signal \N__59743\ : std_logic;
signal \N__59742\ : std_logic;
signal \N__59739\ : std_logic;
signal \N__59738\ : std_logic;
signal \N__59735\ : std_logic;
signal \N__59732\ : std_logic;
signal \N__59729\ : std_logic;
signal \N__59726\ : std_logic;
signal \N__59723\ : std_logic;
signal \N__59720\ : std_logic;
signal \N__59719\ : std_logic;
signal \N__59712\ : std_logic;
signal \N__59709\ : std_logic;
signal \N__59706\ : std_logic;
signal \N__59701\ : std_logic;
signal \N__59700\ : std_logic;
signal \N__59699\ : std_logic;
signal \N__59696\ : std_logic;
signal \N__59693\ : std_logic;
signal \N__59692\ : std_logic;
signal \N__59689\ : std_logic;
signal \N__59688\ : std_logic;
signal \N__59685\ : std_logic;
signal \N__59682\ : std_logic;
signal \N__59679\ : std_logic;
signal \N__59676\ : std_logic;
signal \N__59673\ : std_logic;
signal \N__59670\ : std_logic;
signal \N__59669\ : std_logic;
signal \N__59666\ : std_logic;
signal \N__59663\ : std_logic;
signal \N__59660\ : std_logic;
signal \N__59657\ : std_logic;
signal \N__59654\ : std_logic;
signal \N__59651\ : std_logic;
signal \N__59644\ : std_logic;
signal \N__59639\ : std_logic;
signal \N__59636\ : std_logic;
signal \N__59633\ : std_logic;
signal \N__59630\ : std_logic;
signal \N__59623\ : std_logic;
signal \N__59620\ : std_logic;
signal \N__59617\ : std_logic;
signal \N__59616\ : std_logic;
signal \N__59613\ : std_logic;
signal \N__59612\ : std_logic;
signal \N__59609\ : std_logic;
signal \N__59606\ : std_logic;
signal \N__59603\ : std_logic;
signal \N__59596\ : std_logic;
signal \N__59595\ : std_logic;
signal \N__59592\ : std_logic;
signal \N__59589\ : std_logic;
signal \N__59588\ : std_logic;
signal \N__59585\ : std_logic;
signal \N__59582\ : std_logic;
signal \N__59579\ : std_logic;
signal \N__59576\ : std_logic;
signal \N__59571\ : std_logic;
signal \N__59568\ : std_logic;
signal \N__59565\ : std_logic;
signal \N__59560\ : std_logic;
signal \N__59557\ : std_logic;
signal \N__59556\ : std_logic;
signal \N__59553\ : std_logic;
signal \N__59550\ : std_logic;
signal \N__59549\ : std_logic;
signal \N__59548\ : std_logic;
signal \N__59545\ : std_logic;
signal \N__59540\ : std_logic;
signal \N__59537\ : std_logic;
signal \N__59530\ : std_logic;
signal \N__59527\ : std_logic;
signal \N__59524\ : std_logic;
signal \N__59521\ : std_logic;
signal \N__59518\ : std_logic;
signal \N__59515\ : std_logic;
signal \N__59512\ : std_logic;
signal \N__59511\ : std_logic;
signal \N__59508\ : std_logic;
signal \N__59505\ : std_logic;
signal \N__59504\ : std_logic;
signal \N__59501\ : std_logic;
signal \N__59498\ : std_logic;
signal \N__59495\ : std_logic;
signal \N__59488\ : std_logic;
signal \N__59485\ : std_logic;
signal \N__59482\ : std_logic;
signal \N__59481\ : std_logic;
signal \N__59480\ : std_logic;
signal \N__59479\ : std_logic;
signal \N__59478\ : std_logic;
signal \N__59475\ : std_logic;
signal \N__59472\ : std_logic;
signal \N__59469\ : std_logic;
signal \N__59466\ : std_logic;
signal \N__59463\ : std_logic;
signal \N__59460\ : std_logic;
signal \N__59459\ : std_logic;
signal \N__59456\ : std_logic;
signal \N__59455\ : std_logic;
signal \N__59452\ : std_logic;
signal \N__59449\ : std_logic;
signal \N__59448\ : std_logic;
signal \N__59443\ : std_logic;
signal \N__59440\ : std_logic;
signal \N__59439\ : std_logic;
signal \N__59436\ : std_logic;
signal \N__59433\ : std_logic;
signal \N__59432\ : std_logic;
signal \N__59429\ : std_logic;
signal \N__59426\ : std_logic;
signal \N__59423\ : std_logic;
signal \N__59418\ : std_logic;
signal \N__59415\ : std_logic;
signal \N__59412\ : std_logic;
signal \N__59409\ : std_logic;
signal \N__59406\ : std_logic;
signal \N__59403\ : std_logic;
signal \N__59396\ : std_logic;
signal \N__59393\ : std_logic;
signal \N__59380\ : std_logic;
signal \N__59377\ : std_logic;
signal \N__59374\ : std_logic;
signal \N__59371\ : std_logic;
signal \N__59368\ : std_logic;
signal \N__59365\ : std_logic;
signal \N__59362\ : std_logic;
signal \N__59359\ : std_logic;
signal \N__59358\ : std_logic;
signal \N__59355\ : std_logic;
signal \N__59352\ : std_logic;
signal \N__59349\ : std_logic;
signal \N__59346\ : std_logic;
signal \N__59345\ : std_logic;
signal \N__59340\ : std_logic;
signal \N__59337\ : std_logic;
signal \N__59332\ : std_logic;
signal \N__59329\ : std_logic;
signal \N__59326\ : std_logic;
signal \N__59325\ : std_logic;
signal \N__59324\ : std_logic;
signal \N__59321\ : std_logic;
signal \N__59318\ : std_logic;
signal \N__59315\ : std_logic;
signal \N__59312\ : std_logic;
signal \N__59307\ : std_logic;
signal \N__59302\ : std_logic;
signal \N__59301\ : std_logic;
signal \N__59300\ : std_logic;
signal \N__59297\ : std_logic;
signal \N__59294\ : std_logic;
signal \N__59291\ : std_logic;
signal \N__59288\ : std_logic;
signal \N__59285\ : std_logic;
signal \N__59282\ : std_logic;
signal \N__59279\ : std_logic;
signal \N__59276\ : std_logic;
signal \N__59275\ : std_logic;
signal \N__59274\ : std_logic;
signal \N__59269\ : std_logic;
signal \N__59266\ : std_logic;
signal \N__59261\ : std_logic;
signal \N__59254\ : std_logic;
signal \N__59251\ : std_logic;
signal \N__59250\ : std_logic;
signal \N__59247\ : std_logic;
signal \N__59244\ : std_logic;
signal \N__59241\ : std_logic;
signal \N__59238\ : std_logic;
signal \N__59237\ : std_logic;
signal \N__59232\ : std_logic;
signal \N__59231\ : std_logic;
signal \N__59230\ : std_logic;
signal \N__59227\ : std_logic;
signal \N__59224\ : std_logic;
signal \N__59219\ : std_logic;
signal \N__59212\ : std_logic;
signal \N__59211\ : std_logic;
signal \N__59208\ : std_logic;
signal \N__59205\ : std_logic;
signal \N__59202\ : std_logic;
signal \N__59199\ : std_logic;
signal \N__59196\ : std_logic;
signal \N__59191\ : std_logic;
signal \N__59190\ : std_logic;
signal \N__59187\ : std_logic;
signal \N__59184\ : std_logic;
signal \N__59179\ : std_logic;
signal \N__59178\ : std_logic;
signal \N__59175\ : std_logic;
signal \N__59172\ : std_logic;
signal \N__59169\ : std_logic;
signal \N__59166\ : std_logic;
signal \N__59165\ : std_logic;
signal \N__59162\ : std_logic;
signal \N__59159\ : std_logic;
signal \N__59156\ : std_logic;
signal \N__59149\ : std_logic;
signal \N__59146\ : std_logic;
signal \N__59143\ : std_logic;
signal \N__59140\ : std_logic;
signal \N__59137\ : std_logic;
signal \N__59134\ : std_logic;
signal \N__59133\ : std_logic;
signal \N__59130\ : std_logic;
signal \N__59127\ : std_logic;
signal \N__59126\ : std_logic;
signal \N__59123\ : std_logic;
signal \N__59120\ : std_logic;
signal \N__59117\ : std_logic;
signal \N__59116\ : std_logic;
signal \N__59115\ : std_logic;
signal \N__59112\ : std_logic;
signal \N__59107\ : std_logic;
signal \N__59104\ : std_logic;
signal \N__59101\ : std_logic;
signal \N__59098\ : std_logic;
signal \N__59095\ : std_logic;
signal \N__59086\ : std_logic;
signal \N__59085\ : std_logic;
signal \N__59082\ : std_logic;
signal \N__59079\ : std_logic;
signal \N__59076\ : std_logic;
signal \N__59075\ : std_logic;
signal \N__59074\ : std_logic;
signal \N__59073\ : std_logic;
signal \N__59072\ : std_logic;
signal \N__59069\ : std_logic;
signal \N__59066\ : std_logic;
signal \N__59061\ : std_logic;
signal \N__59056\ : std_logic;
signal \N__59047\ : std_logic;
signal \N__59046\ : std_logic;
signal \N__59043\ : std_logic;
signal \N__59040\ : std_logic;
signal \N__59039\ : std_logic;
signal \N__59036\ : std_logic;
signal \N__59033\ : std_logic;
signal \N__59032\ : std_logic;
signal \N__59029\ : std_logic;
signal \N__59024\ : std_logic;
signal \N__59021\ : std_logic;
signal \N__59014\ : std_logic;
signal \N__59011\ : std_logic;
signal \N__59010\ : std_logic;
signal \N__59009\ : std_logic;
signal \N__59006\ : std_logic;
signal \N__59005\ : std_logic;
signal \N__59004\ : std_logic;
signal \N__59003\ : std_logic;
signal \N__59002\ : std_logic;
signal \N__58999\ : std_logic;
signal \N__58998\ : std_logic;
signal \N__58995\ : std_logic;
signal \N__58992\ : std_logic;
signal \N__58985\ : std_logic;
signal \N__58982\ : std_logic;
signal \N__58979\ : std_logic;
signal \N__58976\ : std_logic;
signal \N__58967\ : std_logic;
signal \N__58962\ : std_logic;
signal \N__58959\ : std_logic;
signal \N__58954\ : std_logic;
signal \N__58951\ : std_logic;
signal \N__58948\ : std_logic;
signal \N__58945\ : std_logic;
signal \N__58942\ : std_logic;
signal \N__58941\ : std_logic;
signal \N__58940\ : std_logic;
signal \N__58937\ : std_logic;
signal \N__58932\ : std_logic;
signal \N__58931\ : std_logic;
signal \N__58926\ : std_logic;
signal \N__58923\ : std_logic;
signal \N__58920\ : std_logic;
signal \N__58917\ : std_logic;
signal \N__58912\ : std_logic;
signal \N__58909\ : std_logic;
signal \N__58906\ : std_logic;
signal \N__58903\ : std_logic;
signal \N__58900\ : std_logic;
signal \N__58899\ : std_logic;
signal \N__58896\ : std_logic;
signal \N__58895\ : std_logic;
signal \N__58892\ : std_logic;
signal \N__58889\ : std_logic;
signal \N__58886\ : std_logic;
signal \N__58883\ : std_logic;
signal \N__58878\ : std_logic;
signal \N__58875\ : std_logic;
signal \N__58872\ : std_logic;
signal \N__58871\ : std_logic;
signal \N__58868\ : std_logic;
signal \N__58865\ : std_logic;
signal \N__58862\ : std_logic;
signal \N__58859\ : std_logic;
signal \N__58856\ : std_logic;
signal \N__58849\ : std_logic;
signal \N__58846\ : std_logic;
signal \N__58843\ : std_logic;
signal \N__58840\ : std_logic;
signal \N__58839\ : std_logic;
signal \N__58836\ : std_logic;
signal \N__58833\ : std_logic;
signal \N__58832\ : std_logic;
signal \N__58829\ : std_logic;
signal \N__58826\ : std_logic;
signal \N__58823\ : std_logic;
signal \N__58822\ : std_logic;
signal \N__58819\ : std_logic;
signal \N__58814\ : std_logic;
signal \N__58811\ : std_logic;
signal \N__58808\ : std_logic;
signal \N__58805\ : std_logic;
signal \N__58798\ : std_logic;
signal \N__58795\ : std_logic;
signal \N__58794\ : std_logic;
signal \N__58791\ : std_logic;
signal \N__58790\ : std_logic;
signal \N__58787\ : std_logic;
signal \N__58784\ : std_logic;
signal \N__58781\ : std_logic;
signal \N__58778\ : std_logic;
signal \N__58775\ : std_logic;
signal \N__58768\ : std_logic;
signal \N__58765\ : std_logic;
signal \N__58762\ : std_logic;
signal \N__58761\ : std_logic;
signal \N__58760\ : std_logic;
signal \N__58757\ : std_logic;
signal \N__58756\ : std_logic;
signal \N__58753\ : std_logic;
signal \N__58750\ : std_logic;
signal \N__58747\ : std_logic;
signal \N__58744\ : std_logic;
signal \N__58741\ : std_logic;
signal \N__58738\ : std_logic;
signal \N__58735\ : std_logic;
signal \N__58726\ : std_logic;
signal \N__58725\ : std_logic;
signal \N__58724\ : std_logic;
signal \N__58719\ : std_logic;
signal \N__58716\ : std_logic;
signal \N__58715\ : std_logic;
signal \N__58712\ : std_logic;
signal \N__58709\ : std_logic;
signal \N__58708\ : std_logic;
signal \N__58705\ : std_logic;
signal \N__58700\ : std_logic;
signal \N__58697\ : std_logic;
signal \N__58694\ : std_logic;
signal \N__58691\ : std_logic;
signal \N__58688\ : std_logic;
signal \N__58685\ : std_logic;
signal \N__58682\ : std_logic;
signal \N__58675\ : std_logic;
signal \N__58672\ : std_logic;
signal \N__58669\ : std_logic;
signal \N__58668\ : std_logic;
signal \N__58667\ : std_logic;
signal \N__58664\ : std_logic;
signal \N__58661\ : std_logic;
signal \N__58658\ : std_logic;
signal \N__58655\ : std_logic;
signal \N__58650\ : std_logic;
signal \N__58649\ : std_logic;
signal \N__58646\ : std_logic;
signal \N__58643\ : std_logic;
signal \N__58640\ : std_logic;
signal \N__58633\ : std_logic;
signal \N__58630\ : std_logic;
signal \N__58629\ : std_logic;
signal \N__58626\ : std_logic;
signal \N__58623\ : std_logic;
signal \N__58620\ : std_logic;
signal \N__58617\ : std_logic;
signal \N__58612\ : std_logic;
signal \N__58609\ : std_logic;
signal \N__58606\ : std_logic;
signal \N__58603\ : std_logic;
signal \N__58600\ : std_logic;
signal \N__58599\ : std_logic;
signal \N__58598\ : std_logic;
signal \N__58595\ : std_logic;
signal \N__58592\ : std_logic;
signal \N__58589\ : std_logic;
signal \N__58582\ : std_logic;
signal \N__58579\ : std_logic;
signal \N__58576\ : std_logic;
signal \N__58573\ : std_logic;
signal \N__58570\ : std_logic;
signal \N__58567\ : std_logic;
signal \N__58564\ : std_logic;
signal \N__58561\ : std_logic;
signal \N__58558\ : std_logic;
signal \N__58555\ : std_logic;
signal \N__58552\ : std_logic;
signal \N__58551\ : std_logic;
signal \N__58550\ : std_logic;
signal \N__58547\ : std_logic;
signal \N__58544\ : std_logic;
signal \N__58541\ : std_logic;
signal \N__58538\ : std_logic;
signal \N__58535\ : std_logic;
signal \N__58532\ : std_logic;
signal \N__58529\ : std_logic;
signal \N__58526\ : std_logic;
signal \N__58523\ : std_logic;
signal \N__58518\ : std_logic;
signal \N__58515\ : std_logic;
signal \N__58510\ : std_logic;
signal \N__58507\ : std_logic;
signal \N__58506\ : std_logic;
signal \N__58503\ : std_logic;
signal \N__58500\ : std_logic;
signal \N__58495\ : std_logic;
signal \N__58492\ : std_logic;
signal \N__58491\ : std_logic;
signal \N__58488\ : std_logic;
signal \N__58485\ : std_logic;
signal \N__58482\ : std_logic;
signal \N__58479\ : std_logic;
signal \N__58476\ : std_logic;
signal \N__58473\ : std_logic;
signal \N__58468\ : std_logic;
signal \N__58467\ : std_logic;
signal \N__58466\ : std_logic;
signal \N__58463\ : std_logic;
signal \N__58462\ : std_logic;
signal \N__58461\ : std_logic;
signal \N__58458\ : std_logic;
signal \N__58455\ : std_logic;
signal \N__58452\ : std_logic;
signal \N__58449\ : std_logic;
signal \N__58446\ : std_logic;
signal \N__58443\ : std_logic;
signal \N__58440\ : std_logic;
signal \N__58433\ : std_logic;
signal \N__58432\ : std_logic;
signal \N__58431\ : std_logic;
signal \N__58428\ : std_logic;
signal \N__58423\ : std_logic;
signal \N__58420\ : std_logic;
signal \N__58417\ : std_logic;
signal \N__58408\ : std_logic;
signal \N__58405\ : std_logic;
signal \N__58404\ : std_logic;
signal \N__58401\ : std_logic;
signal \N__58398\ : std_logic;
signal \N__58395\ : std_logic;
signal \N__58392\ : std_logic;
signal \N__58387\ : std_logic;
signal \N__58384\ : std_logic;
signal \N__58381\ : std_logic;
signal \N__58378\ : std_logic;
signal \N__58375\ : std_logic;
signal \N__58372\ : std_logic;
signal \N__58369\ : std_logic;
signal \N__58368\ : std_logic;
signal \N__58365\ : std_logic;
signal \N__58362\ : std_logic;
signal \N__58359\ : std_logic;
signal \N__58354\ : std_logic;
signal \N__58353\ : std_logic;
signal \N__58350\ : std_logic;
signal \N__58347\ : std_logic;
signal \N__58342\ : std_logic;
signal \N__58339\ : std_logic;
signal \N__58336\ : std_logic;
signal \N__58335\ : std_logic;
signal \N__58330\ : std_logic;
signal \N__58327\ : std_logic;
signal \N__58324\ : std_logic;
signal \N__58321\ : std_logic;
signal \N__58318\ : std_logic;
signal \N__58315\ : std_logic;
signal \N__58312\ : std_logic;
signal \N__58309\ : std_logic;
signal \N__58306\ : std_logic;
signal \N__58305\ : std_logic;
signal \N__58300\ : std_logic;
signal \N__58297\ : std_logic;
signal \N__58294\ : std_logic;
signal \N__58291\ : std_logic;
signal \N__58288\ : std_logic;
signal \N__58287\ : std_logic;
signal \N__58284\ : std_logic;
signal \N__58281\ : std_logic;
signal \N__58276\ : std_logic;
signal \N__58273\ : std_logic;
signal \N__58270\ : std_logic;
signal \N__58267\ : std_logic;
signal \N__58264\ : std_logic;
signal \N__58261\ : std_logic;
signal \N__58258\ : std_logic;
signal \N__58255\ : std_logic;
signal \N__58252\ : std_logic;
signal \N__58249\ : std_logic;
signal \N__58248\ : std_logic;
signal \N__58247\ : std_logic;
signal \N__58244\ : std_logic;
signal \N__58239\ : std_logic;
signal \N__58236\ : std_logic;
signal \N__58233\ : std_logic;
signal \N__58228\ : std_logic;
signal \N__58227\ : std_logic;
signal \N__58224\ : std_logic;
signal \N__58221\ : std_logic;
signal \N__58218\ : std_logic;
signal \N__58217\ : std_logic;
signal \N__58212\ : std_logic;
signal \N__58209\ : std_logic;
signal \N__58204\ : std_logic;
signal \N__58201\ : std_logic;
signal \N__58200\ : std_logic;
signal \N__58199\ : std_logic;
signal \N__58194\ : std_logic;
signal \N__58191\ : std_logic;
signal \N__58186\ : std_logic;
signal \N__58183\ : std_logic;
signal \N__58180\ : std_logic;
signal \N__58177\ : std_logic;
signal \N__58174\ : std_logic;
signal \N__58171\ : std_logic;
signal \N__58168\ : std_logic;
signal \N__58165\ : std_logic;
signal \N__58162\ : std_logic;
signal \N__58159\ : std_logic;
signal \N__58156\ : std_logic;
signal \N__58153\ : std_logic;
signal \N__58150\ : std_logic;
signal \N__58147\ : std_logic;
signal \N__58144\ : std_logic;
signal \N__58141\ : std_logic;
signal \N__58138\ : std_logic;
signal \N__58135\ : std_logic;
signal \N__58132\ : std_logic;
signal \N__58131\ : std_logic;
signal \N__58130\ : std_logic;
signal \N__58127\ : std_logic;
signal \N__58124\ : std_logic;
signal \N__58121\ : std_logic;
signal \N__58114\ : std_logic;
signal \N__58111\ : std_logic;
signal \N__58108\ : std_logic;
signal \N__58105\ : std_logic;
signal \N__58102\ : std_logic;
signal \N__58099\ : std_logic;
signal \N__58098\ : std_logic;
signal \N__58097\ : std_logic;
signal \N__58094\ : std_logic;
signal \N__58089\ : std_logic;
signal \N__58084\ : std_logic;
signal \N__58081\ : std_logic;
signal \N__58078\ : std_logic;
signal \N__58075\ : std_logic;
signal \N__58072\ : std_logic;
signal \N__58069\ : std_logic;
signal \N__58068\ : std_logic;
signal \N__58067\ : std_logic;
signal \N__58064\ : std_logic;
signal \N__58059\ : std_logic;
signal \N__58054\ : std_logic;
signal \N__58053\ : std_logic;
signal \N__58050\ : std_logic;
signal \N__58047\ : std_logic;
signal \N__58042\ : std_logic;
signal \N__58041\ : std_logic;
signal \N__58038\ : std_logic;
signal \N__58037\ : std_logic;
signal \N__58034\ : std_logic;
signal \N__58031\ : std_logic;
signal \N__58028\ : std_logic;
signal \N__58025\ : std_logic;
signal \N__58024\ : std_logic;
signal \N__58017\ : std_logic;
signal \N__58014\ : std_logic;
signal \N__58009\ : std_logic;
signal \N__58006\ : std_logic;
signal \N__58003\ : std_logic;
signal \N__58000\ : std_logic;
signal \N__57997\ : std_logic;
signal \N__57994\ : std_logic;
signal \N__57991\ : std_logic;
signal \N__57988\ : std_logic;
signal \N__57987\ : std_logic;
signal \N__57982\ : std_logic;
signal \N__57979\ : std_logic;
signal \N__57976\ : std_logic;
signal \N__57973\ : std_logic;
signal \N__57970\ : std_logic;
signal \N__57969\ : std_logic;
signal \N__57966\ : std_logic;
signal \N__57963\ : std_logic;
signal \N__57960\ : std_logic;
signal \N__57957\ : std_logic;
signal \N__57952\ : std_logic;
signal \N__57951\ : std_logic;
signal \N__57948\ : std_logic;
signal \N__57945\ : std_logic;
signal \N__57940\ : std_logic;
signal \N__57937\ : std_logic;
signal \N__57934\ : std_logic;
signal \N__57931\ : std_logic;
signal \N__57928\ : std_logic;
signal \N__57925\ : std_logic;
signal \N__57922\ : std_logic;
signal \N__57921\ : std_logic;
signal \N__57916\ : std_logic;
signal \N__57913\ : std_logic;
signal \N__57910\ : std_logic;
signal \N__57909\ : std_logic;
signal \N__57906\ : std_logic;
signal \N__57903\ : std_logic;
signal \N__57900\ : std_logic;
signal \N__57897\ : std_logic;
signal \N__57894\ : std_logic;
signal \N__57889\ : std_logic;
signal \N__57886\ : std_logic;
signal \N__57883\ : std_logic;
signal \N__57882\ : std_logic;
signal \N__57879\ : std_logic;
signal \N__57876\ : std_logic;
signal \N__57871\ : std_logic;
signal \N__57868\ : std_logic;
signal \N__57865\ : std_logic;
signal \N__57862\ : std_logic;
signal \N__57859\ : std_logic;
signal \N__57858\ : std_logic;
signal \N__57857\ : std_logic;
signal \N__57854\ : std_logic;
signal \N__57849\ : std_logic;
signal \N__57846\ : std_logic;
signal \N__57841\ : std_logic;
signal \N__57838\ : std_logic;
signal \N__57837\ : std_logic;
signal \N__57834\ : std_logic;
signal \N__57831\ : std_logic;
signal \N__57828\ : std_logic;
signal \N__57825\ : std_logic;
signal \N__57820\ : std_logic;
signal \N__57819\ : std_logic;
signal \N__57816\ : std_logic;
signal \N__57813\ : std_logic;
signal \N__57810\ : std_logic;
signal \N__57807\ : std_logic;
signal \N__57802\ : std_logic;
signal \N__57799\ : std_logic;
signal \N__57796\ : std_logic;
signal \N__57793\ : std_logic;
signal \N__57790\ : std_logic;
signal \N__57789\ : std_logic;
signal \N__57786\ : std_logic;
signal \N__57783\ : std_logic;
signal \N__57778\ : std_logic;
signal \N__57775\ : std_logic;
signal \N__57772\ : std_logic;
signal \N__57769\ : std_logic;
signal \N__57766\ : std_logic;
signal \N__57763\ : std_logic;
signal \N__57760\ : std_logic;
signal \N__57757\ : std_logic;
signal \N__57754\ : std_logic;
signal \N__57751\ : std_logic;
signal \N__57748\ : std_logic;
signal \N__57747\ : std_logic;
signal \N__57744\ : std_logic;
signal \N__57741\ : std_logic;
signal \N__57736\ : std_logic;
signal \N__57733\ : std_logic;
signal \N__57732\ : std_logic;
signal \N__57729\ : std_logic;
signal \N__57726\ : std_logic;
signal \N__57725\ : std_logic;
signal \N__57724\ : std_logic;
signal \N__57723\ : std_logic;
signal \N__57720\ : std_logic;
signal \N__57717\ : std_logic;
signal \N__57714\ : std_logic;
signal \N__57713\ : std_logic;
signal \N__57710\ : std_logic;
signal \N__57709\ : std_logic;
signal \N__57706\ : std_logic;
signal \N__57701\ : std_logic;
signal \N__57698\ : std_logic;
signal \N__57693\ : std_logic;
signal \N__57692\ : std_logic;
signal \N__57689\ : std_logic;
signal \N__57682\ : std_logic;
signal \N__57679\ : std_logic;
signal \N__57676\ : std_logic;
signal \N__57673\ : std_logic;
signal \N__57670\ : std_logic;
signal \N__57667\ : std_logic;
signal \N__57658\ : std_logic;
signal \N__57657\ : std_logic;
signal \N__57656\ : std_logic;
signal \N__57655\ : std_logic;
signal \N__57652\ : std_logic;
signal \N__57647\ : std_logic;
signal \N__57646\ : std_logic;
signal \N__57645\ : std_logic;
signal \N__57642\ : std_logic;
signal \N__57637\ : std_logic;
signal \N__57634\ : std_logic;
signal \N__57633\ : std_logic;
signal \N__57632\ : std_logic;
signal \N__57629\ : std_logic;
signal \N__57626\ : std_logic;
signal \N__57623\ : std_logic;
signal \N__57620\ : std_logic;
signal \N__57617\ : std_logic;
signal \N__57614\ : std_logic;
signal \N__57611\ : std_logic;
signal \N__57606\ : std_logic;
signal \N__57603\ : std_logic;
signal \N__57600\ : std_logic;
signal \N__57589\ : std_logic;
signal \N__57586\ : std_logic;
signal \N__57583\ : std_logic;
signal \N__57582\ : std_logic;
signal \N__57581\ : std_logic;
signal \N__57578\ : std_logic;
signal \N__57573\ : std_logic;
signal \N__57572\ : std_logic;
signal \N__57571\ : std_logic;
signal \N__57568\ : std_logic;
signal \N__57565\ : std_logic;
signal \N__57562\ : std_logic;
signal \N__57559\ : std_logic;
signal \N__57552\ : std_logic;
signal \N__57547\ : std_logic;
signal \N__57544\ : std_logic;
signal \N__57541\ : std_logic;
signal \N__57538\ : std_logic;
signal \N__57535\ : std_logic;
signal \N__57532\ : std_logic;
signal \N__57529\ : std_logic;
signal \N__57526\ : std_logic;
signal \N__57525\ : std_logic;
signal \N__57522\ : std_logic;
signal \N__57519\ : std_logic;
signal \N__57514\ : std_logic;
signal \N__57511\ : std_logic;
signal \N__57508\ : std_logic;
signal \N__57505\ : std_logic;
signal \N__57502\ : std_logic;
signal \N__57501\ : std_logic;
signal \N__57500\ : std_logic;
signal \N__57499\ : std_logic;
signal \N__57496\ : std_logic;
signal \N__57493\ : std_logic;
signal \N__57490\ : std_logic;
signal \N__57487\ : std_logic;
signal \N__57484\ : std_logic;
signal \N__57481\ : std_logic;
signal \N__57478\ : std_logic;
signal \N__57475\ : std_logic;
signal \N__57472\ : std_logic;
signal \N__57467\ : std_logic;
signal \N__57460\ : std_logic;
signal \N__57457\ : std_logic;
signal \N__57456\ : std_logic;
signal \N__57455\ : std_logic;
signal \N__57454\ : std_logic;
signal \N__57447\ : std_logic;
signal \N__57444\ : std_logic;
signal \N__57443\ : std_logic;
signal \N__57438\ : std_logic;
signal \N__57435\ : std_logic;
signal \N__57434\ : std_logic;
signal \N__57429\ : std_logic;
signal \N__57426\ : std_logic;
signal \N__57423\ : std_logic;
signal \N__57420\ : std_logic;
signal \N__57417\ : std_logic;
signal \N__57412\ : std_logic;
signal \N__57409\ : std_logic;
signal \N__57408\ : std_logic;
signal \N__57405\ : std_logic;
signal \N__57402\ : std_logic;
signal \N__57401\ : std_logic;
signal \N__57398\ : std_logic;
signal \N__57395\ : std_logic;
signal \N__57392\ : std_logic;
signal \N__57389\ : std_logic;
signal \N__57384\ : std_logic;
signal \N__57379\ : std_logic;
signal \N__57376\ : std_logic;
signal \N__57373\ : std_logic;
signal \N__57372\ : std_logic;
signal \N__57371\ : std_logic;
signal \N__57368\ : std_logic;
signal \N__57365\ : std_logic;
signal \N__57362\ : std_logic;
signal \N__57361\ : std_logic;
signal \N__57358\ : std_logic;
signal \N__57355\ : std_logic;
signal \N__57352\ : std_logic;
signal \N__57349\ : std_logic;
signal \N__57346\ : std_logic;
signal \N__57343\ : std_logic;
signal \N__57340\ : std_logic;
signal \N__57331\ : std_logic;
signal \N__57330\ : std_logic;
signal \N__57329\ : std_logic;
signal \N__57328\ : std_logic;
signal \N__57325\ : std_logic;
signal \N__57322\ : std_logic;
signal \N__57317\ : std_logic;
signal \N__57314\ : std_logic;
signal \N__57309\ : std_logic;
signal \N__57308\ : std_logic;
signal \N__57307\ : std_logic;
signal \N__57302\ : std_logic;
signal \N__57299\ : std_logic;
signal \N__57296\ : std_logic;
signal \N__57289\ : std_logic;
signal \N__57286\ : std_logic;
signal \N__57283\ : std_logic;
signal \N__57280\ : std_logic;
signal \N__57277\ : std_logic;
signal \N__57274\ : std_logic;
signal \N__57271\ : std_logic;
signal \N__57268\ : std_logic;
signal \N__57267\ : std_logic;
signal \N__57264\ : std_logic;
signal \N__57261\ : std_logic;
signal \N__57256\ : std_logic;
signal \N__57255\ : std_logic;
signal \N__57252\ : std_logic;
signal \N__57251\ : std_logic;
signal \N__57248\ : std_logic;
signal \N__57245\ : std_logic;
signal \N__57242\ : std_logic;
signal \N__57239\ : std_logic;
signal \N__57236\ : std_logic;
signal \N__57235\ : std_logic;
signal \N__57232\ : std_logic;
signal \N__57229\ : std_logic;
signal \N__57226\ : std_logic;
signal \N__57225\ : std_logic;
signal \N__57222\ : std_logic;
signal \N__57219\ : std_logic;
signal \N__57216\ : std_logic;
signal \N__57213\ : std_logic;
signal \N__57208\ : std_logic;
signal \N__57205\ : std_logic;
signal \N__57196\ : std_logic;
signal \N__57195\ : std_logic;
signal \N__57192\ : std_logic;
signal \N__57191\ : std_logic;
signal \N__57188\ : std_logic;
signal \N__57187\ : std_logic;
signal \N__57184\ : std_logic;
signal \N__57181\ : std_logic;
signal \N__57178\ : std_logic;
signal \N__57175\ : std_logic;
signal \N__57170\ : std_logic;
signal \N__57165\ : std_logic;
signal \N__57162\ : std_logic;
signal \N__57157\ : std_logic;
signal \N__57154\ : std_logic;
signal \N__57153\ : std_logic;
signal \N__57152\ : std_logic;
signal \N__57149\ : std_logic;
signal \N__57144\ : std_logic;
signal \N__57143\ : std_logic;
signal \N__57142\ : std_logic;
signal \N__57139\ : std_logic;
signal \N__57136\ : std_logic;
signal \N__57133\ : std_logic;
signal \N__57130\ : std_logic;
signal \N__57121\ : std_logic;
signal \N__57118\ : std_logic;
signal \N__57115\ : std_logic;
signal \N__57114\ : std_logic;
signal \N__57111\ : std_logic;
signal \N__57108\ : std_logic;
signal \N__57107\ : std_logic;
signal \N__57104\ : std_logic;
signal \N__57103\ : std_logic;
signal \N__57098\ : std_logic;
signal \N__57095\ : std_logic;
signal \N__57092\ : std_logic;
signal \N__57091\ : std_logic;
signal \N__57084\ : std_logic;
signal \N__57081\ : std_logic;
signal \N__57076\ : std_logic;
signal \N__57075\ : std_logic;
signal \N__57072\ : std_logic;
signal \N__57071\ : std_logic;
signal \N__57068\ : std_logic;
signal \N__57065\ : std_logic;
signal \N__57062\ : std_logic;
signal \N__57059\ : std_logic;
signal \N__57056\ : std_logic;
signal \N__57051\ : std_logic;
signal \N__57046\ : std_logic;
signal \N__57045\ : std_logic;
signal \N__57044\ : std_logic;
signal \N__57043\ : std_logic;
signal \N__57040\ : std_logic;
signal \N__57037\ : std_logic;
signal \N__57034\ : std_logic;
signal \N__57031\ : std_logic;
signal \N__57028\ : std_logic;
signal \N__57025\ : std_logic;
signal \N__57024\ : std_logic;
signal \N__57021\ : std_logic;
signal \N__57018\ : std_logic;
signal \N__57013\ : std_logic;
signal \N__57010\ : std_logic;
signal \N__57007\ : std_logic;
signal \N__57006\ : std_logic;
signal \N__57005\ : std_logic;
signal \N__57004\ : std_logic;
signal \N__57001\ : std_logic;
signal \N__56998\ : std_logic;
signal \N__56993\ : std_logic;
signal \N__56988\ : std_logic;
signal \N__56985\ : std_logic;
signal \N__56974\ : std_logic;
signal \N__56971\ : std_logic;
signal \N__56970\ : std_logic;
signal \N__56967\ : std_logic;
signal \N__56964\ : std_logic;
signal \N__56961\ : std_logic;
signal \N__56958\ : std_logic;
signal \N__56957\ : std_logic;
signal \N__56954\ : std_logic;
signal \N__56951\ : std_logic;
signal \N__56948\ : std_logic;
signal \N__56941\ : std_logic;
signal \N__56940\ : std_logic;
signal \N__56939\ : std_logic;
signal \N__56938\ : std_logic;
signal \N__56933\ : std_logic;
signal \N__56930\ : std_logic;
signal \N__56927\ : std_logic;
signal \N__56922\ : std_logic;
signal \N__56917\ : std_logic;
signal \N__56914\ : std_logic;
signal \N__56911\ : std_logic;
signal \N__56908\ : std_logic;
signal \N__56905\ : std_logic;
signal \N__56904\ : std_logic;
signal \N__56903\ : std_logic;
signal \N__56902\ : std_logic;
signal \N__56899\ : std_logic;
signal \N__56896\ : std_logic;
signal \N__56891\ : std_logic;
signal \N__56888\ : std_logic;
signal \N__56881\ : std_logic;
signal \N__56878\ : std_logic;
signal \N__56875\ : std_logic;
signal \N__56872\ : std_logic;
signal \N__56869\ : std_logic;
signal \N__56866\ : std_logic;
signal \N__56863\ : std_logic;
signal \N__56860\ : std_logic;
signal \N__56857\ : std_logic;
signal \N__56854\ : std_logic;
signal \N__56853\ : std_logic;
signal \N__56852\ : std_logic;
signal \N__56849\ : std_logic;
signal \N__56848\ : std_logic;
signal \N__56847\ : std_logic;
signal \N__56846\ : std_logic;
signal \N__56843\ : std_logic;
signal \N__56840\ : std_logic;
signal \N__56837\ : std_logic;
signal \N__56834\ : std_logic;
signal \N__56831\ : std_logic;
signal \N__56830\ : std_logic;
signal \N__56829\ : std_logic;
signal \N__56826\ : std_logic;
signal \N__56825\ : std_logic;
signal \N__56824\ : std_logic;
signal \N__56823\ : std_logic;
signal \N__56818\ : std_logic;
signal \N__56811\ : std_logic;
signal \N__56810\ : std_logic;
signal \N__56807\ : std_logic;
signal \N__56804\ : std_logic;
signal \N__56803\ : std_logic;
signal \N__56802\ : std_logic;
signal \N__56801\ : std_logic;
signal \N__56800\ : std_logic;
signal \N__56797\ : std_logic;
signal \N__56794\ : std_logic;
signal \N__56791\ : std_logic;
signal \N__56788\ : std_logic;
signal \N__56783\ : std_logic;
signal \N__56776\ : std_logic;
signal \N__56771\ : std_logic;
signal \N__56768\ : std_logic;
signal \N__56765\ : std_logic;
signal \N__56758\ : std_logic;
signal \N__56743\ : std_logic;
signal \N__56740\ : std_logic;
signal \N__56737\ : std_logic;
signal \N__56734\ : std_logic;
signal \N__56731\ : std_logic;
signal \N__56728\ : std_logic;
signal \N__56727\ : std_logic;
signal \N__56726\ : std_logic;
signal \N__56723\ : std_logic;
signal \N__56720\ : std_logic;
signal \N__56719\ : std_logic;
signal \N__56716\ : std_logic;
signal \N__56711\ : std_logic;
signal \N__56708\ : std_logic;
signal \N__56707\ : std_logic;
signal \N__56704\ : std_logic;
signal \N__56703\ : std_logic;
signal \N__56700\ : std_logic;
signal \N__56697\ : std_logic;
signal \N__56694\ : std_logic;
signal \N__56691\ : std_logic;
signal \N__56688\ : std_logic;
signal \N__56685\ : std_logic;
signal \N__56682\ : std_logic;
signal \N__56671\ : std_logic;
signal \N__56668\ : std_logic;
signal \N__56665\ : std_logic;
signal \N__56662\ : std_logic;
signal \N__56659\ : std_logic;
signal \N__56656\ : std_logic;
signal \N__56653\ : std_logic;
signal \N__56652\ : std_logic;
signal \N__56651\ : std_logic;
signal \N__56650\ : std_logic;
signal \N__56647\ : std_logic;
signal \N__56646\ : std_logic;
signal \N__56643\ : std_logic;
signal \N__56642\ : std_logic;
signal \N__56637\ : std_logic;
signal \N__56634\ : std_logic;
signal \N__56631\ : std_logic;
signal \N__56630\ : std_logic;
signal \N__56629\ : std_logic;
signal \N__56626\ : std_logic;
signal \N__56623\ : std_logic;
signal \N__56620\ : std_logic;
signal \N__56617\ : std_logic;
signal \N__56614\ : std_logic;
signal \N__56611\ : std_logic;
signal \N__56608\ : std_logic;
signal \N__56605\ : std_logic;
signal \N__56602\ : std_logic;
signal \N__56599\ : std_logic;
signal \N__56594\ : std_logic;
signal \N__56591\ : std_logic;
signal \N__56578\ : std_logic;
signal \N__56575\ : std_logic;
signal \N__56572\ : std_logic;
signal \N__56569\ : std_logic;
signal \N__56566\ : std_logic;
signal \N__56563\ : std_logic;
signal \N__56562\ : std_logic;
signal \N__56561\ : std_logic;
signal \N__56560\ : std_logic;
signal \N__56557\ : std_logic;
signal \N__56552\ : std_logic;
signal \N__56549\ : std_logic;
signal \N__56546\ : std_logic;
signal \N__56543\ : std_logic;
signal \N__56540\ : std_logic;
signal \N__56533\ : std_logic;
signal \N__56530\ : std_logic;
signal \N__56529\ : std_logic;
signal \N__56528\ : std_logic;
signal \N__56525\ : std_logic;
signal \N__56524\ : std_logic;
signal \N__56521\ : std_logic;
signal \N__56518\ : std_logic;
signal \N__56515\ : std_logic;
signal \N__56512\ : std_logic;
signal \N__56509\ : std_logic;
signal \N__56504\ : std_logic;
signal \N__56501\ : std_logic;
signal \N__56498\ : std_logic;
signal \N__56495\ : std_logic;
signal \N__56488\ : std_logic;
signal \N__56485\ : std_logic;
signal \N__56484\ : std_logic;
signal \N__56481\ : std_logic;
signal \N__56478\ : std_logic;
signal \N__56475\ : std_logic;
signal \N__56470\ : std_logic;
signal \N__56467\ : std_logic;
signal \N__56464\ : std_logic;
signal \N__56461\ : std_logic;
signal \N__56458\ : std_logic;
signal \N__56455\ : std_logic;
signal \N__56452\ : std_logic;
signal \N__56451\ : std_logic;
signal \N__56450\ : std_logic;
signal \N__56447\ : std_logic;
signal \N__56442\ : std_logic;
signal \N__56441\ : std_logic;
signal \N__56440\ : std_logic;
signal \N__56437\ : std_logic;
signal \N__56434\ : std_logic;
signal \N__56429\ : std_logic;
signal \N__56426\ : std_logic;
signal \N__56421\ : std_logic;
signal \N__56418\ : std_logic;
signal \N__56413\ : std_logic;
signal \N__56410\ : std_logic;
signal \N__56409\ : std_logic;
signal \N__56406\ : std_logic;
signal \N__56403\ : std_logic;
signal \N__56400\ : std_logic;
signal \N__56399\ : std_logic;
signal \N__56398\ : std_logic;
signal \N__56393\ : std_logic;
signal \N__56390\ : std_logic;
signal \N__56387\ : std_logic;
signal \N__56384\ : std_logic;
signal \N__56379\ : std_logic;
signal \N__56378\ : std_logic;
signal \N__56373\ : std_logic;
signal \N__56370\ : std_logic;
signal \N__56365\ : std_logic;
signal \N__56362\ : std_logic;
signal \N__56359\ : std_logic;
signal \N__56356\ : std_logic;
signal \N__56353\ : std_logic;
signal \N__56352\ : std_logic;
signal \N__56351\ : std_logic;
signal \N__56348\ : std_logic;
signal \N__56345\ : std_logic;
signal \N__56342\ : std_logic;
signal \N__56341\ : std_logic;
signal \N__56338\ : std_logic;
signal \N__56335\ : std_logic;
signal \N__56332\ : std_logic;
signal \N__56329\ : std_logic;
signal \N__56326\ : std_logic;
signal \N__56323\ : std_logic;
signal \N__56314\ : std_logic;
signal \N__56313\ : std_logic;
signal \N__56308\ : std_logic;
signal \N__56305\ : std_logic;
signal \N__56302\ : std_logic;
signal \N__56299\ : std_logic;
signal \N__56296\ : std_logic;
signal \N__56295\ : std_logic;
signal \N__56292\ : std_logic;
signal \N__56291\ : std_logic;
signal \N__56290\ : std_logic;
signal \N__56287\ : std_logic;
signal \N__56284\ : std_logic;
signal \N__56279\ : std_logic;
signal \N__56272\ : std_logic;
signal \N__56269\ : std_logic;
signal \N__56266\ : std_logic;
signal \N__56263\ : std_logic;
signal \N__56260\ : std_logic;
signal \N__56259\ : std_logic;
signal \N__56256\ : std_logic;
signal \N__56253\ : std_logic;
signal \N__56248\ : std_logic;
signal \N__56245\ : std_logic;
signal \N__56242\ : std_logic;
signal \N__56239\ : std_logic;
signal \N__56238\ : std_logic;
signal \N__56237\ : std_logic;
signal \N__56236\ : std_logic;
signal \N__56233\ : std_logic;
signal \N__56230\ : std_logic;
signal \N__56227\ : std_logic;
signal \N__56226\ : std_logic;
signal \N__56225\ : std_logic;
signal \N__56224\ : std_logic;
signal \N__56221\ : std_logic;
signal \N__56214\ : std_logic;
signal \N__56213\ : std_logic;
signal \N__56210\ : std_logic;
signal \N__56207\ : std_logic;
signal \N__56204\ : std_logic;
signal \N__56201\ : std_logic;
signal \N__56200\ : std_logic;
signal \N__56197\ : std_logic;
signal \N__56194\ : std_logic;
signal \N__56193\ : std_logic;
signal \N__56188\ : std_logic;
signal \N__56185\ : std_logic;
signal \N__56182\ : std_logic;
signal \N__56179\ : std_logic;
signal \N__56176\ : std_logic;
signal \N__56173\ : std_logic;
signal \N__56170\ : std_logic;
signal \N__56167\ : std_logic;
signal \N__56164\ : std_logic;
signal \N__56161\ : std_logic;
signal \N__56158\ : std_logic;
signal \N__56155\ : std_logic;
signal \N__56154\ : std_logic;
signal \N__56149\ : std_logic;
signal \N__56146\ : std_logic;
signal \N__56143\ : std_logic;
signal \N__56140\ : std_logic;
signal \N__56135\ : std_logic;
signal \N__56132\ : std_logic;
signal \N__56127\ : std_logic;
signal \N__56126\ : std_logic;
signal \N__56123\ : std_logic;
signal \N__56120\ : std_logic;
signal \N__56117\ : std_logic;
signal \N__56114\ : std_logic;
signal \N__56111\ : std_logic;
signal \N__56108\ : std_logic;
signal \N__56103\ : std_logic;
signal \N__56098\ : std_logic;
signal \N__56093\ : std_logic;
signal \N__56086\ : std_logic;
signal \N__56085\ : std_logic;
signal \N__56084\ : std_logic;
signal \N__56081\ : std_logic;
signal \N__56080\ : std_logic;
signal \N__56077\ : std_logic;
signal \N__56074\ : std_logic;
signal \N__56071\ : std_logic;
signal \N__56068\ : std_logic;
signal \N__56065\ : std_logic;
signal \N__56062\ : std_logic;
signal \N__56059\ : std_logic;
signal \N__56056\ : std_logic;
signal \N__56053\ : std_logic;
signal \N__56048\ : std_logic;
signal \N__56043\ : std_logic;
signal \N__56040\ : std_logic;
signal \N__56035\ : std_logic;
signal \N__56032\ : std_logic;
signal \N__56029\ : std_logic;
signal \N__56028\ : std_logic;
signal \N__56027\ : std_logic;
signal \N__56024\ : std_logic;
signal \N__56021\ : std_logic;
signal \N__56018\ : std_logic;
signal \N__56017\ : std_logic;
signal \N__56014\ : std_logic;
signal \N__56011\ : std_logic;
signal \N__56008\ : std_logic;
signal \N__56005\ : std_logic;
signal \N__56002\ : std_logic;
signal \N__55999\ : std_logic;
signal \N__55996\ : std_logic;
signal \N__55993\ : std_logic;
signal \N__55988\ : std_logic;
signal \N__55985\ : std_logic;
signal \N__55978\ : std_logic;
signal \N__55975\ : std_logic;
signal \N__55972\ : std_logic;
signal \N__55969\ : std_logic;
signal \N__55966\ : std_logic;
signal \N__55963\ : std_logic;
signal \N__55960\ : std_logic;
signal \N__55959\ : std_logic;
signal \N__55956\ : std_logic;
signal \N__55953\ : std_logic;
signal \N__55952\ : std_logic;
signal \N__55951\ : std_logic;
signal \N__55948\ : std_logic;
signal \N__55945\ : std_logic;
signal \N__55942\ : std_logic;
signal \N__55939\ : std_logic;
signal \N__55932\ : std_logic;
signal \N__55929\ : std_logic;
signal \N__55926\ : std_logic;
signal \N__55921\ : std_logic;
signal \N__55920\ : std_logic;
signal \N__55919\ : std_logic;
signal \N__55916\ : std_logic;
signal \N__55913\ : std_logic;
signal \N__55910\ : std_logic;
signal \N__55907\ : std_logic;
signal \N__55904\ : std_logic;
signal \N__55901\ : std_logic;
signal \N__55898\ : std_logic;
signal \N__55893\ : std_logic;
signal \N__55888\ : std_logic;
signal \N__55887\ : std_logic;
signal \N__55886\ : std_logic;
signal \N__55885\ : std_logic;
signal \N__55884\ : std_logic;
signal \N__55883\ : std_logic;
signal \N__55880\ : std_logic;
signal \N__55877\ : std_logic;
signal \N__55876\ : std_logic;
signal \N__55875\ : std_logic;
signal \N__55874\ : std_logic;
signal \N__55873\ : std_logic;
signal \N__55872\ : std_logic;
signal \N__55869\ : std_logic;
signal \N__55868\ : std_logic;
signal \N__55867\ : std_logic;
signal \N__55862\ : std_logic;
signal \N__55859\ : std_logic;
signal \N__55854\ : std_logic;
signal \N__55849\ : std_logic;
signal \N__55842\ : std_logic;
signal \N__55839\ : std_logic;
signal \N__55836\ : std_logic;
signal \N__55833\ : std_logic;
signal \N__55828\ : std_logic;
signal \N__55825\ : std_logic;
signal \N__55820\ : std_logic;
signal \N__55819\ : std_logic;
signal \N__55816\ : std_logic;
signal \N__55813\ : std_logic;
signal \N__55812\ : std_logic;
signal \N__55809\ : std_logic;
signal \N__55806\ : std_logic;
signal \N__55801\ : std_logic;
signal \N__55800\ : std_logic;
signal \N__55797\ : std_logic;
signal \N__55796\ : std_logic;
signal \N__55795\ : std_logic;
signal \N__55792\ : std_logic;
signal \N__55789\ : std_logic;
signal \N__55786\ : std_logic;
signal \N__55783\ : std_logic;
signal \N__55778\ : std_logic;
signal \N__55775\ : std_logic;
signal \N__55768\ : std_logic;
signal \N__55765\ : std_logic;
signal \N__55762\ : std_logic;
signal \N__55757\ : std_logic;
signal \N__55754\ : std_logic;
signal \N__55747\ : std_logic;
signal \N__55742\ : std_logic;
signal \N__55737\ : std_logic;
signal \N__55732\ : std_logic;
signal \N__55729\ : std_logic;
signal \N__55726\ : std_logic;
signal \N__55725\ : std_logic;
signal \N__55724\ : std_logic;
signal \N__55721\ : std_logic;
signal \N__55718\ : std_logic;
signal \N__55715\ : std_logic;
signal \N__55708\ : std_logic;
signal \N__55705\ : std_logic;
signal \N__55704\ : std_logic;
signal \N__55701\ : std_logic;
signal \N__55698\ : std_logic;
signal \N__55697\ : std_logic;
signal \N__55696\ : std_logic;
signal \N__55693\ : std_logic;
signal \N__55690\ : std_logic;
signal \N__55685\ : std_logic;
signal \N__55678\ : std_logic;
signal \N__55675\ : std_logic;
signal \N__55672\ : std_logic;
signal \N__55671\ : std_logic;
signal \N__55670\ : std_logic;
signal \N__55669\ : std_logic;
signal \N__55668\ : std_logic;
signal \N__55665\ : std_logic;
signal \N__55662\ : std_logic;
signal \N__55659\ : std_logic;
signal \N__55656\ : std_logic;
signal \N__55653\ : std_logic;
signal \N__55650\ : std_logic;
signal \N__55647\ : std_logic;
signal \N__55642\ : std_logic;
signal \N__55639\ : std_logic;
signal \N__55636\ : std_logic;
signal \N__55631\ : std_logic;
signal \N__55628\ : std_logic;
signal \N__55623\ : std_logic;
signal \N__55618\ : std_logic;
signal \N__55615\ : std_logic;
signal \N__55614\ : std_logic;
signal \N__55611\ : std_logic;
signal \N__55610\ : std_logic;
signal \N__55607\ : std_logic;
signal \N__55604\ : std_logic;
signal \N__55601\ : std_logic;
signal \N__55598\ : std_logic;
signal \N__55593\ : std_logic;
signal \N__55588\ : std_logic;
signal \N__55587\ : std_logic;
signal \N__55586\ : std_logic;
signal \N__55585\ : std_logic;
signal \N__55584\ : std_logic;
signal \N__55583\ : std_logic;
signal \N__55580\ : std_logic;
signal \N__55575\ : std_logic;
signal \N__55572\ : std_logic;
signal \N__55569\ : std_logic;
signal \N__55566\ : std_logic;
signal \N__55559\ : std_logic;
signal \N__55556\ : std_logic;
signal \N__55549\ : std_logic;
signal \N__55548\ : std_logic;
signal \N__55545\ : std_logic;
signal \N__55544\ : std_logic;
signal \N__55541\ : std_logic;
signal \N__55540\ : std_logic;
signal \N__55537\ : std_logic;
signal \N__55532\ : std_logic;
signal \N__55529\ : std_logic;
signal \N__55526\ : std_logic;
signal \N__55523\ : std_logic;
signal \N__55516\ : std_logic;
signal \N__55515\ : std_logic;
signal \N__55512\ : std_logic;
signal \N__55511\ : std_logic;
signal \N__55510\ : std_logic;
signal \N__55509\ : std_logic;
signal \N__55506\ : std_logic;
signal \N__55505\ : std_logic;
signal \N__55502\ : std_logic;
signal \N__55499\ : std_logic;
signal \N__55496\ : std_logic;
signal \N__55493\ : std_logic;
signal \N__55490\ : std_logic;
signal \N__55487\ : std_logic;
signal \N__55484\ : std_logic;
signal \N__55477\ : std_logic;
signal \N__55468\ : std_logic;
signal \N__55467\ : std_logic;
signal \N__55466\ : std_logic;
signal \N__55465\ : std_logic;
signal \N__55462\ : std_logic;
signal \N__55459\ : std_logic;
signal \N__55454\ : std_logic;
signal \N__55451\ : std_logic;
signal \N__55448\ : std_logic;
signal \N__55445\ : std_logic;
signal \N__55442\ : std_logic;
signal \N__55439\ : std_logic;
signal \N__55436\ : std_logic;
signal \N__55433\ : std_logic;
signal \N__55430\ : std_logic;
signal \N__55425\ : std_logic;
signal \N__55420\ : std_logic;
signal \N__55417\ : std_logic;
signal \N__55414\ : std_logic;
signal \N__55411\ : std_logic;
signal \N__55408\ : std_logic;
signal \N__55405\ : std_logic;
signal \N__55402\ : std_logic;
signal \N__55399\ : std_logic;
signal \N__55396\ : std_logic;
signal \N__55393\ : std_logic;
signal \N__55390\ : std_logic;
signal \N__55387\ : std_logic;
signal \N__55384\ : std_logic;
signal \N__55383\ : std_logic;
signal \N__55382\ : std_logic;
signal \N__55379\ : std_logic;
signal \N__55378\ : std_logic;
signal \N__55377\ : std_logic;
signal \N__55374\ : std_logic;
signal \N__55371\ : std_logic;
signal \N__55368\ : std_logic;
signal \N__55365\ : std_logic;
signal \N__55364\ : std_logic;
signal \N__55361\ : std_logic;
signal \N__55358\ : std_logic;
signal \N__55355\ : std_logic;
signal \N__55350\ : std_logic;
signal \N__55349\ : std_logic;
signal \N__55346\ : std_logic;
signal \N__55345\ : std_logic;
signal \N__55344\ : std_logic;
signal \N__55341\ : std_logic;
signal \N__55338\ : std_logic;
signal \N__55333\ : std_logic;
signal \N__55330\ : std_logic;
signal \N__55327\ : std_logic;
signal \N__55322\ : std_logic;
signal \N__55309\ : std_logic;
signal \N__55308\ : std_logic;
signal \N__55305\ : std_logic;
signal \N__55300\ : std_logic;
signal \N__55297\ : std_logic;
signal \N__55294\ : std_logic;
signal \N__55291\ : std_logic;
signal \N__55288\ : std_logic;
signal \N__55285\ : std_logic;
signal \N__55284\ : std_logic;
signal \N__55281\ : std_logic;
signal \N__55278\ : std_logic;
signal \N__55277\ : std_logic;
signal \N__55272\ : std_logic;
signal \N__55269\ : std_logic;
signal \N__55264\ : std_logic;
signal \N__55263\ : std_logic;
signal \N__55260\ : std_logic;
signal \N__55257\ : std_logic;
signal \N__55254\ : std_logic;
signal \N__55251\ : std_logic;
signal \N__55248\ : std_logic;
signal \N__55245\ : std_logic;
signal \N__55240\ : std_logic;
signal \N__55239\ : std_logic;
signal \N__55236\ : std_logic;
signal \N__55235\ : std_logic;
signal \N__55234\ : std_logic;
signal \N__55231\ : std_logic;
signal \N__55228\ : std_logic;
signal \N__55225\ : std_logic;
signal \N__55222\ : std_logic;
signal \N__55219\ : std_logic;
signal \N__55214\ : std_logic;
signal \N__55213\ : std_logic;
signal \N__55212\ : std_logic;
signal \N__55209\ : std_logic;
signal \N__55206\ : std_logic;
signal \N__55203\ : std_logic;
signal \N__55200\ : std_logic;
signal \N__55197\ : std_logic;
signal \N__55186\ : std_logic;
signal \N__55185\ : std_logic;
signal \N__55184\ : std_logic;
signal \N__55183\ : std_logic;
signal \N__55182\ : std_logic;
signal \N__55181\ : std_logic;
signal \N__55180\ : std_logic;
signal \N__55179\ : std_logic;
signal \N__55178\ : std_logic;
signal \N__55175\ : std_logic;
signal \N__55172\ : std_logic;
signal \N__55169\ : std_logic;
signal \N__55166\ : std_logic;
signal \N__55165\ : std_logic;
signal \N__55164\ : std_logic;
signal \N__55163\ : std_logic;
signal \N__55162\ : std_logic;
signal \N__55157\ : std_logic;
signal \N__55154\ : std_logic;
signal \N__55151\ : std_logic;
signal \N__55148\ : std_logic;
signal \N__55147\ : std_logic;
signal \N__55144\ : std_logic;
signal \N__55137\ : std_logic;
signal \N__55130\ : std_logic;
signal \N__55129\ : std_logic;
signal \N__55128\ : std_logic;
signal \N__55127\ : std_logic;
signal \N__55124\ : std_logic;
signal \N__55121\ : std_logic;
signal \N__55118\ : std_logic;
signal \N__55115\ : std_logic;
signal \N__55110\ : std_logic;
signal \N__55109\ : std_logic;
signal \N__55108\ : std_logic;
signal \N__55105\ : std_logic;
signal \N__55100\ : std_logic;
signal \N__55095\ : std_logic;
signal \N__55092\ : std_logic;
signal \N__55089\ : std_logic;
signal \N__55080\ : std_logic;
signal \N__55077\ : std_logic;
signal \N__55074\ : std_logic;
signal \N__55069\ : std_logic;
signal \N__55054\ : std_logic;
signal \N__55053\ : std_logic;
signal \N__55052\ : std_logic;
signal \N__55049\ : std_logic;
signal \N__55046\ : std_logic;
signal \N__55043\ : std_logic;
signal \N__55040\ : std_logic;
signal \N__55035\ : std_logic;
signal \N__55034\ : std_logic;
signal \N__55033\ : std_logic;
signal \N__55032\ : std_logic;
signal \N__55031\ : std_logic;
signal \N__55028\ : std_logic;
signal \N__55025\ : std_logic;
signal \N__55022\ : std_logic;
signal \N__55017\ : std_logic;
signal \N__55016\ : std_logic;
signal \N__55015\ : std_logic;
signal \N__55014\ : std_logic;
signal \N__55011\ : std_logic;
signal \N__55010\ : std_logic;
signal \N__55007\ : std_logic;
signal \N__55000\ : std_logic;
signal \N__54995\ : std_logic;
signal \N__54992\ : std_logic;
signal \N__54987\ : std_logic;
signal \N__54976\ : std_logic;
signal \N__54973\ : std_logic;
signal \N__54970\ : std_logic;
signal \N__54967\ : std_logic;
signal \N__54966\ : std_logic;
signal \N__54965\ : std_logic;
signal \N__54962\ : std_logic;
signal \N__54957\ : std_logic;
signal \N__54952\ : std_logic;
signal \N__54949\ : std_logic;
signal \N__54946\ : std_logic;
signal \N__54943\ : std_logic;
signal \N__54940\ : std_logic;
signal \N__54937\ : std_logic;
signal \N__54934\ : std_logic;
signal \N__54931\ : std_logic;
signal \N__54928\ : std_logic;
signal \N__54925\ : std_logic;
signal \N__54922\ : std_logic;
signal \N__54919\ : std_logic;
signal \N__54916\ : std_logic;
signal \N__54913\ : std_logic;
signal \N__54910\ : std_logic;
signal \N__54907\ : std_logic;
signal \N__54904\ : std_logic;
signal \N__54901\ : std_logic;
signal \N__54898\ : std_logic;
signal \N__54895\ : std_logic;
signal \N__54894\ : std_logic;
signal \N__54893\ : std_logic;
signal \N__54892\ : std_logic;
signal \N__54889\ : std_logic;
signal \N__54888\ : std_logic;
signal \N__54887\ : std_logic;
signal \N__54884\ : std_logic;
signal \N__54881\ : std_logic;
signal \N__54880\ : std_logic;
signal \N__54877\ : std_logic;
signal \N__54876\ : std_logic;
signal \N__54873\ : std_logic;
signal \N__54868\ : std_logic;
signal \N__54865\ : std_logic;
signal \N__54862\ : std_logic;
signal \N__54859\ : std_logic;
signal \N__54858\ : std_logic;
signal \N__54855\ : std_logic;
signal \N__54852\ : std_logic;
signal \N__54851\ : std_logic;
signal \N__54846\ : std_logic;
signal \N__54843\ : std_logic;
signal \N__54842\ : std_logic;
signal \N__54837\ : std_logic;
signal \N__54836\ : std_logic;
signal \N__54835\ : std_logic;
signal \N__54834\ : std_logic;
signal \N__54831\ : std_logic;
signal \N__54828\ : std_logic;
signal \N__54825\ : std_logic;
signal \N__54822\ : std_logic;
signal \N__54819\ : std_logic;
signal \N__54816\ : std_logic;
signal \N__54813\ : std_logic;
signal \N__54810\ : std_logic;
signal \N__54807\ : std_logic;
signal \N__54800\ : std_logic;
signal \N__54781\ : std_logic;
signal \N__54778\ : std_logic;
signal \N__54775\ : std_logic;
signal \N__54772\ : std_logic;
signal \N__54771\ : std_logic;
signal \N__54770\ : std_logic;
signal \N__54767\ : std_logic;
signal \N__54762\ : std_logic;
signal \N__54757\ : std_logic;
signal \N__54754\ : std_logic;
signal \N__54751\ : std_logic;
signal \N__54750\ : std_logic;
signal \N__54747\ : std_logic;
signal \N__54744\ : std_logic;
signal \N__54741\ : std_logic;
signal \N__54738\ : std_logic;
signal \N__54733\ : std_logic;
signal \N__54732\ : std_logic;
signal \N__54731\ : std_logic;
signal \N__54728\ : std_logic;
signal \N__54727\ : std_logic;
signal \N__54722\ : std_logic;
signal \N__54719\ : std_logic;
signal \N__54716\ : std_logic;
signal \N__54713\ : std_logic;
signal \N__54706\ : std_logic;
signal \N__54703\ : std_logic;
signal \N__54700\ : std_logic;
signal \N__54697\ : std_logic;
signal \N__54694\ : std_logic;
signal \N__54691\ : std_logic;
signal \N__54688\ : std_logic;
signal \N__54685\ : std_logic;
signal \N__54684\ : std_logic;
signal \N__54681\ : std_logic;
signal \N__54680\ : std_logic;
signal \N__54677\ : std_logic;
signal \N__54676\ : std_logic;
signal \N__54675\ : std_logic;
signal \N__54674\ : std_logic;
signal \N__54673\ : std_logic;
signal \N__54672\ : std_logic;
signal \N__54671\ : std_logic;
signal \N__54668\ : std_logic;
signal \N__54665\ : std_logic;
signal \N__54658\ : std_logic;
signal \N__54655\ : std_logic;
signal \N__54652\ : std_logic;
signal \N__54647\ : std_logic;
signal \N__54634\ : std_logic;
signal \N__54631\ : std_logic;
signal \N__54628\ : std_logic;
signal \N__54627\ : std_logic;
signal \N__54624\ : std_logic;
signal \N__54623\ : std_logic;
signal \N__54620\ : std_logic;
signal \N__54617\ : std_logic;
signal \N__54614\ : std_logic;
signal \N__54613\ : std_logic;
signal \N__54612\ : std_logic;
signal \N__54609\ : std_logic;
signal \N__54606\ : std_logic;
signal \N__54603\ : std_logic;
signal \N__54598\ : std_logic;
signal \N__54589\ : std_logic;
signal \N__54586\ : std_logic;
signal \N__54583\ : std_logic;
signal \N__54580\ : std_logic;
signal \N__54579\ : std_logic;
signal \N__54576\ : std_logic;
signal \N__54571\ : std_logic;
signal \N__54568\ : std_logic;
signal \N__54567\ : std_logic;
signal \N__54564\ : std_logic;
signal \N__54561\ : std_logic;
signal \N__54560\ : std_logic;
signal \N__54557\ : std_logic;
signal \N__54556\ : std_logic;
signal \N__54553\ : std_logic;
signal \N__54550\ : std_logic;
signal \N__54547\ : std_logic;
signal \N__54544\ : std_logic;
signal \N__54541\ : std_logic;
signal \N__54532\ : std_logic;
signal \N__54531\ : std_logic;
signal \N__54530\ : std_logic;
signal \N__54525\ : std_logic;
signal \N__54522\ : std_logic;
signal \N__54519\ : std_logic;
signal \N__54518\ : std_logic;
signal \N__54515\ : std_logic;
signal \N__54512\ : std_logic;
signal \N__54509\ : std_logic;
signal \N__54502\ : std_logic;
signal \N__54499\ : std_logic;
signal \N__54496\ : std_logic;
signal \N__54493\ : std_logic;
signal \N__54492\ : std_logic;
signal \N__54489\ : std_logic;
signal \N__54486\ : std_logic;
signal \N__54481\ : std_logic;
signal \N__54480\ : std_logic;
signal \N__54479\ : std_logic;
signal \N__54476\ : std_logic;
signal \N__54473\ : std_logic;
signal \N__54472\ : std_logic;
signal \N__54469\ : std_logic;
signal \N__54468\ : std_logic;
signal \N__54467\ : std_logic;
signal \N__54466\ : std_logic;
signal \N__54463\ : std_logic;
signal \N__54462\ : std_logic;
signal \N__54461\ : std_logic;
signal \N__54460\ : std_logic;
signal \N__54459\ : std_logic;
signal \N__54456\ : std_logic;
signal \N__54453\ : std_logic;
signal \N__54452\ : std_logic;
signal \N__54449\ : std_logic;
signal \N__54446\ : std_logic;
signal \N__54443\ : std_logic;
signal \N__54442\ : std_logic;
signal \N__54439\ : std_logic;
signal \N__54436\ : std_logic;
signal \N__54431\ : std_logic;
signal \N__54428\ : std_logic;
signal \N__54427\ : std_logic;
signal \N__54424\ : std_logic;
signal \N__54423\ : std_logic;
signal \N__54422\ : std_logic;
signal \N__54421\ : std_logic;
signal \N__54418\ : std_logic;
signal \N__54415\ : std_logic;
signal \N__54412\ : std_logic;
signal \N__54411\ : std_logic;
signal \N__54410\ : std_logic;
signal \N__54405\ : std_logic;
signal \N__54402\ : std_logic;
signal \N__54399\ : std_logic;
signal \N__54396\ : std_logic;
signal \N__54395\ : std_logic;
signal \N__54388\ : std_logic;
signal \N__54385\ : std_logic;
signal \N__54384\ : std_logic;
signal \N__54383\ : std_logic;
signal \N__54378\ : std_logic;
signal \N__54373\ : std_logic;
signal \N__54370\ : std_logic;
signal \N__54365\ : std_logic;
signal \N__54360\ : std_logic;
signal \N__54351\ : std_logic;
signal \N__54348\ : std_logic;
signal \N__54343\ : std_logic;
signal \N__54340\ : std_logic;
signal \N__54337\ : std_logic;
signal \N__54316\ : std_logic;
signal \N__54315\ : std_logic;
signal \N__54312\ : std_logic;
signal \N__54309\ : std_logic;
signal \N__54308\ : std_logic;
signal \N__54305\ : std_logic;
signal \N__54302\ : std_logic;
signal \N__54299\ : std_logic;
signal \N__54298\ : std_logic;
signal \N__54297\ : std_logic;
signal \N__54296\ : std_logic;
signal \N__54291\ : std_logic;
signal \N__54288\ : std_logic;
signal \N__54285\ : std_logic;
signal \N__54280\ : std_logic;
signal \N__54271\ : std_logic;
signal \N__54268\ : std_logic;
signal \N__54267\ : std_logic;
signal \N__54266\ : std_logic;
signal \N__54263\ : std_logic;
signal \N__54262\ : std_logic;
signal \N__54261\ : std_logic;
signal \N__54258\ : std_logic;
signal \N__54255\ : std_logic;
signal \N__54254\ : std_logic;
signal \N__54251\ : std_logic;
signal \N__54246\ : std_logic;
signal \N__54243\ : std_logic;
signal \N__54242\ : std_logic;
signal \N__54239\ : std_logic;
signal \N__54236\ : std_logic;
signal \N__54233\ : std_logic;
signal \N__54230\ : std_logic;
signal \N__54227\ : std_logic;
signal \N__54224\ : std_logic;
signal \N__54211\ : std_logic;
signal \N__54210\ : std_logic;
signal \N__54205\ : std_logic;
signal \N__54202\ : std_logic;
signal \N__54199\ : std_logic;
signal \N__54198\ : std_logic;
signal \N__54195\ : std_logic;
signal \N__54192\ : std_logic;
signal \N__54187\ : std_logic;
signal \N__54186\ : std_logic;
signal \N__54185\ : std_logic;
signal \N__54178\ : std_logic;
signal \N__54175\ : std_logic;
signal \N__54172\ : std_logic;
signal \N__54169\ : std_logic;
signal \N__54166\ : std_logic;
signal \N__54163\ : std_logic;
signal \N__54162\ : std_logic;
signal \N__54159\ : std_logic;
signal \N__54156\ : std_logic;
signal \N__54155\ : std_logic;
signal \N__54152\ : std_logic;
signal \N__54149\ : std_logic;
signal \N__54146\ : std_logic;
signal \N__54143\ : std_logic;
signal \N__54136\ : std_logic;
signal \N__54135\ : std_logic;
signal \N__54134\ : std_logic;
signal \N__54131\ : std_logic;
signal \N__54130\ : std_logic;
signal \N__54127\ : std_logic;
signal \N__54126\ : std_logic;
signal \N__54123\ : std_logic;
signal \N__54122\ : std_logic;
signal \N__54119\ : std_logic;
signal \N__54116\ : std_logic;
signal \N__54115\ : std_logic;
signal \N__54112\ : std_logic;
signal \N__54109\ : std_logic;
signal \N__54106\ : std_logic;
signal \N__54103\ : std_logic;
signal \N__54098\ : std_logic;
signal \N__54097\ : std_logic;
signal \N__54096\ : std_logic;
signal \N__54095\ : std_logic;
signal \N__54094\ : std_logic;
signal \N__54091\ : std_logic;
signal \N__54088\ : std_logic;
signal \N__54079\ : std_logic;
signal \N__54070\ : std_logic;
signal \N__54067\ : std_logic;
signal \N__54058\ : std_logic;
signal \N__54055\ : std_logic;
signal \N__54054\ : std_logic;
signal \N__54051\ : std_logic;
signal \N__54048\ : std_logic;
signal \N__54045\ : std_logic;
signal \N__54042\ : std_logic;
signal \N__54039\ : std_logic;
signal \N__54036\ : std_logic;
signal \N__54031\ : std_logic;
signal \N__54028\ : std_logic;
signal \N__54025\ : std_logic;
signal \N__54022\ : std_logic;
signal \N__54021\ : std_logic;
signal \N__54020\ : std_logic;
signal \N__54017\ : std_logic;
signal \N__54014\ : std_logic;
signal \N__54011\ : std_logic;
signal \N__54008\ : std_logic;
signal \N__54005\ : std_logic;
signal \N__54002\ : std_logic;
signal \N__53999\ : std_logic;
signal \N__53996\ : std_logic;
signal \N__53993\ : std_logic;
signal \N__53986\ : std_logic;
signal \N__53983\ : std_logic;
signal \N__53980\ : std_logic;
signal \N__53977\ : std_logic;
signal \N__53974\ : std_logic;
signal \N__53973\ : std_logic;
signal \N__53970\ : std_logic;
signal \N__53967\ : std_logic;
signal \N__53964\ : std_logic;
signal \N__53963\ : std_logic;
signal \N__53960\ : std_logic;
signal \N__53957\ : std_logic;
signal \N__53954\ : std_logic;
signal \N__53947\ : std_logic;
signal \N__53944\ : std_logic;
signal \N__53943\ : std_logic;
signal \N__53942\ : std_logic;
signal \N__53939\ : std_logic;
signal \N__53936\ : std_logic;
signal \N__53933\ : std_logic;
signal \N__53930\ : std_logic;
signal \N__53927\ : std_logic;
signal \N__53924\ : std_logic;
signal \N__53921\ : std_logic;
signal \N__53918\ : std_logic;
signal \N__53911\ : std_logic;
signal \N__53908\ : std_logic;
signal \N__53907\ : std_logic;
signal \N__53904\ : std_logic;
signal \N__53901\ : std_logic;
signal \N__53898\ : std_logic;
signal \N__53895\ : std_logic;
signal \N__53892\ : std_logic;
signal \N__53889\ : std_logic;
signal \N__53884\ : std_logic;
signal \N__53881\ : std_logic;
signal \N__53878\ : std_logic;
signal \N__53875\ : std_logic;
signal \N__53874\ : std_logic;
signal \N__53871\ : std_logic;
signal \N__53870\ : std_logic;
signal \N__53869\ : std_logic;
signal \N__53868\ : std_logic;
signal \N__53865\ : std_logic;
signal \N__53862\ : std_logic;
signal \N__53859\ : std_logic;
signal \N__53854\ : std_logic;
signal \N__53851\ : std_logic;
signal \N__53842\ : std_logic;
signal \N__53839\ : std_logic;
signal \N__53838\ : std_logic;
signal \N__53837\ : std_logic;
signal \N__53834\ : std_logic;
signal \N__53829\ : std_logic;
signal \N__53824\ : std_logic;
signal \N__53821\ : std_logic;
signal \N__53818\ : std_logic;
signal \N__53815\ : std_logic;
signal \N__53812\ : std_logic;
signal \N__53809\ : std_logic;
signal \N__53808\ : std_logic;
signal \N__53805\ : std_logic;
signal \N__53804\ : std_logic;
signal \N__53801\ : std_logic;
signal \N__53798\ : std_logic;
signal \N__53795\ : std_logic;
signal \N__53794\ : std_logic;
signal \N__53791\ : std_logic;
signal \N__53786\ : std_logic;
signal \N__53783\ : std_logic;
signal \N__53780\ : std_logic;
signal \N__53777\ : std_logic;
signal \N__53770\ : std_logic;
signal \N__53769\ : std_logic;
signal \N__53768\ : std_logic;
signal \N__53765\ : std_logic;
signal \N__53760\ : std_logic;
signal \N__53755\ : std_logic;
signal \N__53752\ : std_logic;
signal \N__53751\ : std_logic;
signal \N__53748\ : std_logic;
signal \N__53745\ : std_logic;
signal \N__53744\ : std_logic;
signal \N__53741\ : std_logic;
signal \N__53738\ : std_logic;
signal \N__53735\ : std_logic;
signal \N__53732\ : std_logic;
signal \N__53729\ : std_logic;
signal \N__53722\ : std_logic;
signal \N__53721\ : std_logic;
signal \N__53720\ : std_logic;
signal \N__53715\ : std_logic;
signal \N__53714\ : std_logic;
signal \N__53711\ : std_logic;
signal \N__53710\ : std_logic;
signal \N__53709\ : std_logic;
signal \N__53706\ : std_logic;
signal \N__53703\ : std_logic;
signal \N__53702\ : std_logic;
signal \N__53699\ : std_logic;
signal \N__53694\ : std_logic;
signal \N__53693\ : std_logic;
signal \N__53688\ : std_logic;
signal \N__53685\ : std_logic;
signal \N__53682\ : std_logic;
signal \N__53679\ : std_logic;
signal \N__53676\ : std_logic;
signal \N__53671\ : std_logic;
signal \N__53662\ : std_logic;
signal \N__53659\ : std_logic;
signal \N__53658\ : std_logic;
signal \N__53657\ : std_logic;
signal \N__53654\ : std_logic;
signal \N__53651\ : std_logic;
signal \N__53648\ : std_logic;
signal \N__53645\ : std_logic;
signal \N__53642\ : std_logic;
signal \N__53639\ : std_logic;
signal \N__53636\ : std_logic;
signal \N__53633\ : std_logic;
signal \N__53626\ : std_logic;
signal \N__53623\ : std_logic;
signal \N__53622\ : std_logic;
signal \N__53619\ : std_logic;
signal \N__53618\ : std_logic;
signal \N__53615\ : std_logic;
signal \N__53612\ : std_logic;
signal \N__53609\ : std_logic;
signal \N__53602\ : std_logic;
signal \N__53601\ : std_logic;
signal \N__53598\ : std_logic;
signal \N__53595\ : std_logic;
signal \N__53592\ : std_logic;
signal \N__53587\ : std_logic;
signal \N__53586\ : std_logic;
signal \N__53585\ : std_logic;
signal \N__53582\ : std_logic;
signal \N__53579\ : std_logic;
signal \N__53576\ : std_logic;
signal \N__53573\ : std_logic;
signal \N__53570\ : std_logic;
signal \N__53563\ : std_logic;
signal \N__53560\ : std_logic;
signal \N__53557\ : std_logic;
signal \N__53556\ : std_logic;
signal \N__53553\ : std_logic;
signal \N__53550\ : std_logic;
signal \N__53545\ : std_logic;
signal \N__53542\ : std_logic;
signal \N__53539\ : std_logic;
signal \N__53538\ : std_logic;
signal \N__53537\ : std_logic;
signal \N__53532\ : std_logic;
signal \N__53529\ : std_logic;
signal \N__53526\ : std_logic;
signal \N__53523\ : std_logic;
signal \N__53520\ : std_logic;
signal \N__53517\ : std_logic;
signal \N__53512\ : std_logic;
signal \N__53511\ : std_logic;
signal \N__53510\ : std_logic;
signal \N__53507\ : std_logic;
signal \N__53506\ : std_logic;
signal \N__53501\ : std_logic;
signal \N__53498\ : std_logic;
signal \N__53495\ : std_logic;
signal \N__53494\ : std_logic;
signal \N__53491\ : std_logic;
signal \N__53488\ : std_logic;
signal \N__53485\ : std_logic;
signal \N__53482\ : std_logic;
signal \N__53473\ : std_logic;
signal \N__53470\ : std_logic;
signal \N__53469\ : std_logic;
signal \N__53466\ : std_logic;
signal \N__53463\ : std_logic;
signal \N__53460\ : std_logic;
signal \N__53459\ : std_logic;
signal \N__53456\ : std_logic;
signal \N__53453\ : std_logic;
signal \N__53450\ : std_logic;
signal \N__53443\ : std_logic;
signal \N__53442\ : std_logic;
signal \N__53439\ : std_logic;
signal \N__53436\ : std_logic;
signal \N__53433\ : std_logic;
signal \N__53430\ : std_logic;
signal \N__53425\ : std_logic;
signal \N__53422\ : std_logic;
signal \N__53421\ : std_logic;
signal \N__53418\ : std_logic;
signal \N__53415\ : std_logic;
signal \N__53414\ : std_logic;
signal \N__53409\ : std_logic;
signal \N__53406\ : std_logic;
signal \N__53403\ : std_logic;
signal \N__53400\ : std_logic;
signal \N__53395\ : std_logic;
signal \N__53392\ : std_logic;
signal \N__53391\ : std_logic;
signal \N__53386\ : std_logic;
signal \N__53383\ : std_logic;
signal \N__53380\ : std_logic;
signal \N__53379\ : std_logic;
signal \N__53376\ : std_logic;
signal \N__53375\ : std_logic;
signal \N__53372\ : std_logic;
signal \N__53369\ : std_logic;
signal \N__53366\ : std_logic;
signal \N__53363\ : std_logic;
signal \N__53358\ : std_logic;
signal \N__53353\ : std_logic;
signal \N__53350\ : std_logic;
signal \N__53347\ : std_logic;
signal \N__53344\ : std_logic;
signal \N__53343\ : std_logic;
signal \N__53342\ : std_logic;
signal \N__53339\ : std_logic;
signal \N__53334\ : std_logic;
signal \N__53333\ : std_logic;
signal \N__53330\ : std_logic;
signal \N__53327\ : std_logic;
signal \N__53326\ : std_logic;
signal \N__53325\ : std_logic;
signal \N__53322\ : std_logic;
signal \N__53319\ : std_logic;
signal \N__53316\ : std_logic;
signal \N__53311\ : std_logic;
signal \N__53302\ : std_logic;
signal \N__53299\ : std_logic;
signal \N__53298\ : std_logic;
signal \N__53297\ : std_logic;
signal \N__53294\ : std_logic;
signal \N__53289\ : std_logic;
signal \N__53284\ : std_logic;
signal \N__53281\ : std_logic;
signal \N__53280\ : std_logic;
signal \N__53275\ : std_logic;
signal \N__53272\ : std_logic;
signal \N__53271\ : std_logic;
signal \N__53266\ : std_logic;
signal \N__53263\ : std_logic;
signal \N__53260\ : std_logic;
signal \N__53259\ : std_logic;
signal \N__53256\ : std_logic;
signal \N__53255\ : std_logic;
signal \N__53252\ : std_logic;
signal \N__53249\ : std_logic;
signal \N__53246\ : std_logic;
signal \N__53243\ : std_logic;
signal \N__53238\ : std_logic;
signal \N__53235\ : std_logic;
signal \N__53230\ : std_logic;
signal \N__53229\ : std_logic;
signal \N__53228\ : std_logic;
signal \N__53227\ : std_logic;
signal \N__53226\ : std_logic;
signal \N__53225\ : std_logic;
signal \N__53224\ : std_logic;
signal \N__53223\ : std_logic;
signal \N__53222\ : std_logic;
signal \N__53221\ : std_logic;
signal \N__53220\ : std_logic;
signal \N__53219\ : std_logic;
signal \N__53218\ : std_logic;
signal \N__53217\ : std_logic;
signal \N__53216\ : std_logic;
signal \N__53215\ : std_logic;
signal \N__53212\ : std_logic;
signal \N__53211\ : std_logic;
signal \N__53210\ : std_logic;
signal \N__53209\ : std_logic;
signal \N__53208\ : std_logic;
signal \N__53205\ : std_logic;
signal \N__53202\ : std_logic;
signal \N__53199\ : std_logic;
signal \N__53196\ : std_logic;
signal \N__53195\ : std_logic;
signal \N__53192\ : std_logic;
signal \N__53189\ : std_logic;
signal \N__53188\ : std_logic;
signal \N__53187\ : std_logic;
signal \N__53180\ : std_logic;
signal \N__53179\ : std_logic;
signal \N__53178\ : std_logic;
signal \N__53177\ : std_logic;
signal \N__53176\ : std_logic;
signal \N__53175\ : std_logic;
signal \N__53174\ : std_logic;
signal \N__53173\ : std_logic;
signal \N__53172\ : std_logic;
signal \N__53165\ : std_logic;
signal \N__53160\ : std_logic;
signal \N__53157\ : std_logic;
signal \N__53154\ : std_logic;
signal \N__53145\ : std_logic;
signal \N__53136\ : std_logic;
signal \N__53135\ : std_logic;
signal \N__53132\ : std_logic;
signal \N__53129\ : std_logic;
signal \N__53122\ : std_logic;
signal \N__53119\ : std_logic;
signal \N__53118\ : std_logic;
signal \N__53115\ : std_logic;
signal \N__53112\ : std_logic;
signal \N__53109\ : std_logic;
signal \N__53106\ : std_logic;
signal \N__53103\ : std_logic;
signal \N__53100\ : std_logic;
signal \N__53095\ : std_logic;
signal \N__53092\ : std_logic;
signal \N__53087\ : std_logic;
signal \N__53080\ : std_logic;
signal \N__53079\ : std_logic;
signal \N__53076\ : std_logic;
signal \N__53071\ : std_logic;
signal \N__53066\ : std_logic;
signal \N__53063\ : std_logic;
signal \N__53060\ : std_logic;
signal \N__53055\ : std_logic;
signal \N__53040\ : std_logic;
signal \N__53037\ : std_logic;
signal \N__53036\ : std_logic;
signal \N__53033\ : std_logic;
signal \N__53030\ : std_logic;
signal \N__53027\ : std_logic;
signal \N__53024\ : std_logic;
signal \N__53015\ : std_logic;
signal \N__53012\ : std_logic;
signal \N__53011\ : std_logic;
signal \N__53008\ : std_logic;
signal \N__53005\ : std_logic;
signal \N__53000\ : std_logic;
signal \N__52997\ : std_logic;
signal \N__52996\ : std_logic;
signal \N__52993\ : std_logic;
signal \N__52990\ : std_logic;
signal \N__52987\ : std_logic;
signal \N__52984\ : std_logic;
signal \N__52981\ : std_logic;
signal \N__52978\ : std_logic;
signal \N__52975\ : std_logic;
signal \N__52960\ : std_logic;
signal \N__52957\ : std_logic;
signal \N__52956\ : std_logic;
signal \N__52953\ : std_logic;
signal \N__52950\ : std_logic;
signal \N__52949\ : std_logic;
signal \N__52946\ : std_logic;
signal \N__52943\ : std_logic;
signal \N__52942\ : std_logic;
signal \N__52939\ : std_logic;
signal \N__52936\ : std_logic;
signal \N__52933\ : std_logic;
signal \N__52930\ : std_logic;
signal \N__52921\ : std_logic;
signal \N__52920\ : std_logic;
signal \N__52919\ : std_logic;
signal \N__52916\ : std_logic;
signal \N__52913\ : std_logic;
signal \N__52910\ : std_logic;
signal \N__52907\ : std_logic;
signal \N__52904\ : std_logic;
signal \N__52903\ : std_logic;
signal \N__52900\ : std_logic;
signal \N__52895\ : std_logic;
signal \N__52892\ : std_logic;
signal \N__52889\ : std_logic;
signal \N__52886\ : std_logic;
signal \N__52879\ : std_logic;
signal \N__52876\ : std_logic;
signal \N__52875\ : std_logic;
signal \N__52872\ : std_logic;
signal \N__52869\ : std_logic;
signal \N__52864\ : std_logic;
signal \N__52863\ : std_logic;
signal \N__52862\ : std_logic;
signal \N__52859\ : std_logic;
signal \N__52854\ : std_logic;
signal \N__52849\ : std_logic;
signal \N__52846\ : std_logic;
signal \N__52843\ : std_logic;
signal \N__52840\ : std_logic;
signal \N__52837\ : std_logic;
signal \N__52834\ : std_logic;
signal \N__52831\ : std_logic;
signal \N__52828\ : std_logic;
signal \N__52827\ : std_logic;
signal \N__52824\ : std_logic;
signal \N__52821\ : std_logic;
signal \N__52818\ : std_logic;
signal \N__52815\ : std_logic;
signal \N__52812\ : std_logic;
signal \N__52809\ : std_logic;
signal \N__52804\ : std_logic;
signal \N__52801\ : std_logic;
signal \N__52798\ : std_logic;
signal \N__52795\ : std_logic;
signal \N__52794\ : std_logic;
signal \N__52791\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52785\ : std_logic;
signal \N__52782\ : std_logic;
signal \N__52779\ : std_logic;
signal \N__52774\ : std_logic;
signal \N__52771\ : std_logic;
signal \N__52768\ : std_logic;
signal \N__52765\ : std_logic;
signal \N__52762\ : std_logic;
signal \N__52759\ : std_logic;
signal \N__52758\ : std_logic;
signal \N__52755\ : std_logic;
signal \N__52752\ : std_logic;
signal \N__52749\ : std_logic;
signal \N__52746\ : std_logic;
signal \N__52743\ : std_logic;
signal \N__52740\ : std_logic;
signal \N__52735\ : std_logic;
signal \N__52734\ : std_logic;
signal \N__52729\ : std_logic;
signal \N__52726\ : std_logic;
signal \N__52723\ : std_logic;
signal \N__52722\ : std_logic;
signal \N__52719\ : std_logic;
signal \N__52716\ : std_logic;
signal \N__52711\ : std_logic;
signal \N__52708\ : std_logic;
signal \N__52707\ : std_logic;
signal \N__52706\ : std_logic;
signal \N__52703\ : std_logic;
signal \N__52698\ : std_logic;
signal \N__52693\ : std_logic;
signal \N__52690\ : std_logic;
signal \N__52689\ : std_logic;
signal \N__52686\ : std_logic;
signal \N__52683\ : std_logic;
signal \N__52678\ : std_logic;
signal \N__52675\ : std_logic;
signal \N__52672\ : std_logic;
signal \N__52671\ : std_logic;
signal \N__52668\ : std_logic;
signal \N__52665\ : std_logic;
signal \N__52662\ : std_logic;
signal \N__52657\ : std_logic;
signal \N__52654\ : std_logic;
signal \N__52651\ : std_logic;
signal \N__52648\ : std_logic;
signal \N__52647\ : std_logic;
signal \N__52646\ : std_logic;
signal \N__52645\ : std_logic;
signal \N__52642\ : std_logic;
signal \N__52637\ : std_logic;
signal \N__52634\ : std_logic;
signal \N__52629\ : std_logic;
signal \N__52626\ : std_logic;
signal \N__52623\ : std_logic;
signal \N__52620\ : std_logic;
signal \N__52615\ : std_logic;
signal \N__52612\ : std_logic;
signal \N__52609\ : std_logic;
signal \N__52606\ : std_logic;
signal \N__52603\ : std_logic;
signal \N__52600\ : std_logic;
signal \N__52599\ : std_logic;
signal \N__52596\ : std_logic;
signal \N__52593\ : std_logic;
signal \N__52588\ : std_logic;
signal \N__52585\ : std_logic;
signal \N__52582\ : std_logic;
signal \N__52579\ : std_logic;
signal \N__52576\ : std_logic;
signal \N__52573\ : std_logic;
signal \N__52570\ : std_logic;
signal \N__52567\ : std_logic;
signal \N__52564\ : std_logic;
signal \N__52563\ : std_logic;
signal \N__52560\ : std_logic;
signal \N__52559\ : std_logic;
signal \N__52556\ : std_logic;
signal \N__52553\ : std_logic;
signal \N__52550\ : std_logic;
signal \N__52547\ : std_logic;
signal \N__52544\ : std_logic;
signal \N__52543\ : std_logic;
signal \N__52540\ : std_logic;
signal \N__52535\ : std_logic;
signal \N__52532\ : std_logic;
signal \N__52525\ : std_logic;
signal \N__52522\ : std_logic;
signal \N__52519\ : std_logic;
signal \N__52516\ : std_logic;
signal \N__52513\ : std_logic;
signal \N__52510\ : std_logic;
signal \N__52507\ : std_logic;
signal \N__52506\ : std_logic;
signal \N__52505\ : std_logic;
signal \N__52500\ : std_logic;
signal \N__52497\ : std_logic;
signal \N__52492\ : std_logic;
signal \N__52491\ : std_logic;
signal \N__52490\ : std_logic;
signal \N__52489\ : std_logic;
signal \N__52486\ : std_logic;
signal \N__52483\ : std_logic;
signal \N__52482\ : std_logic;
signal \N__52479\ : std_logic;
signal \N__52476\ : std_logic;
signal \N__52473\ : std_logic;
signal \N__52470\ : std_logic;
signal \N__52467\ : std_logic;
signal \N__52462\ : std_logic;
signal \N__52459\ : std_logic;
signal \N__52454\ : std_logic;
signal \N__52447\ : std_logic;
signal \N__52446\ : std_logic;
signal \N__52445\ : std_logic;
signal \N__52444\ : std_logic;
signal \N__52441\ : std_logic;
signal \N__52438\ : std_logic;
signal \N__52435\ : std_logic;
signal \N__52432\ : std_logic;
signal \N__52423\ : std_logic;
signal \N__52420\ : std_logic;
signal \N__52417\ : std_logic;
signal \N__52416\ : std_logic;
signal \N__52413\ : std_logic;
signal \N__52410\ : std_logic;
signal \N__52405\ : std_logic;
signal \N__52402\ : std_logic;
signal \N__52399\ : std_logic;
signal \N__52398\ : std_logic;
signal \N__52397\ : std_logic;
signal \N__52394\ : std_logic;
signal \N__52391\ : std_logic;
signal \N__52388\ : std_logic;
signal \N__52385\ : std_logic;
signal \N__52378\ : std_logic;
signal \N__52375\ : std_logic;
signal \N__52372\ : std_logic;
signal \N__52369\ : std_logic;
signal \N__52366\ : std_logic;
signal \N__52363\ : std_logic;
signal \N__52362\ : std_logic;
signal \N__52359\ : std_logic;
signal \N__52356\ : std_logic;
signal \N__52351\ : std_logic;
signal \N__52350\ : std_logic;
signal \N__52347\ : std_logic;
signal \N__52346\ : std_logic;
signal \N__52345\ : std_logic;
signal \N__52342\ : std_logic;
signal \N__52339\ : std_logic;
signal \N__52338\ : std_logic;
signal \N__52335\ : std_logic;
signal \N__52332\ : std_logic;
signal \N__52331\ : std_logic;
signal \N__52328\ : std_logic;
signal \N__52325\ : std_logic;
signal \N__52322\ : std_logic;
signal \N__52319\ : std_logic;
signal \N__52316\ : std_logic;
signal \N__52313\ : std_logic;
signal \N__52308\ : std_logic;
signal \N__52305\ : std_logic;
signal \N__52300\ : std_logic;
signal \N__52297\ : std_logic;
signal \N__52294\ : std_logic;
signal \N__52289\ : std_logic;
signal \N__52282\ : std_logic;
signal \N__52279\ : std_logic;
signal \N__52276\ : std_logic;
signal \N__52275\ : std_logic;
signal \N__52272\ : std_logic;
signal \N__52269\ : std_logic;
signal \N__52264\ : std_logic;
signal \N__52261\ : std_logic;
signal \N__52258\ : std_logic;
signal \N__52255\ : std_logic;
signal \N__52252\ : std_logic;
signal \N__52249\ : std_logic;
signal \N__52246\ : std_logic;
signal \N__52243\ : std_logic;
signal \N__52240\ : std_logic;
signal \N__52237\ : std_logic;
signal \N__52234\ : std_logic;
signal \N__52231\ : std_logic;
signal \N__52228\ : std_logic;
signal \N__52225\ : std_logic;
signal \N__52222\ : std_logic;
signal \N__52219\ : std_logic;
signal \N__52216\ : std_logic;
signal \N__52213\ : std_logic;
signal \N__52210\ : std_logic;
signal \N__52207\ : std_logic;
signal \N__52206\ : std_logic;
signal \N__52203\ : std_logic;
signal \N__52200\ : std_logic;
signal \N__52195\ : std_logic;
signal \N__52192\ : std_logic;
signal \N__52189\ : std_logic;
signal \N__52186\ : std_logic;
signal \N__52185\ : std_logic;
signal \N__52184\ : std_logic;
signal \N__52181\ : std_logic;
signal \N__52176\ : std_logic;
signal \N__52171\ : std_logic;
signal \N__52168\ : std_logic;
signal \N__52167\ : std_logic;
signal \N__52166\ : std_logic;
signal \N__52163\ : std_logic;
signal \N__52160\ : std_logic;
signal \N__52159\ : std_logic;
signal \N__52158\ : std_logic;
signal \N__52155\ : std_logic;
signal \N__52152\ : std_logic;
signal \N__52149\ : std_logic;
signal \N__52144\ : std_logic;
signal \N__52135\ : std_logic;
signal \N__52134\ : std_logic;
signal \N__52131\ : std_logic;
signal \N__52130\ : std_logic;
signal \N__52127\ : std_logic;
signal \N__52124\ : std_logic;
signal \N__52121\ : std_logic;
signal \N__52118\ : std_logic;
signal \N__52115\ : std_logic;
signal \N__52108\ : std_logic;
signal \N__52107\ : std_logic;
signal \N__52104\ : std_logic;
signal \N__52103\ : std_logic;
signal \N__52100\ : std_logic;
signal \N__52097\ : std_logic;
signal \N__52094\ : std_logic;
signal \N__52093\ : std_logic;
signal \N__52092\ : std_logic;
signal \N__52089\ : std_logic;
signal \N__52084\ : std_logic;
signal \N__52081\ : std_logic;
signal \N__52078\ : std_logic;
signal \N__52075\ : std_logic;
signal \N__52070\ : std_logic;
signal \N__52067\ : std_logic;
signal \N__52060\ : std_logic;
signal \N__52057\ : std_logic;
signal \N__52054\ : std_logic;
signal \N__52053\ : std_logic;
signal \N__52050\ : std_logic;
signal \N__52047\ : std_logic;
signal \N__52044\ : std_logic;
signal \N__52041\ : std_logic;
signal \N__52040\ : std_logic;
signal \N__52037\ : std_logic;
signal \N__52034\ : std_logic;
signal \N__52031\ : std_logic;
signal \N__52024\ : std_logic;
signal \N__52021\ : std_logic;
signal \N__52020\ : std_logic;
signal \N__52019\ : std_logic;
signal \N__52016\ : std_logic;
signal \N__52015\ : std_logic;
signal \N__52012\ : std_logic;
signal \N__52009\ : std_logic;
signal \N__52006\ : std_logic;
signal \N__52003\ : std_logic;
signal \N__52000\ : std_logic;
signal \N__51997\ : std_logic;
signal \N__51992\ : std_logic;
signal \N__51991\ : std_logic;
signal \N__51986\ : std_logic;
signal \N__51983\ : std_logic;
signal \N__51980\ : std_logic;
signal \N__51973\ : std_logic;
signal \N__51972\ : std_logic;
signal \N__51969\ : std_logic;
signal \N__51966\ : std_logic;
signal \N__51963\ : std_logic;
signal \N__51960\ : std_logic;
signal \N__51957\ : std_logic;
signal \N__51954\ : std_logic;
signal \N__51951\ : std_logic;
signal \N__51946\ : std_logic;
signal \N__51943\ : std_logic;
signal \N__51942\ : std_logic;
signal \N__51939\ : std_logic;
signal \N__51936\ : std_logic;
signal \N__51933\ : std_logic;
signal \N__51930\ : std_logic;
signal \N__51927\ : std_logic;
signal \N__51924\ : std_logic;
signal \N__51919\ : std_logic;
signal \N__51916\ : std_logic;
signal \N__51913\ : std_logic;
signal \N__51912\ : std_logic;
signal \N__51909\ : std_logic;
signal \N__51906\ : std_logic;
signal \N__51903\ : std_logic;
signal \N__51900\ : std_logic;
signal \N__51895\ : std_logic;
signal \N__51892\ : std_logic;
signal \N__51889\ : std_logic;
signal \N__51886\ : std_logic;
signal \N__51885\ : std_logic;
signal \N__51882\ : std_logic;
signal \N__51879\ : std_logic;
signal \N__51874\ : std_logic;
signal \N__51871\ : std_logic;
signal \N__51868\ : std_logic;
signal \N__51865\ : std_logic;
signal \N__51862\ : std_logic;
signal \N__51859\ : std_logic;
signal \N__51856\ : std_logic;
signal \N__51853\ : std_logic;
signal \N__51850\ : std_logic;
signal \N__51847\ : std_logic;
signal \N__51846\ : std_logic;
signal \N__51843\ : std_logic;
signal \N__51840\ : std_logic;
signal \N__51837\ : std_logic;
signal \N__51834\ : std_logic;
signal \N__51833\ : std_logic;
signal \N__51830\ : std_logic;
signal \N__51827\ : std_logic;
signal \N__51824\ : std_logic;
signal \N__51821\ : std_logic;
signal \N__51818\ : std_logic;
signal \N__51811\ : std_logic;
signal \N__51808\ : std_logic;
signal \N__51807\ : std_logic;
signal \N__51804\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51798\ : std_logic;
signal \N__51795\ : std_logic;
signal \N__51792\ : std_logic;
signal \N__51787\ : std_logic;
signal \N__51786\ : std_logic;
signal \N__51785\ : std_logic;
signal \N__51782\ : std_logic;
signal \N__51777\ : std_logic;
signal \N__51776\ : std_logic;
signal \N__51775\ : std_logic;
signal \N__51770\ : std_logic;
signal \N__51765\ : std_logic;
signal \N__51760\ : std_logic;
signal \N__51759\ : std_logic;
signal \N__51756\ : std_logic;
signal \N__51753\ : std_logic;
signal \N__51750\ : std_logic;
signal \N__51747\ : std_logic;
signal \N__51744\ : std_logic;
signal \N__51741\ : std_logic;
signal \N__51736\ : std_logic;
signal \N__51733\ : std_logic;
signal \N__51730\ : std_logic;
signal \N__51729\ : std_logic;
signal \N__51726\ : std_logic;
signal \N__51723\ : std_logic;
signal \N__51718\ : std_logic;
signal \N__51715\ : std_logic;
signal \N__51712\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51708\ : std_logic;
signal \N__51707\ : std_logic;
signal \N__51706\ : std_logic;
signal \N__51703\ : std_logic;
signal \N__51700\ : std_logic;
signal \N__51695\ : std_logic;
signal \N__51688\ : std_logic;
signal \N__51687\ : std_logic;
signal \N__51686\ : std_logic;
signal \N__51685\ : std_logic;
signal \N__51682\ : std_logic;
signal \N__51675\ : std_logic;
signal \N__51674\ : std_logic;
signal \N__51673\ : std_logic;
signal \N__51672\ : std_logic;
signal \N__51669\ : std_logic;
signal \N__51666\ : std_logic;
signal \N__51663\ : std_logic;
signal \N__51658\ : std_logic;
signal \N__51649\ : std_logic;
signal \N__51646\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51640\ : std_logic;
signal \N__51637\ : std_logic;
signal \N__51636\ : std_logic;
signal \N__51633\ : std_logic;
signal \N__51630\ : std_logic;
signal \N__51627\ : std_logic;
signal \N__51624\ : std_logic;
signal \N__51623\ : std_logic;
signal \N__51618\ : std_logic;
signal \N__51617\ : std_logic;
signal \N__51614\ : std_logic;
signal \N__51611\ : std_logic;
signal \N__51608\ : std_logic;
signal \N__51601\ : std_logic;
signal \N__51598\ : std_logic;
signal \N__51595\ : std_logic;
signal \N__51592\ : std_logic;
signal \N__51589\ : std_logic;
signal \N__51588\ : std_logic;
signal \N__51583\ : std_logic;
signal \N__51582\ : std_logic;
signal \N__51579\ : std_logic;
signal \N__51576\ : std_logic;
signal \N__51573\ : std_logic;
signal \N__51570\ : std_logic;
signal \N__51567\ : std_logic;
signal \N__51562\ : std_logic;
signal \N__51559\ : std_logic;
signal \N__51556\ : std_logic;
signal \N__51553\ : std_logic;
signal \N__51550\ : std_logic;
signal \N__51547\ : std_logic;
signal \N__51544\ : std_logic;
signal \N__51541\ : std_logic;
signal \N__51540\ : std_logic;
signal \N__51539\ : std_logic;
signal \N__51538\ : std_logic;
signal \N__51535\ : std_logic;
signal \N__51532\ : std_logic;
signal \N__51527\ : std_logic;
signal \N__51520\ : std_logic;
signal \N__51519\ : std_logic;
signal \N__51518\ : std_logic;
signal \N__51515\ : std_logic;
signal \N__51514\ : std_logic;
signal \N__51513\ : std_logic;
signal \N__51510\ : std_logic;
signal \N__51507\ : std_logic;
signal \N__51504\ : std_logic;
signal \N__51501\ : std_logic;
signal \N__51498\ : std_logic;
signal \N__51495\ : std_logic;
signal \N__51492\ : std_logic;
signal \N__51489\ : std_logic;
signal \N__51484\ : std_logic;
signal \N__51479\ : std_logic;
signal \N__51478\ : std_logic;
signal \N__51475\ : std_logic;
signal \N__51472\ : std_logic;
signal \N__51469\ : std_logic;
signal \N__51466\ : std_logic;
signal \N__51457\ : std_logic;
signal \N__51456\ : std_logic;
signal \N__51453\ : std_logic;
signal \N__51450\ : std_logic;
signal \N__51445\ : std_logic;
signal \N__51442\ : std_logic;
signal \N__51439\ : std_logic;
signal \N__51436\ : std_logic;
signal \N__51433\ : std_logic;
signal \N__51432\ : std_logic;
signal \N__51429\ : std_logic;
signal \N__51426\ : std_logic;
signal \N__51421\ : std_logic;
signal \N__51418\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51414\ : std_logic;
signal \N__51411\ : std_logic;
signal \N__51410\ : std_logic;
signal \N__51407\ : std_logic;
signal \N__51406\ : std_logic;
signal \N__51403\ : std_logic;
signal \N__51400\ : std_logic;
signal \N__51399\ : std_logic;
signal \N__51396\ : std_logic;
signal \N__51393\ : std_logic;
signal \N__51390\ : std_logic;
signal \N__51387\ : std_logic;
signal \N__51386\ : std_logic;
signal \N__51383\ : std_logic;
signal \N__51380\ : std_logic;
signal \N__51377\ : std_logic;
signal \N__51374\ : std_logic;
signal \N__51371\ : std_logic;
signal \N__51368\ : std_logic;
signal \N__51365\ : std_logic;
signal \N__51362\ : std_logic;
signal \N__51349\ : std_logic;
signal \N__51346\ : std_logic;
signal \N__51345\ : std_logic;
signal \N__51342\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51338\ : std_logic;
signal \N__51335\ : std_logic;
signal \N__51332\ : std_logic;
signal \N__51331\ : std_logic;
signal \N__51330\ : std_logic;
signal \N__51327\ : std_logic;
signal \N__51324\ : std_logic;
signal \N__51321\ : std_logic;
signal \N__51318\ : std_logic;
signal \N__51315\ : std_logic;
signal \N__51312\ : std_logic;
signal \N__51301\ : std_logic;
signal \N__51298\ : std_logic;
signal \N__51295\ : std_logic;
signal \N__51292\ : std_logic;
signal \N__51291\ : std_logic;
signal \N__51288\ : std_logic;
signal \N__51287\ : std_logic;
signal \N__51284\ : std_logic;
signal \N__51283\ : std_logic;
signal \N__51282\ : std_logic;
signal \N__51279\ : std_logic;
signal \N__51276\ : std_logic;
signal \N__51273\ : std_logic;
signal \N__51270\ : std_logic;
signal \N__51267\ : std_logic;
signal \N__51266\ : std_logic;
signal \N__51261\ : std_logic;
signal \N__51260\ : std_logic;
signal \N__51259\ : std_logic;
signal \N__51258\ : std_logic;
signal \N__51257\ : std_logic;
signal \N__51256\ : std_logic;
signal \N__51255\ : std_logic;
signal \N__51252\ : std_logic;
signal \N__51249\ : std_logic;
signal \N__51244\ : std_logic;
signal \N__51241\ : std_logic;
signal \N__51234\ : std_logic;
signal \N__51227\ : std_logic;
signal \N__51214\ : std_logic;
signal \N__51211\ : std_logic;
signal \N__51208\ : std_logic;
signal \N__51207\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51201\ : std_logic;
signal \N__51200\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51194\ : std_logic;
signal \N__51191\ : std_logic;
signal \N__51188\ : std_logic;
signal \N__51185\ : std_logic;
signal \N__51178\ : std_logic;
signal \N__51175\ : std_logic;
signal \N__51172\ : std_logic;
signal \N__51171\ : std_logic;
signal \N__51168\ : std_logic;
signal \N__51165\ : std_logic;
signal \N__51162\ : std_logic;
signal \N__51157\ : std_logic;
signal \N__51154\ : std_logic;
signal \N__51153\ : std_logic;
signal \N__51150\ : std_logic;
signal \N__51147\ : std_logic;
signal \N__51142\ : std_logic;
signal \N__51139\ : std_logic;
signal \N__51136\ : std_logic;
signal \N__51133\ : std_logic;
signal \N__51130\ : std_logic;
signal \N__51129\ : std_logic;
signal \N__51126\ : std_logic;
signal \N__51123\ : std_logic;
signal \N__51122\ : std_logic;
signal \N__51119\ : std_logic;
signal \N__51114\ : std_logic;
signal \N__51109\ : std_logic;
signal \N__51108\ : std_logic;
signal \N__51105\ : std_logic;
signal \N__51104\ : std_logic;
signal \N__51101\ : std_logic;
signal \N__51098\ : std_logic;
signal \N__51097\ : std_logic;
signal \N__51094\ : std_logic;
signal \N__51091\ : std_logic;
signal \N__51090\ : std_logic;
signal \N__51087\ : std_logic;
signal \N__51084\ : std_logic;
signal \N__51081\ : std_logic;
signal \N__51078\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51070\ : std_logic;
signal \N__51061\ : std_logic;
signal \N__51058\ : std_logic;
signal \N__51055\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51051\ : std_logic;
signal \N__51048\ : std_logic;
signal \N__51043\ : std_logic;
signal \N__51040\ : std_logic;
signal \N__51037\ : std_logic;
signal \N__51034\ : std_logic;
signal \N__51033\ : std_logic;
signal \N__51030\ : std_logic;
signal \N__51027\ : std_logic;
signal \N__51022\ : std_logic;
signal \N__51019\ : std_logic;
signal \N__51016\ : std_logic;
signal \N__51015\ : std_logic;
signal \N__51012\ : std_logic;
signal \N__51009\ : std_logic;
signal \N__51006\ : std_logic;
signal \N__51003\ : std_logic;
signal \N__51000\ : std_logic;
signal \N__50997\ : std_logic;
signal \N__50992\ : std_logic;
signal \N__50989\ : std_logic;
signal \N__50988\ : std_logic;
signal \N__50985\ : std_logic;
signal \N__50984\ : std_logic;
signal \N__50981\ : std_logic;
signal \N__50978\ : std_logic;
signal \N__50977\ : std_logic;
signal \N__50974\ : std_logic;
signal \N__50971\ : std_logic;
signal \N__50968\ : std_logic;
signal \N__50965\ : std_logic;
signal \N__50962\ : std_logic;
signal \N__50959\ : std_logic;
signal \N__50956\ : std_logic;
signal \N__50953\ : std_logic;
signal \N__50944\ : std_logic;
signal \N__50941\ : std_logic;
signal \N__50938\ : std_logic;
signal \N__50937\ : std_logic;
signal \N__50934\ : std_logic;
signal \N__50933\ : std_logic;
signal \N__50930\ : std_logic;
signal \N__50927\ : std_logic;
signal \N__50924\ : std_logic;
signal \N__50921\ : std_logic;
signal \N__50918\ : std_logic;
signal \N__50915\ : std_logic;
signal \N__50908\ : std_logic;
signal \N__50905\ : std_logic;
signal \N__50904\ : std_logic;
signal \N__50903\ : std_logic;
signal \N__50900\ : std_logic;
signal \N__50897\ : std_logic;
signal \N__50894\ : std_logic;
signal \N__50891\ : std_logic;
signal \N__50888\ : std_logic;
signal \N__50885\ : std_logic;
signal \N__50882\ : std_logic;
signal \N__50879\ : std_logic;
signal \N__50872\ : std_logic;
signal \N__50869\ : std_logic;
signal \N__50866\ : std_logic;
signal \N__50863\ : std_logic;
signal \N__50860\ : std_logic;
signal \N__50857\ : std_logic;
signal \N__50854\ : std_logic;
signal \N__50853\ : std_logic;
signal \N__50852\ : std_logic;
signal \N__50849\ : std_logic;
signal \N__50844\ : std_logic;
signal \N__50839\ : std_logic;
signal \N__50836\ : std_logic;
signal \N__50833\ : std_logic;
signal \N__50830\ : std_logic;
signal \N__50829\ : std_logic;
signal \N__50826\ : std_logic;
signal \N__50823\ : std_logic;
signal \N__50822\ : std_logic;
signal \N__50819\ : std_logic;
signal \N__50816\ : std_logic;
signal \N__50813\ : std_logic;
signal \N__50810\ : std_logic;
signal \N__50807\ : std_logic;
signal \N__50804\ : std_logic;
signal \N__50797\ : std_logic;
signal \N__50796\ : std_logic;
signal \N__50793\ : std_logic;
signal \N__50790\ : std_logic;
signal \N__50785\ : std_logic;
signal \N__50784\ : std_logic;
signal \N__50781\ : std_logic;
signal \N__50778\ : std_logic;
signal \N__50775\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50769\ : std_logic;
signal \N__50766\ : std_logic;
signal \N__50763\ : std_logic;
signal \N__50760\ : std_logic;
signal \N__50757\ : std_logic;
signal \N__50754\ : std_logic;
signal \N__50749\ : std_logic;
signal \N__50746\ : std_logic;
signal \N__50743\ : std_logic;
signal \N__50740\ : std_logic;
signal \N__50739\ : std_logic;
signal \N__50736\ : std_logic;
signal \N__50733\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50727\ : std_logic;
signal \N__50722\ : std_logic;
signal \N__50719\ : std_logic;
signal \N__50716\ : std_logic;
signal \N__50713\ : std_logic;
signal \N__50710\ : std_logic;
signal \N__50707\ : std_logic;
signal \N__50704\ : std_logic;
signal \N__50701\ : std_logic;
signal \N__50698\ : std_logic;
signal \N__50695\ : std_logic;
signal \N__50692\ : std_logic;
signal \N__50691\ : std_logic;
signal \N__50688\ : std_logic;
signal \N__50685\ : std_logic;
signal \N__50680\ : std_logic;
signal \N__50679\ : std_logic;
signal \N__50678\ : std_logic;
signal \N__50675\ : std_logic;
signal \N__50674\ : std_logic;
signal \N__50673\ : std_logic;
signal \N__50672\ : std_logic;
signal \N__50669\ : std_logic;
signal \N__50666\ : std_logic;
signal \N__50663\ : std_logic;
signal \N__50660\ : std_logic;
signal \N__50659\ : std_logic;
signal \N__50654\ : std_logic;
signal \N__50651\ : std_logic;
signal \N__50648\ : std_logic;
signal \N__50645\ : std_logic;
signal \N__50642\ : std_logic;
signal \N__50641\ : std_logic;
signal \N__50640\ : std_logic;
signal \N__50639\ : std_logic;
signal \N__50636\ : std_logic;
signal \N__50633\ : std_logic;
signal \N__50624\ : std_logic;
signal \N__50621\ : std_logic;
signal \N__50616\ : std_logic;
signal \N__50605\ : std_logic;
signal \N__50604\ : std_logic;
signal \N__50603\ : std_logic;
signal \N__50602\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50600\ : std_logic;
signal \N__50599\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50593\ : std_logic;
signal \N__50592\ : std_logic;
signal \N__50589\ : std_logic;
signal \N__50586\ : std_logic;
signal \N__50583\ : std_logic;
signal \N__50582\ : std_logic;
signal \N__50579\ : std_logic;
signal \N__50576\ : std_logic;
signal \N__50573\ : std_logic;
signal \N__50570\ : std_logic;
signal \N__50567\ : std_logic;
signal \N__50566\ : std_logic;
signal \N__50563\ : std_logic;
signal \N__50558\ : std_logic;
signal \N__50555\ : std_logic;
signal \N__50554\ : std_logic;
signal \N__50553\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50550\ : std_logic;
signal \N__50545\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50530\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50518\ : std_logic;
signal \N__50515\ : std_logic;
signal \N__50500\ : std_logic;
signal \N__50497\ : std_logic;
signal \N__50496\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50487\ : std_logic;
signal \N__50486\ : std_logic;
signal \N__50485\ : std_logic;
signal \N__50482\ : std_logic;
signal \N__50479\ : std_logic;
signal \N__50474\ : std_logic;
signal \N__50467\ : std_logic;
signal \N__50464\ : std_logic;
signal \N__50461\ : std_logic;
signal \N__50458\ : std_logic;
signal \N__50457\ : std_logic;
signal \N__50456\ : std_logic;
signal \N__50453\ : std_logic;
signal \N__50450\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50442\ : std_logic;
signal \N__50439\ : std_logic;
signal \N__50434\ : std_logic;
signal \N__50433\ : std_logic;
signal \N__50432\ : std_logic;
signal \N__50429\ : std_logic;
signal \N__50426\ : std_logic;
signal \N__50425\ : std_logic;
signal \N__50422\ : std_logic;
signal \N__50419\ : std_logic;
signal \N__50412\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50406\ : std_logic;
signal \N__50405\ : std_logic;
signal \N__50402\ : std_logic;
signal \N__50399\ : std_logic;
signal \N__50396\ : std_logic;
signal \N__50395\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50387\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50379\ : std_logic;
signal \N__50376\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50361\ : std_logic;
signal \N__50360\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50356\ : std_logic;
signal \N__50353\ : std_logic;
signal \N__50350\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50347\ : std_logic;
signal \N__50346\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50340\ : std_logic;
signal \N__50339\ : std_logic;
signal \N__50336\ : std_logic;
signal \N__50333\ : std_logic;
signal \N__50332\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50313\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50300\ : std_logic;
signal \N__50297\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50279\ : std_logic;
signal \N__50272\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50226\ : std_logic;
signal \N__50223\ : std_logic;
signal \N__50220\ : std_logic;
signal \N__50217\ : std_logic;
signal \N__50214\ : std_logic;
signal \N__50209\ : std_logic;
signal \N__50206\ : std_logic;
signal \N__50203\ : std_logic;
signal \N__50200\ : std_logic;
signal \N__50197\ : std_logic;
signal \N__50194\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50188\ : std_logic;
signal \N__50185\ : std_logic;
signal \N__50182\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50176\ : std_logic;
signal \N__50175\ : std_logic;
signal \N__50172\ : std_logic;
signal \N__50169\ : std_logic;
signal \N__50164\ : std_logic;
signal \N__50161\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50150\ : std_logic;
signal \N__50149\ : std_logic;
signal \N__50146\ : std_logic;
signal \N__50143\ : std_logic;
signal \N__50140\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50129\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__50123\ : std_logic;
signal \N__50120\ : std_logic;
signal \N__50113\ : std_logic;
signal \N__50110\ : std_logic;
signal \N__50109\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50105\ : std_logic;
signal \N__50102\ : std_logic;
signal \N__50099\ : std_logic;
signal \N__50092\ : std_logic;
signal \N__50089\ : std_logic;
signal \N__50086\ : std_logic;
signal \N__50083\ : std_logic;
signal \N__50082\ : std_logic;
signal \N__50081\ : std_logic;
signal \N__50078\ : std_logic;
signal \N__50077\ : std_logic;
signal \N__50076\ : std_logic;
signal \N__50073\ : std_logic;
signal \N__50070\ : std_logic;
signal \N__50067\ : std_logic;
signal \N__50064\ : std_logic;
signal \N__50063\ : std_logic;
signal \N__50060\ : std_logic;
signal \N__50057\ : std_logic;
signal \N__50054\ : std_logic;
signal \N__50049\ : std_logic;
signal \N__50046\ : std_logic;
signal \N__50043\ : std_logic;
signal \N__50038\ : std_logic;
signal \N__50033\ : std_logic;
signal \N__50026\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50022\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49995\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49984\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49980\ : std_logic;
signal \N__49979\ : std_logic;
signal \N__49976\ : std_logic;
signal \N__49975\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49968\ : std_logic;
signal \N__49965\ : std_logic;
signal \N__49960\ : std_logic;
signal \N__49951\ : std_logic;
signal \N__49948\ : std_logic;
signal \N__49945\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49933\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49927\ : std_logic;
signal \N__49924\ : std_logic;
signal \N__49921\ : std_logic;
signal \N__49918\ : std_logic;
signal \N__49917\ : std_logic;
signal \N__49916\ : std_logic;
signal \N__49913\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49907\ : std_logic;
signal \N__49906\ : std_logic;
signal \N__49903\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49886\ : std_logic;
signal \N__49879\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49869\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49863\ : std_logic;
signal \N__49858\ : std_logic;
signal \N__49855\ : std_logic;
signal \N__49852\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49844\ : std_logic;
signal \N__49841\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49828\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49822\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49816\ : std_logic;
signal \N__49813\ : std_logic;
signal \N__49810\ : std_logic;
signal \N__49809\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49802\ : std_logic;
signal \N__49799\ : std_logic;
signal \N__49794\ : std_logic;
signal \N__49789\ : std_logic;
signal \N__49786\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49781\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49775\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49765\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49754\ : std_logic;
signal \N__49751\ : std_logic;
signal \N__49748\ : std_logic;
signal \N__49745\ : std_logic;
signal \N__49744\ : std_logic;
signal \N__49741\ : std_logic;
signal \N__49738\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49731\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49717\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49696\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49692\ : std_logic;
signal \N__49691\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49683\ : std_logic;
signal \N__49678\ : std_logic;
signal \N__49677\ : std_logic;
signal \N__49676\ : std_logic;
signal \N__49673\ : std_logic;
signal \N__49672\ : std_logic;
signal \N__49669\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49665\ : std_logic;
signal \N__49662\ : std_logic;
signal \N__49659\ : std_logic;
signal \N__49656\ : std_logic;
signal \N__49655\ : std_logic;
signal \N__49652\ : std_logic;
signal \N__49649\ : std_logic;
signal \N__49644\ : std_logic;
signal \N__49641\ : std_logic;
signal \N__49638\ : std_logic;
signal \N__49633\ : std_logic;
signal \N__49630\ : std_logic;
signal \N__49627\ : std_logic;
signal \N__49624\ : std_logic;
signal \N__49619\ : std_logic;
signal \N__49618\ : std_logic;
signal \N__49615\ : std_logic;
signal \N__49612\ : std_logic;
signal \N__49609\ : std_logic;
signal \N__49606\ : std_logic;
signal \N__49597\ : std_logic;
signal \N__49594\ : std_logic;
signal \N__49591\ : std_logic;
signal \N__49588\ : std_logic;
signal \N__49585\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49581\ : std_logic;
signal \N__49578\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49571\ : std_logic;
signal \N__49566\ : std_logic;
signal \N__49563\ : std_logic;
signal \N__49560\ : std_logic;
signal \N__49559\ : std_logic;
signal \N__49558\ : std_logic;
signal \N__49553\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49540\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49535\ : std_logic;
signal \N__49532\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49522\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49516\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49510\ : std_logic;
signal \N__49507\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49502\ : std_logic;
signal \N__49499\ : std_logic;
signal \N__49498\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49492\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49487\ : std_logic;
signal \N__49484\ : std_logic;
signal \N__49479\ : std_logic;
signal \N__49476\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49458\ : std_logic;
signal \N__49455\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49448\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49441\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49401\ : std_logic;
signal \N__49398\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49396\ : std_logic;
signal \N__49393\ : std_logic;
signal \N__49390\ : std_logic;
signal \N__49387\ : std_logic;
signal \N__49384\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49371\ : std_logic;
signal \N__49368\ : std_logic;
signal \N__49365\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49357\ : std_logic;
signal \N__49354\ : std_logic;
signal \N__49351\ : std_logic;
signal \N__49348\ : std_logic;
signal \N__49347\ : std_logic;
signal \N__49346\ : std_logic;
signal \N__49343\ : std_logic;
signal \N__49340\ : std_logic;
signal \N__49337\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49329\ : std_logic;
signal \N__49328\ : std_logic;
signal \N__49327\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49320\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49312\ : std_logic;
signal \N__49303\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49301\ : std_logic;
signal \N__49298\ : std_logic;
signal \N__49295\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49288\ : std_logic;
signal \N__49285\ : std_logic;
signal \N__49282\ : std_logic;
signal \N__49279\ : std_logic;
signal \N__49276\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49266\ : std_logic;
signal \N__49261\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49259\ : std_logic;
signal \N__49258\ : std_logic;
signal \N__49257\ : std_logic;
signal \N__49252\ : std_logic;
signal \N__49249\ : std_logic;
signal \N__49246\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49240\ : std_logic;
signal \N__49231\ : std_logic;
signal \N__49230\ : std_logic;
signal \N__49229\ : std_logic;
signal \N__49228\ : std_logic;
signal \N__49227\ : std_logic;
signal \N__49222\ : std_logic;
signal \N__49219\ : std_logic;
signal \N__49214\ : std_logic;
signal \N__49213\ : std_logic;
signal \N__49210\ : std_logic;
signal \N__49205\ : std_logic;
signal \N__49202\ : std_logic;
signal \N__49199\ : std_logic;
signal \N__49196\ : std_logic;
signal \N__49193\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49183\ : std_logic;
signal \N__49182\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49178\ : std_logic;
signal \N__49175\ : std_logic;
signal \N__49172\ : std_logic;
signal \N__49169\ : std_logic;
signal \N__49166\ : std_logic;
signal \N__49161\ : std_logic;
signal \N__49160\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49152\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49136\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49127\ : std_logic;
signal \N__49124\ : std_logic;
signal \N__49121\ : std_logic;
signal \N__49118\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49098\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49092\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49084\ : std_logic;
signal \N__49081\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49079\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49073\ : std_logic;
signal \N__49070\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49068\ : std_logic;
signal \N__49065\ : std_logic;
signal \N__49062\ : std_logic;
signal \N__49059\ : std_logic;
signal \N__49056\ : std_logic;
signal \N__49053\ : std_logic;
signal \N__49050\ : std_logic;
signal \N__49045\ : std_logic;
signal \N__49040\ : std_logic;
signal \N__49037\ : std_logic;
signal \N__49034\ : std_logic;
signal \N__49031\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49017\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49011\ : std_logic;
signal \N__49006\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48997\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48985\ : std_logic;
signal \N__48982\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48973\ : std_logic;
signal \N__48970\ : std_logic;
signal \N__48967\ : std_logic;
signal \N__48964\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48960\ : std_logic;
signal \N__48957\ : std_logic;
signal \N__48954\ : std_logic;
signal \N__48949\ : std_logic;
signal \N__48946\ : std_logic;
signal \N__48943\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48934\ : std_logic;
signal \N__48933\ : std_logic;
signal \N__48932\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48930\ : std_logic;
signal \N__48927\ : std_logic;
signal \N__48924\ : std_logic;
signal \N__48921\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48907\ : std_logic;
signal \N__48904\ : std_logic;
signal \N__48901\ : std_logic;
signal \N__48898\ : std_logic;
signal \N__48895\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48885\ : std_logic;
signal \N__48880\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48873\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48869\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48860\ : std_logic;
signal \N__48855\ : std_logic;
signal \N__48852\ : std_logic;
signal \N__48849\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48838\ : std_logic;
signal \N__48837\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48831\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48829\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48823\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48814\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48808\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48799\ : std_logic;
signal \N__48790\ : std_logic;
signal \N__48789\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48785\ : std_logic;
signal \N__48782\ : std_logic;
signal \N__48779\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48772\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48757\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48730\ : std_logic;
signal \N__48727\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48711\ : std_logic;
signal \N__48708\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48694\ : std_logic;
signal \N__48691\ : std_logic;
signal \N__48688\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48679\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48661\ : std_logic;
signal \N__48658\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48650\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48644\ : std_logic;
signal \N__48641\ : std_logic;
signal \N__48634\ : std_logic;
signal \N__48631\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48618\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48605\ : std_logic;
signal \N__48602\ : std_logic;
signal \N__48599\ : std_logic;
signal \N__48596\ : std_logic;
signal \N__48595\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48584\ : std_logic;
signal \N__48581\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48553\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48541\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48531\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48524\ : std_logic;
signal \N__48521\ : std_logic;
signal \N__48518\ : std_logic;
signal \N__48511\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48496\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48490\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48477\ : std_logic;
signal \N__48474\ : std_logic;
signal \N__48471\ : std_logic;
signal \N__48468\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48444\ : std_logic;
signal \N__48441\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48423\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48391\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48382\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48377\ : std_logic;
signal \N__48374\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48366\ : std_logic;
signal \N__48363\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48327\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48319\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48311\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48301\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48248\ : std_logic;
signal \N__48243\ : std_logic;
signal \N__48240\ : std_logic;
signal \N__48237\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48219\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48192\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48184\ : std_logic;
signal \N__48181\ : std_logic;
signal \N__48178\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48145\ : std_logic;
signal \N__48142\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48136\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48127\ : std_logic;
signal \N__48120\ : std_logic;
signal \N__48117\ : std_logic;
signal \N__48114\ : std_logic;
signal \N__48111\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48102\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48082\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48068\ : std_logic;
signal \N__48065\ : std_logic;
signal \N__48062\ : std_logic;
signal \N__48059\ : std_logic;
signal \N__48052\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48046\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48040\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48034\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48015\ : std_logic;
signal \N__48012\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__48001\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47980\ : std_logic;
signal \N__47977\ : std_logic;
signal \N__47976\ : std_logic;
signal \N__47975\ : std_logic;
signal \N__47972\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47953\ : std_logic;
signal \N__47950\ : std_logic;
signal \N__47947\ : std_logic;
signal \N__47944\ : std_logic;
signal \N__47941\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47935\ : std_logic;
signal \N__47932\ : std_logic;
signal \N__47929\ : std_logic;
signal \N__47926\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47900\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47845\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47812\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47773\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47767\ : std_logic;
signal \N__47764\ : std_logic;
signal \N__47761\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47755\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47749\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47739\ : std_logic;
signal \N__47734\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47709\ : std_logic;
signal \N__47704\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47670\ : std_logic;
signal \N__47667\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47646\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47623\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47614\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47597\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47593\ : std_logic;
signal \N__47588\ : std_logic;
signal \N__47585\ : std_logic;
signal \N__47582\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47560\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47552\ : std_logic;
signal \N__47549\ : std_logic;
signal \N__47548\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47539\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47526\ : std_logic;
signal \N__47521\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47491\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47479\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47467\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47370\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47266\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47239\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47216\ : std_logic;
signal \N__47213\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47207\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47205\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47192\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47176\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47170\ : std_logic;
signal \N__47167\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47161\ : std_logic;
signal \N__47158\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47145\ : std_logic;
signal \N__47142\ : std_logic;
signal \N__47139\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47125\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47104\ : std_logic;
signal \N__47101\ : std_logic;
signal \N__47098\ : std_logic;
signal \N__47095\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47086\ : std_logic;
signal \N__47083\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47079\ : std_logic;
signal \N__47076\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47065\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47059\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47046\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47038\ : std_logic;
signal \N__47035\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47032\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47026\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47010\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46984\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46954\ : std_logic;
signal \N__46951\ : std_logic;
signal \N__46948\ : std_logic;
signal \N__46945\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46938\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46933\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46865\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46803\ : std_logic;
signal \N__46800\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46797\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46756\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46739\ : std_logic;
signal \N__46738\ : std_logic;
signal \N__46737\ : std_logic;
signal \N__46736\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46732\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46730\ : std_logic;
signal \N__46729\ : std_logic;
signal \N__46728\ : std_logic;
signal \N__46727\ : std_logic;
signal \N__46726\ : std_logic;
signal \N__46725\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46704\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46692\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46645\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46636\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46582\ : std_logic;
signal \N__46577\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46569\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46505\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46495\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46473\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46368\ : std_logic;
signal \N__46365\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46338\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46334\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46330\ : std_logic;
signal \N__46327\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46283\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46266\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46262\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46251\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46241\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46207\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46203\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46167\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46138\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45985\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45969\ : std_logic;
signal \N__45966\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45880\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45868\ : std_logic;
signal \N__45865\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45853\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45847\ : std_logic;
signal \N__45844\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45829\ : std_logic;
signal \N__45826\ : std_logic;
signal \N__45825\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45814\ : std_logic;
signal \N__45811\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45793\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45780\ : std_logic;
signal \N__45777\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45766\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45738\ : std_logic;
signal \N__45733\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45713\ : std_logic;
signal \N__45710\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45703\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45685\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45660\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45612\ : std_logic;
signal \N__45609\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45565\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45509\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45475\ : std_logic;
signal \N__45472\ : std_logic;
signal \N__45469\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45379\ : std_logic;
signal \N__45376\ : std_logic;
signal \N__45373\ : std_logic;
signal \N__45370\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45334\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45326\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45316\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45307\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45291\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45287\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45274\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45259\ : std_logic;
signal \N__45256\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45217\ : std_logic;
signal \N__45214\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45199\ : std_logic;
signal \N__45196\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45189\ : std_logic;
signal \N__45188\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45179\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45170\ : std_logic;
signal \N__45163\ : std_logic;
signal \N__45154\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45142\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45124\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44996\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44945\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44897\ : std_logic;
signal \N__44894\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44855\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44809\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44804\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44795\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44782\ : std_logic;
signal \N__44779\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44752\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44743\ : std_logic;
signal \N__44740\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44704\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44693\ : std_logic;
signal \N__44690\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44681\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44668\ : std_logic;
signal \N__44665\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44651\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44638\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44634\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44616\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44571\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44562\ : std_logic;
signal \N__44559\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44538\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44524\ : std_logic;
signal \N__44521\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44511\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44472\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44413\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44384\ : std_logic;
signal \N__44383\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44344\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44287\ : std_logic;
signal \N__44284\ : std_logic;
signal \N__44281\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44240\ : std_logic;
signal \N__44237\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44215\ : std_logic;
signal \N__44212\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44137\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44125\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44117\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44048\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44030\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44005\ : std_logic;
signal \N__44002\ : std_logic;
signal \N__43999\ : std_logic;
signal \N__43996\ : std_logic;
signal \N__43993\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43975\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43972\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43961\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43942\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43918\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43912\ : std_logic;
signal \N__43909\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43906\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43883\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43877\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43802\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43791\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43783\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43738\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43695\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43674\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43659\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43627\ : std_logic;
signal \N__43624\ : std_logic;
signal \N__43621\ : std_logic;
signal \N__43618\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43551\ : std_logic;
signal \N__43548\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43541\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43531\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43522\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43503\ : std_logic;
signal \N__43498\ : std_logic;
signal \N__43495\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43454\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43434\ : std_logic;
signal \N__43431\ : std_logic;
signal \N__43428\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43404\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43389\ : std_logic;
signal \N__43386\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43326\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43247\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43234\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43207\ : std_logic;
signal \N__43204\ : std_logic;
signal \N__43201\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43195\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43137\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43084\ : std_logic;
signal \N__43081\ : std_logic;
signal \N__43078\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43057\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43045\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43015\ : std_logic;
signal \N__43012\ : std_logic;
signal \N__43009\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42901\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42868\ : std_logic;
signal \N__42865\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42802\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42756\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42750\ : std_logic;
signal \N__42747\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42700\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42676\ : std_logic;
signal \N__42673\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42668\ : std_logic;
signal \N__42665\ : std_logic;
signal \N__42662\ : std_logic;
signal \N__42659\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42599\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42586\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42565\ : std_logic;
signal \N__42562\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42547\ : std_logic;
signal \N__42544\ : std_logic;
signal \N__42541\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42536\ : std_logic;
signal \N__42533\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42520\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42506\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42497\ : std_logic;
signal \N__42496\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42479\ : std_logic;
signal \N__42476\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42464\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42427\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42418\ : std_logic;
signal \N__42415\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42361\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42355\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42349\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42343\ : std_logic;
signal \N__42338\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42329\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42251\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42210\ : std_logic;
signal \N__42207\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42178\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42142\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42133\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42127\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42121\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42085\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41977\ : std_logic;
signal \N__41974\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41971\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41965\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41942\ : std_logic;
signal \N__41939\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41929\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41926\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41915\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41878\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41830\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41823\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41776\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41761\ : std_logic;
signal \N__41758\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41725\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41721\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41710\ : std_logic;
signal \N__41707\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41677\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41659\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41644\ : std_logic;
signal \N__41641\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41632\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41533\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41518\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41486\ : std_logic;
signal \N__41483\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41460\ : std_logic;
signal \N__41459\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41456\ : std_logic;
signal \N__41453\ : std_logic;
signal \N__41450\ : std_logic;
signal \N__41449\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41404\ : std_logic;
signal \N__41403\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41384\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41352\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41310\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41236\ : std_logic;
signal \N__41233\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41216\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41176\ : std_logic;
signal \N__41173\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41155\ : std_logic;
signal \N__41152\ : std_logic;
signal \N__41149\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41131\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41110\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41080\ : std_logic;
signal \N__41077\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41029\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41027\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40972\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40963\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40927\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40904\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40897\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40883\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40826\ : std_logic;
signal \N__40825\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40823\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40554\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40286\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40187\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40165\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40149\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40137\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40071\ : std_logic;
signal \N__40068\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40062\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40026\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39955\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39934\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39913\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39868\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39865\ : std_logic;
signal \N__39862\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39740\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39487\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39409\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39250\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39194\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38997\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38695\ : std_logic;
signal \N__38692\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38663\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38362\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38354\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37799\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37684\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37182\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37056\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37023\ : std_logic;
signal \N__37020\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36730\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36493\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36424\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36373\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35263\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal tx_enable : std_logic;
signal \LED_c\ : std_logic;
signal \c0.n18673\ : std_logic;
signal \c0.n18661\ : std_logic;
signal n39 : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \quad_counter0.n17222\ : std_logic;
signal \quad_counter0.n17223\ : std_logic;
signal \quad_counter0.n17224\ : std_logic;
signal \quad_counter0.n17225\ : std_logic;
signal \quad_counter0.n17226\ : std_logic;
signal \quad_counter0.n17227\ : std_logic;
signal \quad_counter0.n17228\ : std_logic;
signal \quad_counter0.n17229\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \quad_counter0.n17230\ : std_logic;
signal \quad_counter0.n17231\ : std_logic;
signal \quad_counter0.n17232\ : std_logic;
signal \quad_counter0.n17233\ : std_logic;
signal \quad_counter0.n17234\ : std_logic;
signal \quad_counter0.n17235\ : std_logic;
signal \quad_counter0.n17236\ : std_logic;
signal data_out_frame_6_6 : std_logic;
signal data_out_frame_5_1 : std_logic;
signal data_out_frame_7_6 : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \quad_counter0.b_delay_counter_1\ : std_logic;
signal \quad_counter0.n13182\ : std_logic;
signal \quad_counter0.n17207\ : std_logic;
signal \quad_counter0.n17208\ : std_logic;
signal \quad_counter0.n17209\ : std_logic;
signal \quad_counter0.b_delay_counter_4\ : std_logic;
signal \quad_counter0.n13197\ : std_logic;
signal \quad_counter0.n17210\ : std_logic;
signal \quad_counter0.n17211\ : std_logic;
signal \quad_counter0.n17212\ : std_logic;
signal \quad_counter0.b_delay_counter_7\ : std_logic;
signal \quad_counter0.n13214\ : std_logic;
signal \quad_counter0.n17213\ : std_logic;
signal \quad_counter0.n17214\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \quad_counter0.n17215\ : std_logic;
signal \quad_counter0.n17216\ : std_logic;
signal \quad_counter0.b_delay_counter_11\ : std_logic;
signal \quad_counter0.n13257\ : std_logic;
signal \quad_counter0.n17217\ : std_logic;
signal \quad_counter0.n17218\ : std_logic;
signal \quad_counter0.b_delay_counter_13\ : std_logic;
signal \quad_counter0.n13263\ : std_logic;
signal \quad_counter0.n17219\ : std_logic;
signal \quad_counter0.n17220\ : std_logic;
signal \quad_counter0.n17221\ : std_logic;
signal \quad_counter0.n13260\ : std_logic;
signal \quad_counter0.b_delay_counter_12\ : std_logic;
signal \quad_counter0.n13444\ : std_logic;
signal \quad_counter0.n13266\ : std_logic;
signal \quad_counter0.b_delay_counter_14\ : std_logic;
signal \quad_counter0.n13248\ : std_logic;
signal \quad_counter0.b_delay_counter_8\ : std_logic;
signal \quad_counter0.n13203\ : std_logic;
signal \quad_counter0.b_delay_counter_6\ : std_logic;
signal \quad_counter0.b_delay_counter_0\ : std_logic;
signal \quad_counter0.n13251\ : std_logic;
signal \quad_counter0.b_delay_counter_9\ : std_logic;
signal \quad_counter0.n13194\ : std_logic;
signal \quad_counter0.b_delay_counter_3\ : std_logic;
signal \quad_counter0.n13200\ : std_logic;
signal \quad_counter0.b_delay_counter_5\ : std_logic;
signal \c0.n18649\ : std_logic;
signal \c0.n18639\ : std_logic;
signal \c0.n18663\ : std_logic;
signal \a_delay_counter_15__N_2916\ : std_logic;
signal n12447 : std_logic;
signal \PIN_7_c\ : std_logic;
signal \quadA_delayed\ : std_logic;
signal \quad_counter0.a_delay_counter_15\ : std_logic;
signal \quad_counter0.a_delay_counter_8\ : std_logic;
signal \quad_counter0.a_delay_counter_1\ : std_logic;
signal \quad_counter0.a_delay_counter_6\ : std_logic;
signal \quad_counter0.a_delay_counter_9\ : std_logic;
signal \quad_counter0.a_delay_counter_7\ : std_logic;
signal \quad_counter0.n18_cascade_\ : std_logic;
signal a_delay_counter_0 : std_logic;
signal \quad_counter0.n20_cascade_\ : std_logic;
signal \quad_counter0.a_delay_counter_2\ : std_logic;
signal n11349 : std_logic;
signal \quad_counter0.a_delay_counter_5\ : std_logic;
signal \quad_counter0.a_delay_counter_10\ : std_logic;
signal \quad_counter0.a_delay_counter_12\ : std_logic;
signal \quad_counter0.a_delay_counter_3\ : std_logic;
signal \quad_counter0.n20954\ : std_logic;
signal \quad_counter0.a_delay_counter_4\ : std_logic;
signal \quad_counter0.a_delay_counter_11\ : std_logic;
signal \quad_counter0.a_delay_counter_14\ : std_logic;
signal \quad_counter0.a_delay_counter_13\ : std_logic;
signal \quad_counter0.n19\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \quad_counter0.count_direction\ : std_logic;
signal n2279 : std_logic;
signal \quad_counter0.n17282\ : std_logic;
signal n2278 : std_logic;
signal \quad_counter0.n17283\ : std_logic;
signal encoder0_position_2 : std_logic;
signal n2277 : std_logic;
signal \quad_counter0.n17284\ : std_logic;
signal encoder0_position_3 : std_logic;
signal n2276 : std_logic;
signal \quad_counter0.n17285\ : std_logic;
signal \quad_counter0.n17286\ : std_logic;
signal \quad_counter0.n17287\ : std_logic;
signal \quad_counter0.n17288\ : std_logic;
signal \quad_counter0.n17289\ : std_logic;
signal \bfn_10_10_0_\ : std_logic;
signal \quad_counter0.n17290\ : std_logic;
signal \quad_counter0.n17291\ : std_logic;
signal \quad_counter0.n17292\ : std_logic;
signal \quad_counter0.n17293\ : std_logic;
signal \quad_counter0.n17294\ : std_logic;
signal \quad_counter0.n17295\ : std_logic;
signal \quad_counter0.n17296\ : std_logic;
signal \quad_counter0.n17297\ : std_logic;
signal \bfn_10_11_0_\ : std_logic;
signal \quad_counter0.n17298\ : std_logic;
signal \quad_counter0.n17299\ : std_logic;
signal n2261 : std_logic;
signal \quad_counter0.n17300\ : std_logic;
signal n2260 : std_logic;
signal \quad_counter0.n17301\ : std_logic;
signal n2259 : std_logic;
signal \quad_counter0.n17302\ : std_logic;
signal n2258 : std_logic;
signal \quad_counter0.n17303\ : std_logic;
signal encoder0_position_22 : std_logic;
signal n2257 : std_logic;
signal \quad_counter0.n17304\ : std_logic;
signal \quad_counter0.n17305\ : std_logic;
signal n2256 : std_logic;
signal \bfn_10_12_0_\ : std_logic;
signal n2255 : std_logic;
signal \quad_counter0.n17306\ : std_logic;
signal n2254 : std_logic;
signal \quad_counter0.n17307\ : std_logic;
signal \quad_counter0.n17308\ : std_logic;
signal \quad_counter0.n17309\ : std_logic;
signal \quad_counter0.n17310\ : std_logic;
signal \quad_counter0.n17311\ : std_logic;
signal \quad_counter0.n17312\ : std_logic;
signal \quad_counter0.n17313\ : std_logic;
signal \quad_counter0.n2228\ : std_logic;
signal \bfn_10_13_0_\ : std_logic;
signal n2275 : std_logic;
signal n2272 : std_logic;
signal n2274 : std_logic;
signal n2248 : std_logic;
signal \c0.n5_adj_3471\ : std_logic;
signal encoder0_position_5 : std_logic;
signal data_out_frame_9_6 : std_logic;
signal \quad_counter0.n13254\ : std_logic;
signal \quad_counter0.b_delay_counter_10\ : std_logic;
signal \quad_counter0.n13269\ : std_logic;
signal \quad_counter0.b_delay_counter_15\ : std_logic;
signal \quad_counter0.n26_adj_2991\ : std_logic;
signal \quad_counter0.n27_adj_2992\ : std_logic;
signal \quad_counter0.n28_adj_2990\ : std_logic;
signal \quad_counter0.n25_adj_2993\ : std_logic;
signal n11347 : std_logic;
signal \n11347_cascade_\ : std_logic;
signal \quad_counter0.n21603\ : std_logic;
signal data_out_frame_10_6 : std_logic;
signal \c0.n21629\ : std_logic;
signal \PIN_8_c\ : std_logic;
signal \quadB_delayed\ : std_logic;
signal \quad_counter0.n13187\ : std_logic;
signal \quad_counter0.b_delay_counter_2\ : std_logic;
signal \c0.n21331_cascade_\ : std_logic;
signal \c0.n17354_cascade_\ : std_logic;
signal \c0.n21521\ : std_logic;
signal \c0.tx.n6_cascade_\ : std_logic;
signal \c0.n15938_cascade_\ : std_logic;
signal \c0.tx.r_Clock_Count_0\ : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \c0.tx.r_Clock_Count_1\ : std_logic;
signal \c0.tx.n17274\ : std_logic;
signal \c0.tx.r_Clock_Count_2\ : std_logic;
signal \c0.tx.n17275\ : std_logic;
signal \c0.tx.r_Clock_Count_3\ : std_logic;
signal \c0.tx.n17276\ : std_logic;
signal \c0.tx.r_Clock_Count_4\ : std_logic;
signal \c0.tx.n17277\ : std_logic;
signal \c0.tx.r_Clock_Count_5\ : std_logic;
signal \c0.tx.n17278\ : std_logic;
signal \c0.tx.r_Clock_Count_6\ : std_logic;
signal \c0.tx.n17279\ : std_logic;
signal \c0.tx.r_Clock_Count_7\ : std_logic;
signal \c0.tx.n17280\ : std_logic;
signal \c0.tx.n17281\ : std_logic;
signal \bfn_10_19_0_\ : std_logic;
signal \c0.n18671\ : std_logic;
signal \c0.n18617\ : std_logic;
signal \quad_counter1.n25_adj_3577_cascade_\ : std_logic;
signal \n11343_cascade_\ : std_logic;
signal \n12417_cascade_\ : std_logic;
signal \quad_counter1.n28_adj_3574\ : std_logic;
signal \PIN_13_c\ : std_logic;
signal n11343 : std_logic;
signal \quadB_delayed_adj_3585\ : std_logic;
signal \quad_counter1.n26_adj_3575\ : std_logic;
signal \quad_counter1.n27_adj_3576\ : std_logic;
signal \quad_counter1.n16_cascade_\ : std_logic;
signal \quad_counter1.n24_adj_3578_cascade_\ : std_logic;
signal n11351 : std_logic;
signal \B_filtered\ : std_logic;
signal \quad_counter0.B_delayed\ : std_logic;
signal \quad_counter1.n6\ : std_logic;
signal \A_filtered\ : std_logic;
signal \quad_counter0.A_delayed\ : std_logic;
signal \quad_counter1.n22\ : std_logic;
signal n2269 : std_logic;
signal n2268 : std_logic;
signal n2267 : std_logic;
signal n2266 : std_logic;
signal n2265 : std_logic;
signal n2264 : std_logic;
signal encoder0_position_15 : std_logic;
signal n2263 : std_logic;
signal n2262 : std_logic;
signal data_out_frame_6_4 : std_logic;
signal encoder0_position_25 : std_logic;
signal encoder0_position_10 : std_logic;
signal encoder0_position_20 : std_logic;
signal data_out_frame_7_4 : std_logic;
signal n2253 : std_logic;
signal n2249 : std_logic;
signal encoder0_position_30 : std_logic;
signal data_out_frame_6_1 : std_logic;
signal encoder0_position_1 : std_logic;
signal n2251 : std_logic;
signal encoder0_position_28 : std_logic;
signal encoder0_position_16 : std_logic;
signal encoder0_position_14 : std_logic;
signal data_out_frame_8_6 : std_logic;
signal encoder0_position_4 : std_logic;
signal \c0.n21632\ : std_logic;
signal \c0.n21299\ : std_logic;
signal data_out_frame_8_7 : std_logic;
signal \c0.n21626_cascade_\ : std_logic;
signal encoder0_position_7 : std_logic;
signal data_out_frame_9_7 : std_logic;
signal \c0.n11_adj_3472\ : std_logic;
signal \c0.n11_adj_3479\ : std_logic;
signal \c0.n11_adj_3444_cascade_\ : std_logic;
signal \c0.n21289_cascade_\ : std_logic;
signal \c0.n55_cascade_\ : std_logic;
signal \c0.n14301_cascade_\ : std_logic;
signal \c0.n15942\ : std_logic;
signal n6866 : std_logic;
signal data_out_frame_10_4 : std_logic;
signal \c0.n21288\ : std_logic;
signal n2273 : std_logic;
signal encoder0_position_6 : std_logic;
signal \c0.n21517\ : std_logic;
signal \c0.n21506_cascade_\ : std_logic;
signal \c0.n55\ : std_logic;
signal \c0.r_Bit_Index_2\ : std_logic;
signal \c0.n21414_cascade_\ : std_logic;
signal \c0.n11\ : std_logic;
signal \c0.n15938\ : std_logic;
signal \c0.tx.n8\ : std_logic;
signal \c0.tx.n4\ : std_logic;
signal \c0.tx.n21179_cascade_\ : std_logic;
signal \c0.r_Clock_Count_8\ : std_logic;
signal \c0.tx.n12759\ : std_logic;
signal \c0.FRAME_MATCHER_state_15\ : std_logic;
signal \c0.FRAME_MATCHER_state_10\ : std_logic;
signal \c0.FRAME_MATCHER_state_11\ : std_logic;
signal \c0.n18669\ : std_logic;
signal \c0.n18679\ : std_logic;
signal \c0.n18637\ : std_logic;
signal \c0.FRAME_MATCHER_state_22\ : std_logic;
signal \c0.n18635\ : std_logic;
signal \c0.FRAME_MATCHER_state_26\ : std_logic;
signal \c0.n18623\ : std_logic;
signal \c0.FRAME_MATCHER_state_13\ : std_logic;
signal \c0.n18665\ : std_logic;
signal \c0.FRAME_MATCHER_state_23\ : std_logic;
signal \c0.FRAME_MATCHER_state_20\ : std_logic;
signal \c0.n18651\ : std_logic;
signal \c0.n18625\ : std_logic;
signal \c0.n18641\ : std_logic;
signal b_delay_counter_0 : std_logic;
signal n187 : std_logic;
signal \bfn_12_5_0_\ : std_logic;
signal \quad_counter1.b_delay_counter_1\ : std_logic;
signal \quad_counter1.n17237\ : std_logic;
signal \quad_counter1.b_delay_counter_2\ : std_logic;
signal \quad_counter1.n17238\ : std_logic;
signal \quad_counter1.b_delay_counter_3\ : std_logic;
signal \quad_counter1.n17239\ : std_logic;
signal \quad_counter1.b_delay_counter_4\ : std_logic;
signal \quad_counter1.n17240\ : std_logic;
signal \quad_counter1.b_delay_counter_5\ : std_logic;
signal \quad_counter1.n17241\ : std_logic;
signal \quad_counter1.b_delay_counter_6\ : std_logic;
signal \quad_counter1.n17242\ : std_logic;
signal \quad_counter1.b_delay_counter_7\ : std_logic;
signal \quad_counter1.n17243\ : std_logic;
signal \quad_counter1.n17244\ : std_logic;
signal \quad_counter1.b_delay_counter_8\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \quad_counter1.b_delay_counter_9\ : std_logic;
signal \quad_counter1.n17245\ : std_logic;
signal \quad_counter1.b_delay_counter_10\ : std_logic;
signal \quad_counter1.n17246\ : std_logic;
signal \quad_counter1.b_delay_counter_11\ : std_logic;
signal \quad_counter1.n17247\ : std_logic;
signal \quad_counter1.b_delay_counter_12\ : std_logic;
signal \quad_counter1.n17248\ : std_logic;
signal \quad_counter1.b_delay_counter_13\ : std_logic;
signal \quad_counter1.n17249\ : std_logic;
signal \quad_counter1.b_delay_counter_14\ : std_logic;
signal \quad_counter1.n17250\ : std_logic;
signal \quad_counter1.n17251\ : std_logic;
signal \quad_counter1.b_delay_counter_15\ : std_logic;
signal n12417 : std_logic;
signal \b_delay_counter_15__N_2933\ : std_logic;
signal \PIN_12_c\ : std_logic;
signal \quadA_delayed_adj_3584\ : std_logic;
signal \a_delay_counter_15__N_2916_adj_3589_cascade_\ : std_logic;
signal \quad_counter1.n20\ : std_logic;
signal a_delay_counter_0_adj_3583 : std_logic;
signal n39_adj_3587 : std_logic;
signal \bfn_12_8_0_\ : std_logic;
signal \quad_counter1.a_delay_counter_1\ : std_logic;
signal \quad_counter1.n17252\ : std_logic;
signal \quad_counter1.a_delay_counter_2\ : std_logic;
signal \quad_counter1.n17253\ : std_logic;
signal \quad_counter1.a_delay_counter_3\ : std_logic;
signal \quad_counter1.n17254\ : std_logic;
signal \quad_counter1.a_delay_counter_4\ : std_logic;
signal \quad_counter1.n17255\ : std_logic;
signal \quad_counter1.a_delay_counter_5\ : std_logic;
signal \quad_counter1.n17256\ : std_logic;
signal \quad_counter1.a_delay_counter_6\ : std_logic;
signal \quad_counter1.n17257\ : std_logic;
signal \quad_counter1.a_delay_counter_7\ : std_logic;
signal \quad_counter1.n17258\ : std_logic;
signal \quad_counter1.n17259\ : std_logic;
signal \quad_counter1.a_delay_counter_8\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \quad_counter1.a_delay_counter_9\ : std_logic;
signal \quad_counter1.n17260\ : std_logic;
signal \quad_counter1.a_delay_counter_10\ : std_logic;
signal \quad_counter1.n17261\ : std_logic;
signal \quad_counter1.a_delay_counter_11\ : std_logic;
signal \quad_counter1.n17262\ : std_logic;
signal \quad_counter1.a_delay_counter_12\ : std_logic;
signal \quad_counter1.n17263\ : std_logic;
signal \quad_counter1.a_delay_counter_13\ : std_logic;
signal \quad_counter1.n17264\ : std_logic;
signal \quad_counter1.a_delay_counter_14\ : std_logic;
signal \quad_counter1.n17265\ : std_logic;
signal \quad_counter1.n17266\ : std_logic;
signal \quad_counter1.a_delay_counter_15\ : std_logic;
signal n12477 : std_logic;
signal \a_delay_counter_15__N_2916_adj_3589\ : std_logic;
signal data_out_frame_9_2 : std_logic;
signal data_out_frame_8_2 : std_logic;
signal \c0.n21650\ : std_logic;
signal \c0.n21564_cascade_\ : std_logic;
signal n2270 : std_logic;
signal n2250 : std_logic;
signal encoder0_position_13 : std_logic;
signal data_out_frame_11_6 : std_logic;
signal n2271 : std_logic;
signal data_out_frame_11_4 : std_logic;
signal \c0.n5_adj_3033\ : std_logic;
signal data_out_frame_12_6 : std_logic;
signal encoder0_position_17 : std_logic;
signal data_out_frame_7_1 : std_logic;
signal \c0.n6_adj_3324\ : std_logic;
signal data_out_frame_13_3 : std_logic;
signal data_out_frame_12_7 : std_logic;
signal data_out_frame_11_3 : std_logic;
signal data_out_frame_10_3 : std_logic;
signal encoder0_position_12 : std_logic;
signal data_out_frame_13_6 : std_logic;
signal \c0.n21301\ : std_logic;
signal \c0.n21653\ : std_logic;
signal \c0.n21305\ : std_logic;
signal \c0.n21570\ : std_logic;
signal \c0.n21307_cascade_\ : std_logic;
signal \c0.n21577\ : std_logic;
signal \n21578_cascade_\ : std_logic;
signal n21656 : std_logic;
signal data_out_frame_13_7 : std_logic;
signal \c0.n21467\ : std_logic;
signal \c0.tx.n21330\ : std_logic;
signal n9_adj_3588 : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal \c0.n9753_cascade_\ : std_logic;
signal data_out_frame_12_3 : std_logic;
signal \c0.n21456\ : std_logic;
signal \c0.r_Bit_Index_1\ : std_logic;
signal \c0.n21614\ : std_logic;
signal \c0.n32\ : std_logic;
signal \c0.n2_adj_3556_cascade_\ : std_logic;
signal \c0.n7_adj_3557\ : std_logic;
signal \c0.n21329\ : std_logic;
signal \c0.n19001_cascade_\ : std_logic;
signal \c0.n30_adj_3559\ : std_logic;
signal \c0.n12498\ : std_logic;
signal \c0.n15920\ : std_logic;
signal \r_SM_Main_1_adj_3592\ : std_logic;
signal n4_adj_3580 : std_logic;
signal n9_adj_3591 : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal \c0.n12512\ : std_logic;
signal \c0.r_SM_Main_0\ : std_logic;
signal \c0.n19023\ : std_logic;
signal \c0.n18609\ : std_logic;
signal \c0.FRAME_MATCHER_state_14\ : std_logic;
signal \c0.FRAME_MATCHER_state_9\ : std_logic;
signal \c0.n10_adj_3488\ : std_logic;
signal \c0.n15850_cascade_\ : std_logic;
signal \c0.n11427_cascade_\ : std_logic;
signal \c0.n16_adj_3484\ : std_logic;
signal \c0.FRAME_MATCHER_state_31\ : std_logic;
signal \c0.n19045_cascade_\ : std_logic;
signal \c0.n4_adj_3046\ : std_logic;
signal \c0.n19045\ : std_logic;
signal \c0.FRAME_MATCHER_state_25\ : std_logic;
signal \c0.FRAME_MATCHER_state_28\ : std_logic;
signal \c0.n10_adj_3438\ : std_logic;
signal \c0.n19050\ : std_logic;
signal \c0.FRAME_MATCHER_state_6\ : std_logic;
signal \c0.n63\ : std_logic;
signal \c0.rx.r_Rx_Data_R\ : std_logic;
signal \c0.FRAME_MATCHER_state_16\ : std_logic;
signal \c0.n18659\ : std_logic;
signal \c0.n19146\ : std_logic;
signal \c0.FRAME_MATCHER_state_3\ : std_logic;
signal \c0.n18633\ : std_logic;
signal \c0.FRAME_MATCHER_state_27\ : std_logic;
signal \c0.FRAME_MATCHER_state_19\ : std_logic;
signal \c0.FRAME_MATCHER_state_24\ : std_logic;
signal \c0.n17_adj_3486\ : std_logic;
signal \c0.FRAME_MATCHER_state_7\ : std_logic;
signal \c0.n18677\ : std_logic;
signal \c0.FRAME_MATCHER_state_30\ : std_logic;
signal \c0.n18601\ : std_logic;
signal \c0.n6_adj_3143_cascade_\ : std_logic;
signal \c0.n4_adj_3227\ : std_logic;
signal \quad_counter1.A_delayed\ : std_logic;
signal \B_filtered_adj_3582\ : std_logic;
signal \quad_counter1.B_delayed\ : std_logic;
signal \A_filtered_adj_3581\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \quad_counter1.count_direction\ : std_logic;
signal \quad_counter1.n17314\ : std_logic;
signal \quad_counter1.n17315\ : std_logic;
signal n2343 : std_logic;
signal \quad_counter1.n17316\ : std_logic;
signal \quad_counter1.n17317\ : std_logic;
signal n2341 : std_logic;
signal \quad_counter1.n17318\ : std_logic;
signal \quad_counter1.n17319\ : std_logic;
signal encoder1_position_6 : std_logic;
signal n2339 : std_logic;
signal \quad_counter1.n17320\ : std_logic;
signal \quad_counter1.n17321\ : std_logic;
signal encoder1_position_7 : std_logic;
signal n2338 : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal n2337 : std_logic;
signal \quad_counter1.n17322\ : std_logic;
signal n2336 : std_logic;
signal \quad_counter1.n17323\ : std_logic;
signal encoder1_position_10 : std_logic;
signal n2335 : std_logic;
signal \quad_counter1.n17324\ : std_logic;
signal encoder1_position_11 : std_logic;
signal n2334 : std_logic;
signal \quad_counter1.n17325\ : std_logic;
signal \quad_counter1.n17326\ : std_logic;
signal encoder1_position_13 : std_logic;
signal n2332 : std_logic;
signal \quad_counter1.n17327\ : std_logic;
signal encoder1_position_14 : std_logic;
signal n2331 : std_logic;
signal \quad_counter1.n17328\ : std_logic;
signal \quad_counter1.n17329\ : std_logic;
signal encoder1_position_15 : std_logic;
signal n2330 : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal encoder1_position_16 : std_logic;
signal n2329 : std_logic;
signal \quad_counter1.n17330\ : std_logic;
signal n2328 : std_logic;
signal \quad_counter1.n17331\ : std_logic;
signal n2327 : std_logic;
signal \quad_counter1.n17332\ : std_logic;
signal encoder1_position_19 : std_logic;
signal n2326 : std_logic;
signal \quad_counter1.n17333\ : std_logic;
signal encoder1_position_20 : std_logic;
signal n2325 : std_logic;
signal \quad_counter1.n17334\ : std_logic;
signal \quad_counter1.n17335\ : std_logic;
signal encoder1_position_22 : std_logic;
signal n2323 : std_logic;
signal \quad_counter1.n17336\ : std_logic;
signal \quad_counter1.n17337\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal n2321 : std_logic;
signal \quad_counter1.n17338\ : std_logic;
signal \quad_counter1.n17339\ : std_logic;
signal n2319 : std_logic;
signal \quad_counter1.n17340\ : std_logic;
signal encoder1_position_27 : std_logic;
signal n2318 : std_logic;
signal \quad_counter1.n17341\ : std_logic;
signal \quad_counter1.n17342\ : std_logic;
signal \quad_counter1.n17343\ : std_logic;
signal encoder1_position_30 : std_logic;
signal n2315 : std_logic;
signal \quad_counter1.n17344\ : std_logic;
signal \quad_counter1.n17345\ : std_logic;
signal \quad_counter1.n2301\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal n2314 : std_logic;
signal n2345 : std_logic;
signal data_out_frame_12_5 : std_logic;
signal encoder1_position_4 : std_logic;
signal data_out_frame_13_4 : std_logic;
signal encoder1_position_31 : std_logic;
signal n2320 : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal data_out_frame_9_4 : std_logic;
signal data_out_frame_8_4 : std_logic;
signal \c0.n21287\ : std_logic;
signal encoder0_position_9 : std_logic;
signal encoder1_position_24 : std_logic;
signal \c0.data_out_frame_0_4\ : std_logic;
signal encoder0_position_8 : std_logic;
signal encoder0_position_0 : std_logic;
signal encoder1_position_25 : std_logic;
signal encoder1_position_2 : std_logic;
signal encoder1_position_17 : std_logic;
signal data_out_frame_13_2 : std_logic;
signal data_out_frame_12_2 : std_logic;
signal \c0.n11_adj_3108\ : std_logic;
signal data_out_frame_10_1 : std_logic;
signal data_out_frame_11_1 : std_logic;
signal data_out_frame_13_5 : std_logic;
signal \c0.r_SM_Main_2_N_2547_0\ : std_logic;
signal tx_active : std_logic;
signal \c0.n15842\ : std_logic;
signal \c0.n11_adj_3404\ : std_logic;
signal \c0.n7_adj_3333\ : std_logic;
signal data_out_frame_9_1 : std_logic;
signal \c0.n21605\ : std_logic;
signal data_out_frame_8_1 : std_logic;
signal \c0.n21608_cascade_\ : std_logic;
signal \c0.r_Tx_Data_0\ : std_logic;
signal \c0.n21466\ : std_logic;
signal encoder1_position_9 : std_logic;
signal \c0.n21566\ : std_logic;
signal \n10_cascade_\ : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal data_out_frame_12_1 : std_logic;
signal \c0.n11_adj_3104\ : std_logic;
signal n10_adj_3593 : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \c0.n17346\ : std_logic;
signal \c0.n17347\ : std_logic;
signal \c0.n17348\ : std_logic;
signal \c0.n17349\ : std_logic;
signal \c0.n17350\ : std_logic;
signal \c0.n17351\ : std_logic;
signal \c0.n17352\ : std_logic;
signal \c0.n19052\ : std_logic;
signal \c0.n6_adj_3338\ : std_logic;
signal \c0.n12326\ : std_logic;
signal \c0.n12326_cascade_\ : std_logic;
signal \c0.n12758\ : std_logic;
signal \c0.n4_adj_3263_cascade_\ : std_logic;
signal \c0.n936_cascade_\ : std_logic;
signal \c0.tx_transmit_N_2443\ : std_logic;
signal \c0.n21420\ : std_logic;
signal \c0.FRAME_MATCHER_state_21\ : std_logic;
signal \c0.n18627\ : std_logic;
signal \c0.n19650\ : std_logic;
signal \c0.n19638_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_31_N_1864_2\ : std_logic;
signal \c0.n6_adj_3521_cascade_\ : std_logic;
signal \c0.n936\ : std_logic;
signal \c0.n11_adj_3370\ : std_logic;
signal \c0.n19638\ : std_logic;
signal \c0.n6_adj_3515_cascade_\ : std_logic;
signal \c0.n5_adj_3516\ : std_logic;
signal \c0.FRAME_MATCHER_state_5\ : std_logic;
signal \c0.n18681\ : std_logic;
signal \c0.FRAME_MATCHER_state_17\ : std_logic;
signal \c0.n18657\ : std_logic;
signal \c0.FRAME_MATCHER_state_4\ : std_logic;
signal \c0.n18629\ : std_logic;
signal \bfn_14_5_0_\ : std_logic;
signal \c0.n17176\ : std_logic;
signal \c0.n2_adj_3144\ : std_logic;
signal \c0.n17177\ : std_logic;
signal \c0.n2_adj_3145\ : std_logic;
signal \c0.n17178\ : std_logic;
signal \c0.n17179\ : std_logic;
signal \c0.n17180\ : std_logic;
signal \c0.n17180_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17180_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17180_THRU_CRY_2_THRU_CO\ : std_logic;
signal \bfn_14_6_0_\ : std_logic;
signal \c0.n17181\ : std_logic;
signal \c0.n17181_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17181_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17181_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17181_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17181_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17181_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17181_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \c0.n17182\ : std_logic;
signal \c0.n17182_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17182_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17182_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17182_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17182_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17182_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17182_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \c0.n17183\ : std_logic;
signal \c0.n17183_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17183_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17183_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17183_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17183_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17183_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17183_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \c0.n17184\ : std_logic;
signal \c0.n17184_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17184_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17184_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17184_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17184_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17184_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17184_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \c0.n17185\ : std_logic;
signal \c0.n17185_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17185_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17185_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17185_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17185_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17185_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17185_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \c0.n17186\ : std_logic;
signal \c0.n17186_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17186_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17186_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17186_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17186_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17186_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17186_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \c0.n17187\ : std_logic;
signal \c0.n17187_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17187_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17187_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17187_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17187_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17187_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17187_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \c0.n17188\ : std_logic;
signal \c0.n17188_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17188_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17188_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17188_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17188_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17188_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17188_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \c0.n6_adj_3162\ : std_logic;
signal \c0.n17189\ : std_logic;
signal \c0.n17189_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17189_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17189_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17189_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17189_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17189_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17189_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \c0.n17190\ : std_logic;
signal \c0.n17190_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17190_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17190_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17190_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17190_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17190_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17190_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \c0.n17191\ : std_logic;
signal \c0.n17191_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17191_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17191_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17191_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17191_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17191_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17191_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \c0.n17192\ : std_logic;
signal \c0.n17192_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17192_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17192_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17192_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17192_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17192_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17192_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \c0.n6_adj_3188\ : std_logic;
signal \c0.n17193\ : std_logic;
signal \c0.n17193_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17193_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17193_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17193_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17193_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17193_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17193_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \c0.n6_adj_3186\ : std_logic;
signal \c0.n17194\ : std_logic;
signal \c0.n17194_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17194_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17194_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17194_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17194_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17194_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17194_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \c0.n6_adj_3184\ : std_logic;
signal \c0.n17195\ : std_logic;
signal \c0.n17195_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17195_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17195_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17195_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17195_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17195_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17195_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \c0.n6_adj_3182\ : std_logic;
signal \c0.n17196\ : std_logic;
signal \c0.n17196_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17196_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17196_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17196_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17196_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17196_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17196_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal \c0.n6_adj_3180\ : std_logic;
signal \c0.n17197\ : std_logic;
signal \c0.n17197_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17197_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17197_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17197_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17197_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17197_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17197_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_23_0_\ : std_logic;
signal \c0.n6_adj_3178\ : std_logic;
signal \c0.n17198\ : std_logic;
signal \c0.n17198_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17198_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17198_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17198_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17198_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17198_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17198_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal \c0.n17199\ : std_logic;
signal \c0.n17199_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17199_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17199_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17199_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17199_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17199_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17199_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_25_0_\ : std_logic;
signal \c0.n17200\ : std_logic;
signal \c0.n17200_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17200_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17200_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17200_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17200_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17200_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17200_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_26_0_\ : std_logic;
signal \c0.n17201\ : std_logic;
signal \c0.n17201_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17201_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17201_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17201_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17201_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17201_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17201_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_27_0_\ : std_logic;
signal \c0.n17202\ : std_logic;
signal \c0.n17202_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17202_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17202_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17202_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17202_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17202_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17202_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_28_0_\ : std_logic;
signal \c0.n17203\ : std_logic;
signal \c0.n17203_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17203_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17203_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17203_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17203_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17203_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17203_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_29_0_\ : std_logic;
signal \c0.n17204\ : std_logic;
signal \c0.n17204_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17204_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17204_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17204_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17204_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17204_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17204_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_30_0_\ : std_logic;
signal \c0.n17205\ : std_logic;
signal \c0.n17205_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17205_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17205_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17205_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17205_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n17205_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17205_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_31_0_\ : std_logic;
signal \c0.n17206\ : std_logic;
signal \c0.n17206_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n17206_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n17206_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n17206_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n17206_THRU_CRY_4_THRU_CO\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \c0.n17206_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n17206_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_14_32_0_\ : std_logic;
signal n20764 : std_logic;
signal n16 : std_logic;
signal \c0.n6_adj_3155\ : std_logic;
signal encoder0_position_24 : std_logic;
signal n2340 : std_logic;
signal encoder1_position_5 : std_logic;
signal \c0.n21647\ : std_logic;
signal encoder1_position_26 : std_logic;
signal data_out_frame_10_2 : std_logic;
signal \c0.n6_adj_3154\ : std_logic;
signal data_out_frame_6_0 : std_logic;
signal \c0.n6_adj_3321\ : std_logic;
signal n2344 : std_logic;
signal data_out_frame_28_4 : std_logic;
signal n2342 : std_logic;
signal encoder1_position_3 : std_logic;
signal encoder0_position_19 : std_logic;
signal \c0.n6_adj_3379_cascade_\ : std_logic;
signal n2324 : std_logic;
signal encoder1_position_21 : std_logic;
signal \c0.n21559\ : std_logic;
signal \c0.n5_adj_3102\ : std_logic;
signal n2322 : std_logic;
signal encoder0_position_11 : std_logic;
signal data_out_frame_10_7 : std_logic;
signal \c0.n21623\ : std_logic;
signal data_out_frame_9_3 : std_logic;
signal \c0.n21641\ : std_logic;
signal data_out_frame_8_3 : std_logic;
signal \c0.n21644\ : std_logic;
signal data_out_frame_11_5 : std_logic;
signal data_out_frame_8_5 : std_logic;
signal \c0.n21635_cascade_\ : std_logic;
signal data_out_frame_9_5 : std_logic;
signal data_out_frame_5_3 : std_logic;
signal \c0.n21470\ : std_logic;
signal \c0.n21542\ : std_logic;
signal n2316 : std_logic;
signal \c0.n6_adj_3156\ : std_logic;
signal encoder1_position_29 : std_logic;
signal data_out_frame_10_5 : std_logic;
signal encoder0_position_29 : std_logic;
signal \c0.data_out_frame_7_0\ : std_logic;
signal \c0.n17150\ : std_logic;
signal encoder1_position_18 : std_logic;
signal data_out_frame_11_2 : std_logic;
signal data_out_frame_10_0 : std_logic;
signal data_out_frame_11_0 : std_logic;
signal data_out_frame_8_0 : std_logic;
signal \c0.n21617_cascade_\ : std_logic;
signal data_out_frame_9_0 : std_logic;
signal \c0.n21620_cascade_\ : std_logic;
signal \c0.n21574\ : std_logic;
signal \c0.byte_transmit_counter_6\ : std_logic;
signal \c0.byte_transmit_counter_7\ : std_logic;
signal \c0.n7235\ : std_logic;
signal \c0.n2_adj_3147\ : std_logic;
signal \c0.n6_adj_3151\ : std_logic;
signal encoder0_position_21 : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal data_out_frame_7_5 : std_logic;
signal data_out_frame_6_5 : std_logic;
signal \c0.n5_adj_3447\ : std_logic;
signal byte_transmit_counter_5 : std_logic;
signal n9377 : std_logic;
signal data_out_frame_5_5 : std_logic;
signal \c0.n21546\ : std_logic;
signal \c0.n6_adj_3192\ : std_logic;
signal encoder1_position_1 : std_logic;
signal data_out_frame_13_1 : std_logic;
signal \c0.n6_adj_3190\ : std_logic;
signal \c0.rx.n14601_cascade_\ : std_logic;
signal n12301 : std_logic;
signal \c0.n15685\ : std_logic;
signal \c0.rx.n6\ : std_logic;
signal \n12492_cascade_\ : std_logic;
signal \c0.r_Bit_Index_0\ : std_logic;
signal tx_o : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal \c0.r_SM_Main_2\ : std_logic;
signal \c0.n21611\ : std_logic;
signal encoder0_position_23 : std_logic;
signal data_out_frame_7_7 : std_logic;
signal n13179 : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal \c0.rx.n17267\ : std_logic;
signal n12908 : std_logic;
signal \c0.rx.n17268\ : std_logic;
signal \c0.rx.n17269\ : std_logic;
signal \c0.rx.n17270\ : std_logic;
signal \c0.rx.n17271\ : std_logic;
signal \c0.rx.n17272\ : std_logic;
signal \c0.rx.n3\ : std_logic;
signal \c0.rx.n17273\ : std_logic;
signal \c0.rx.n7\ : std_logic;
signal \c0.FRAME_MATCHER_i_8\ : std_logic;
signal \c0.FRAME_MATCHER_i_19\ : std_logic;
signal \c0.n6_adj_3161\ : std_logic;
signal \c0.FRAME_MATCHER_i_25\ : std_logic;
signal \c0.n6_adj_3172\ : std_logic;
signal \c0.n6_adj_3194\ : std_logic;
signal \c0.FRAME_MATCHER_i_12\ : std_logic;
signal \c0.FRAME_MATCHER_i_20\ : std_logic;
signal \c0.FRAME_MATCHER_i_14\ : std_logic;
signal \c0.FRAME_MATCHER_i_7\ : std_logic;
signal \c0.n6_adj_3160\ : std_logic;
signal \c0.FRAME_MATCHER_i_22\ : std_logic;
signal \c0.FRAME_MATCHER_i_16\ : std_logic;
signal \c0.FRAME_MATCHER_i_11\ : std_logic;
signal \c0.n41_adj_3258_cascade_\ : std_logic;
signal \c0.n43_adj_3257\ : std_logic;
signal \c0.FRAME_MATCHER_i_10\ : std_logic;
signal \c0.FRAME_MATCHER_i_15\ : std_logic;
signal \c0.FRAME_MATCHER_i_13\ : std_logic;
signal \c0.FRAME_MATCHER_i_9\ : std_logic;
signal \c0.n40_adj_3259\ : std_logic;
signal \c0.n45_adj_3262\ : std_logic;
signal \c0.n39_adj_3260_cascade_\ : std_logic;
signal \c0.n50_adj_3261\ : std_logic;
signal \c0.n11432\ : std_logic;
signal \c0.n14_adj_3080_cascade_\ : std_logic;
signal \c0.n10_adj_3081\ : std_logic;
signal \c0.n4812\ : std_logic;
signal \c0.n19119\ : std_logic;
signal \c0.n19119_cascade_\ : std_logic;
signal \c0.n21273\ : std_logic;
signal \c0.n5_adj_3306_cascade_\ : std_logic;
signal \c0.n2_adj_3302\ : std_logic;
signal \c0.n11433_cascade_\ : std_logic;
signal \c0.n8_adj_3228_cascade_\ : std_logic;
signal \c0.n2103\ : std_logic;
signal \c0.n2103_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_29\ : std_logic;
signal \c0.n18653\ : std_logic;
signal \c0.FRAME_MATCHER_state_31_N_1736_2\ : std_logic;
signal \c0.FRAME_MATCHER_state_31_N_1736_1\ : std_logic;
signal \c0.n6_adj_3176\ : std_logic;
signal \c0.n11433\ : std_logic;
signal \c0.n700\ : std_logic;
signal \c0.n1\ : std_logic;
signal \c0.FRAME_MATCHER_i_21\ : std_logic;
signal \c0.FRAME_MATCHER_i_17\ : std_logic;
signal \c0.n44_adj_3255\ : std_logic;
signal \c0.FRAME_MATCHER_i_24\ : std_logic;
signal \c0.n6_adj_3174\ : std_logic;
signal \c0.FRAME_MATCHER_state_8\ : std_logic;
signal \c0.n18675\ : std_logic;
signal n11289 : std_logic;
signal \c0.FRAME_MATCHER_i_26\ : std_logic;
signal \n2108_cascade_\ : std_logic;
signal \c0.n6_adj_3170\ : std_logic;
signal \c0.n6_adj_3165\ : std_logic;
signal \c0.FRAME_MATCHER_i_27\ : std_logic;
signal \c0.n6_adj_3168\ : std_logic;
signal \c0.FRAME_MATCHER_i_28\ : std_logic;
signal \c0.n6_adj_3166\ : std_logic;
signal \c0.n6_adj_3159\ : std_logic;
signal \c0.FRAME_MATCHER_i_30\ : std_logic;
signal \c0.n6_adj_3164\ : std_logic;
signal \c0.n6_adj_3150\ : std_logic;
signal n2333 : std_logic;
signal \c0.n21319\ : std_logic;
signal encoder0_position_18 : std_logic;
signal \c0.n21317\ : std_logic;
signal count_enable : std_logic;
signal n2252 : std_logic;
signal encoder0_position_27 : std_logic;
signal data_out_frame_7_3 : std_logic;
signal data_out_frame_6_3 : std_logic;
signal \c0.n5_adj_3380\ : std_logic;
signal \c0.n21320\ : std_logic;
signal \c0.n21562\ : std_logic;
signal \c0.n21322_cascade_\ : std_logic;
signal n10_adj_3594 : std_logic;
signal data_out_frame_7_2 : std_logic;
signal \c0.n5_adj_3106\ : std_logic;
signal encoder0_position_26 : std_logic;
signal data_out_frame_6_2 : std_logic;
signal \c0.data_out_frame_0_2\ : std_logic;
signal \c0.n21473_cascade_\ : std_logic;
signal \c0.n6_adj_3105\ : std_logic;
signal data_out_frame_28_6 : std_logic;
signal \c0.data_out_frame_0_3\ : std_logic;
signal \c0.n11_adj_3325\ : std_logic;
signal encoder1_position_8 : std_logic;
signal data_out_frame_12_0 : std_logic;
signal encoder1_position_23 : std_logic;
signal data_out_frame_11_7 : std_logic;
signal n2317 : std_logic;
signal count_enable_adj_3586 : std_logic;
signal encoder1_position_28 : std_logic;
signal data_out_frame_5_6 : std_logic;
signal data_out_frame_29_3 : std_logic;
signal \c0.data_out_frame_28_3\ : std_logic;
signal \c0.n9753\ : std_logic;
signal \c0.n26_adj_3382_cascade_\ : std_logic;
signal \c0.n21314\ : std_logic;
signal \c0.n21316\ : std_logic;
signal data_out_frame_5_4 : std_logic;
signal \c0.n21465\ : std_logic;
signal \c0.data_out_frame_5_0\ : std_logic;
signal control_mode_5 : std_logic;
signal \c0.n21638\ : std_logic;
signal \c0.n11_adj_3462\ : std_logic;
signal data_out_frame_5_2 : std_logic;
signal \c0.rx.n9\ : std_logic;
signal n12920 : std_logic;
signal \c0.n70\ : std_logic;
signal \c0.n15850\ : std_logic;
signal \c0.n21231\ : std_logic;
signal \c0.n12254\ : std_logic;
signal encoder1_position_12 : std_logic;
signal data_out_frame_12_4 : std_logic;
signal data_out_frame_5_7 : std_logic;
signal \c0.n5_adj_3475\ : std_logic;
signal \c0.byte_transmit_counter_2\ : std_logic;
signal \c0.n21576_cascade_\ : std_logic;
signal \c0.byte_transmit_counter_1\ : std_logic;
signal \c0.n21302_cascade_\ : std_logic;
signal \c0.n21304_cascade_\ : std_logic;
signal \c0.n21572\ : std_logic;
signal n9 : std_logic;
signal \c0.n9755\ : std_logic;
signal data_out_frame_28_5 : std_logic;
signal \c0.n21308\ : std_logic;
signal byte_transmit_counter_4 : std_logic;
signal byte_transmit_counter_3 : std_logic;
signal \c0.n21310_cascade_\ : std_logic;
signal \c0.n21568\ : std_logic;
signal n9_adj_3590 : std_logic;
signal \c0.rx.n11302\ : std_logic;
signal \c0.rx.n11302_cascade_\ : std_logic;
signal encoder1_position_0 : std_logic;
signal data_out_frame_13_0 : std_logic;
signal \c0.rx.n21451_cascade_\ : std_logic;
signal \c0.rx.n15906_cascade_\ : std_logic;
signal \c0.rx.n20851\ : std_logic;
signal \c0.rx.n32\ : std_logic;
signal \c0.rx.n20964\ : std_logic;
signal \c0.rx.n15906\ : std_logic;
signal \r_SM_Main_2_N_2473_2_cascade_\ : std_logic;
signal \c0.rx.n15926\ : std_logic;
signal \c0.rx.n35_cascade_\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal \c0.rx.n12_cascade_\ : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal \c0.rx.n21406_cascade_\ : std_logic;
signal \r_SM_Main_2_N_2473_2\ : std_logic;
signal \c0.rx.r_Clock_Count_6\ : std_logic;
signal \c0.rx.r_Clock_Count_2\ : std_logic;
signal \c0.rx.r_Clock_Count_0\ : std_logic;
signal \c0.rx.r_Clock_Count_1\ : std_logic;
signal \c0.rx.n8\ : std_logic;
signal n12914 : std_logic;
signal n12917 : std_logic;
signal \c0.n11440\ : std_logic;
signal \c0.n11317_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31\ : std_logic;
signal \c0.rx.r_Clock_Count_4\ : std_logic;
signal \c0.rx.r_Clock_Count_5\ : std_logic;
signal \c0.rx.n21267\ : std_logic;
signal \c0.FRAME_MATCHER_i_18\ : std_logic;
signal \c0.FRAME_MATCHER_i_23\ : std_logic;
signal \c0.FRAME_MATCHER_i_29\ : std_logic;
signal \c0.n42_adj_3256\ : std_logic;
signal \c0.n1_adj_3002\ : std_logic;
signal \c0.n21053\ : std_logic;
signal \c0.n11_adj_3093\ : std_logic;
signal \c0.n15701_cascade_\ : std_logic;
signal \n11421_cascade_\ : std_logic;
signal \c0.n11422\ : std_logic;
signal \c0.n3632\ : std_logic;
signal \c0.n9389\ : std_logic;
signal \c0.n3\ : std_logic;
signal \c0.n11427\ : std_logic;
signal \c0.n15874\ : std_logic;
signal \c0.n121\ : std_logic;
signal \c0.n103\ : std_logic;
signal \c0.n63_adj_3084\ : std_logic;
signal \c0.n19_adj_3252\ : std_logic;
signal \c0.n21_adj_3253\ : std_logic;
signal \c0.n19_adj_3252_cascade_\ : std_logic;
signal \c0.n63_adj_3083\ : std_logic;
signal \c0.n7804\ : std_logic;
signal \c0.n21281_cascade_\ : std_logic;
signal \c0.n108\ : std_logic;
signal \c0.n108_cascade_\ : std_logic;
signal \c0.n92_adj_3254\ : std_logic;
signal data_in_1_2 : std_logic;
signal \c0.n26_adj_3107\ : std_logic;
signal \c0.n38_adj_3328\ : std_logic;
signal \c0.n21279_cascade_\ : std_logic;
signal \c0.n21255_cascade_\ : std_logic;
signal \c0.n37_adj_3332\ : std_logic;
signal \c0.n63_adj_3417_cascade_\ : std_logic;
signal \c0.n5_adj_3040_cascade_\ : std_logic;
signal \c0.n30_adj_3264\ : std_logic;
signal \c0.data_in_frame_5_0\ : std_logic;
signal \c0.data_in_frame_9_7\ : std_logic;
signal \c0.n19115_cascade_\ : std_logic;
signal \c0.data_in_frame_10_1\ : std_logic;
signal \c0.n63_adj_3146\ : std_logic;
signal \c0.n20_adj_3437_cascade_\ : std_logic;
signal \n21222_cascade_\ : std_logic;
signal control_mode_6 : std_logic;
signal control_mode_2 : std_logic;
signal control_mode_4 : std_logic;
signal control_mode_3 : std_logic;
signal control_mode_7 : std_logic;
signal \c0.n9_cascade_\ : std_logic;
signal \c0.n16_adj_3008_cascade_\ : std_logic;
signal \c0.n9\ : std_logic;
signal \c0.n19449_cascade_\ : std_logic;
signal control_mode_0 : std_logic;
signal \FRAME_MATCHER_state_31_N_1800_2\ : std_logic;
signal \FRAME_MATCHER_state_2\ : std_logic;
signal \c0.n15499\ : std_logic;
signal \c0.n13_adj_3016\ : std_logic;
signal \c0.FRAME_MATCHER_rx_data_ready_prev\ : std_logic;
signal \c0.n19111_cascade_\ : std_logic;
signal \c0.n19493\ : std_logic;
signal \c0.n16\ : std_logic;
signal \c0.n24\ : std_logic;
signal \c0.n28_cascade_\ : std_logic;
signal \c0.n12026_cascade_\ : std_logic;
signal \c0.n10_cascade_\ : std_logic;
signal \c0.n21104\ : std_logic;
signal \n3846_cascade_\ : std_logic;
signal \c0.rx.r_Clock_Count_7\ : std_logic;
signal \c0.rx.n6_adj_2995\ : std_logic;
signal \c0.rx.n11455\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_2479_0\ : std_logic;
signal n3792 : std_logic;
signal n12911 : std_logic;
signal \c0.rx.r_Clock_Count_3\ : std_logic;
signal \c0.rx.n15860\ : std_logic;
signal \c0.n19449\ : std_logic;
signal n12492 : std_logic;
signal n12835 : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal \c0.n22_adj_3276_cascade_\ : std_logic;
signal \c0.n36_adj_3277_cascade_\ : std_logic;
signal \c0.n20415_cascade_\ : std_logic;
signal \c0.n14_adj_3407_cascade_\ : std_logic;
signal \c0.n100_adj_3403\ : std_logic;
signal \c0.n18_adj_3412\ : std_logic;
signal \c0.n20300_cascade_\ : std_logic;
signal \c0.n20300\ : std_logic;
signal \c0.FRAME_MATCHER_state_0\ : std_logic;
signal \c0.n3235\ : std_logic;
signal \c0.data_in_frame_28_6\ : std_logic;
signal \c0.n17947_cascade_\ : std_logic;
signal \c0.n20793\ : std_logic;
signal \c0.n10_adj_3242_cascade_\ : std_logic;
signal data_in_0_2 : std_logic;
signal \c0.n14_adj_3243\ : std_logic;
signal \c0.n105\ : std_logic;
signal data_in_3_3 : std_logic;
signal data_in_3_1 : std_logic;
signal data_in_0_7 : std_logic;
signal data_in_1_6 : std_logic;
signal \c0.n18_adj_3229\ : std_logic;
signal \c0.n11446\ : std_logic;
signal \c0.n21108_cascade_\ : std_logic;
signal \c0.n12_adj_3248\ : std_logic;
signal data_in_3_5 : std_logic;
signal \c0.n20_adj_3250\ : std_logic;
signal data_in_2_3 : std_logic;
signal data_in_1_3 : std_logic;
signal data_in_0_6 : std_logic;
signal data_in_0_3 : std_logic;
signal \c0.n18_adj_3246\ : std_logic;
signal \c0.n20_cascade_\ : std_logic;
signal \c0.n16_adj_3247\ : std_logic;
signal \c0.n11311\ : std_logic;
signal data_in_3_2 : std_logic;
signal data_in_0_5 : std_logic;
signal \c0.n5_adj_2999\ : std_logic;
signal \c0.FRAME_MATCHER_state_18\ : std_logic;
signal \c0.n18655\ : std_logic;
signal \c0.FRAME_MATCHER_i_4\ : std_logic;
signal \c0.FRAME_MATCHER_i_6\ : std_logic;
signal \c0.FRAME_MATCHER_i_3\ : std_logic;
signal \c0.n20224_cascade_\ : std_logic;
signal \c0.n19_cascade_\ : std_logic;
signal \c0.n20246_cascade_\ : std_logic;
signal \c0.n24_adj_3327\ : std_logic;
signal \c0.n23_adj_3039_cascade_\ : std_logic;
signal \c0.n23_adj_3039\ : std_logic;
signal \c0.n30_adj_3042\ : std_logic;
signal data_out_frame_29_2 : std_logic;
signal \c0.n18428_cascade_\ : std_logic;
signal \c0.n29_adj_3446\ : std_logic;
signal data_out_frame_28_2 : std_logic;
signal \c0.data_out_frame_28__0__N_708_cascade_\ : std_logic;
signal \c0.data_out_frame_28__0__N_708\ : std_logic;
signal \c0.data_out_frame_29_0\ : std_logic;
signal \c0.data_out_frame_29_1\ : std_logic;
signal data_out_frame_28_1 : std_logic;
signal \c0.byte_transmit_counter_0\ : std_logic;
signal \c0.n26_adj_3103\ : std_logic;
signal \c0.n20209\ : std_logic;
signal \c0.n20204\ : std_logic;
signal \c0.n19217_cascade_\ : std_logic;
signal \c0.n66\ : std_logic;
signal n21222 : std_logic;
signal control_mode_1 : std_logic;
signal \c0.n16_adj_3018\ : std_logic;
signal \c0.n32_adj_3493_cascade_\ : std_logic;
signal \c0.n36_adj_3547_cascade_\ : std_logic;
signal \c0.n63_adj_3417\ : std_logic;
signal \c0.n38_adj_3548_cascade_\ : std_logic;
signal \c0.n34_adj_3411\ : std_logic;
signal \c0.n18443_cascade_\ : std_logic;
signal \c0.n25_adj_3495\ : std_logic;
signal \c0.data_in_frame_9_4\ : std_logic;
signal \c0.n25_adj_3495_cascade_\ : std_logic;
signal \c0.n6_adj_3005\ : std_logic;
signal \c0.n13\ : std_logic;
signal \c0.n20_adj_3539\ : std_logic;
signal \c0.n12_adj_3001_cascade_\ : std_logic;
signal \c0.n20403_cascade_\ : std_logic;
signal \c0.n10_adj_3514\ : std_logic;
signal \c0.n20398_cascade_\ : std_logic;
signal \c0.n4_adj_3071\ : std_logic;
signal \c0.n5_adj_3003\ : std_logic;
signal \c0.n36_adj_3267_cascade_\ : std_logic;
signal \c0.n94\ : std_logic;
signal \c0.n12_adj_3004\ : std_logic;
signal data_in_frame_18_6 : std_logic;
signal n4_adj_3595 : std_logic;
signal \c0.n14_adj_3434\ : std_logic;
signal \c0.FRAME_MATCHER_state_12\ : std_logic;
signal \c0.n14\ : std_logic;
signal \c0.n18667\ : std_logic;
signal \c0.n61_cascade_\ : std_logic;
signal \c0.n50\ : std_logic;
signal \c0.n61\ : std_logic;
signal \c0.n86_adj_3393_cascade_\ : std_logic;
signal \c0.n95_cascade_\ : std_logic;
signal \c0.n15_adj_3441\ : std_logic;
signal data_in_3_7 : std_logic;
signal data_in_frame_16_6 : std_logic;
signal \c0.data_in_frame_28_4\ : std_logic;
signal \c0.n20931\ : std_logic;
signal \c0.n18537\ : std_logic;
signal \c0.n20370\ : std_logic;
signal \c0.data_in_frame_29_7\ : std_logic;
signal \c0.data_in_frame_29_6\ : std_logic;
signal \c0.n10_adj_3152_cascade_\ : std_logic;
signal \c0.n21117\ : std_logic;
signal \c0.data_in_frame_29_0\ : std_logic;
signal \c0.n21117_cascade_\ : std_logic;
signal \c0.n18\ : std_logic;
signal \c0.n5_adj_3142\ : std_logic;
signal \c0.n5_adj_3142_cascade_\ : std_logic;
signal \c0.n22_adj_3305_cascade_\ : std_logic;
signal \c0.n37_adj_3309_cascade_\ : std_logic;
signal \c0.n21099_cascade_\ : std_logic;
signal \c0.n18_adj_3314\ : std_logic;
signal \c0.n10_adj_3353_cascade_\ : std_logic;
signal \c0.n21111\ : std_logic;
signal \c0.n9_adj_3352_cascade_\ : std_logic;
signal \c0.n21051\ : std_logic;
signal \c0.data_in_frame_27_7\ : std_logic;
signal \c0.data_in_frame_27_6\ : std_logic;
signal \c0.data_in_frame_26_4\ : std_logic;
signal data_in_2_2 : std_logic;
signal \c0.n10_adj_3238\ : std_logic;
signal \c0.n110\ : std_logic;
signal data_in_2_5 : std_logic;
signal data_in_1_5 : std_logic;
signal \c0.n160\ : std_logic;
signal data_in_2_0 : std_logic;
signal data_in_1_0 : std_logic;
signal \c0.n12_adj_3230\ : std_logic;
signal data_in_2_7 : std_logic;
signal \c0.n11443\ : std_logic;
signal data_in_0_1 : std_logic;
signal \FRAME_MATCHER_state_1\ : std_logic;
signal n4_adj_3596 : std_logic;
signal n11421 : std_logic;
signal n1295 : std_logic;
signal \c0.n26\ : std_logic;
signal \c0.n5_adj_3044\ : std_logic;
signal \c0.n25_adj_3045\ : std_logic;
signal \c0.n14_adj_3073_cascade_\ : std_logic;
signal \c0.n10_adj_3068\ : std_logic;
signal \c0.n22_adj_3041\ : std_logic;
signal \c0.n21079\ : std_logic;
signal \c0.n11516\ : std_logic;
signal \c0.n14_adj_3480\ : std_logic;
signal \c0.n13_adj_3490_cascade_\ : std_logic;
signal \c0.n13_adj_3546\ : std_logic;
signal \c0.n15497\ : std_logic;
signal \c0.n14_adj_3459\ : std_logic;
signal \c0.n6_adj_3453\ : std_logic;
signal \c0.n39_adj_3398_cascade_\ : std_logic;
signal \c0.n13_adj_3526\ : std_logic;
signal \c0.n14_adj_3525\ : std_logic;
signal \c0.n15_adj_3543\ : std_logic;
signal \c0.n13_adj_3526_cascade_\ : std_logic;
signal \c0.n11_adj_3394\ : std_logic;
signal \c0.n28_adj_3519\ : std_logic;
signal \c0.n16_adj_3416_cascade_\ : std_logic;
signal \c0.n16_adj_3542\ : std_logic;
signal \c0.n5_adj_3528\ : std_logic;
signal \c0.n78_cascade_\ : std_logic;
signal \c0.n30_adj_3119_cascade_\ : std_logic;
signal \c0.n20088\ : std_logic;
signal \c0.n20055_cascade_\ : std_logic;
signal \c0.n5_adj_3099\ : std_logic;
signal \c0.n37_adj_3110_cascade_\ : std_logic;
signal \c0.n22_adj_3115\ : std_logic;
signal \c0.n6_adj_3024_cascade_\ : std_logic;
signal \c0.n18435_cascade_\ : std_logic;
signal \c0.data_in_frame_10_2\ : std_logic;
signal \c0.n14_adj_3007\ : std_logic;
signal \c0.n31_adj_3121\ : std_logic;
signal \c0.n27\ : std_logic;
signal \c0.n28_adj_3120_cascade_\ : std_logic;
signal \c0.n33_adj_3122\ : std_logic;
signal \c0.n20052_cascade_\ : std_logic;
signal \c0.n10_adj_3129_cascade_\ : std_logic;
signal \c0.n18400_cascade_\ : std_logic;
signal \c0.n5_adj_3040\ : std_logic;
signal \c0.n42_adj_3560\ : std_logic;
signal \c0.n35_adj_3342_cascade_\ : std_logic;
signal \c0.n39_adj_3339\ : std_logic;
signal \c0.n12_adj_3015\ : std_logic;
signal \c0.n44_adj_3561_cascade_\ : std_logic;
signal \c0.n13_adj_3017\ : std_logic;
signal \c0.n21118\ : std_logic;
signal data_in_frame_18_2 : std_logic;
signal \c0.n21118_cascade_\ : std_logic;
signal \c0.n13_adj_3139\ : std_logic;
signal \c0.n36_adj_3267\ : std_logic;
signal \c0.n96_adj_3418_cascade_\ : std_logic;
signal \c0.n99_adj_3424\ : std_logic;
signal \c0.n77_adj_3415\ : std_logic;
signal \c0.n20801_cascade_\ : std_logic;
signal \c0.n96_adj_3401_cascade_\ : std_logic;
signal \c0.n99\ : std_logic;
signal \c0.n47_adj_3408\ : std_logic;
signal \c0.n18435\ : std_logic;
signal \c0.n42_adj_3064_cascade_\ : std_logic;
signal \c0.n15489_cascade_\ : std_logic;
signal \c0.data_in_frame_15_2\ : std_logic;
signal encoder0_position_31 : std_logic;
signal data_out_frame_6_7 : std_logic;
signal data_in_frame_23_2 : std_logic;
signal \c0.n13_adj_3405_cascade_\ : std_logic;
signal \c0.data_in_frame_27_0\ : std_logic;
signal \c0.n17880_cascade_\ : std_logic;
signal \c0.n19342_cascade_\ : std_logic;
signal \c0.n12035\ : std_logic;
signal \c0.n19496_cascade_\ : std_logic;
signal \c0.n15_adj_3395\ : std_logic;
signal \c0.n19342\ : std_logic;
signal \c0.n36_adj_3307_cascade_\ : std_logic;
signal \c0.n39_adj_3312\ : std_logic;
signal \c0.n29_adj_3148\ : std_logic;
signal \c0.n78_adj_3357\ : std_logic;
signal \c0.n75_cascade_\ : std_logic;
signal \c0.n93_adj_3373_cascade_\ : std_logic;
signal \c0.n96_adj_3419\ : std_logic;
signal \c0.n23_adj_3222_cascade_\ : std_logic;
signal \c0.n76\ : std_logic;
signal \c0.n34\ : std_logic;
signal \c0.n19403\ : std_logic;
signal \c0.data_in_frame_26_6\ : std_logic;
signal \c0.n38_adj_3051\ : std_logic;
signal \c0.n38_adj_3051_cascade_\ : std_logic;
signal \c0.n19496\ : std_logic;
signal \c0.n17947\ : std_logic;
signal \c0.n60_adj_3065\ : std_logic;
signal \c0.n64\ : std_logic;
signal \c0.n51_cascade_\ : std_logic;
signal \c0.n32_adj_3052\ : std_logic;
signal \c0.n45_adj_3284\ : std_logic;
signal \c0.n40_adj_3282\ : std_logic;
signal \c0.n20930\ : std_logic;
signal \c0.n15_adj_3297_cascade_\ : std_logic;
signal \c0.n21003\ : std_logic;
signal \c0.n21_adj_3300_cascade_\ : std_logic;
signal \c0.n23_adj_3304\ : std_logic;
signal \c0.n21247_cascade_\ : std_logic;
signal \c0.n24_adj_3298\ : std_logic;
signal \c0.n14_adj_3354\ : std_logic;
signal data_in_3_4 : std_logic;
signal data_in_0_0 : std_logic;
signal data_in_1_7 : std_logic;
signal \c0.n10_adj_3231\ : std_logic;
signal data_in_2_1 : std_logic;
signal data_in_1_1 : std_logic;
signal \r_Bit_Index_2\ : std_logic;
signal \r_Bit_Index_1\ : std_logic;
signal n4 : std_logic;
signal n4_adj_3579 : std_logic;
signal \c0.n9_adj_3025\ : std_logic;
signal \c0.data_in_frame_2_7\ : std_logic;
signal \c0.n9_adj_3351\ : std_logic;
signal \c0.data_in_frame_4_6\ : std_logic;
signal \c0.n11_adj_3507\ : std_logic;
signal \c0.n13_adj_3504\ : std_logic;
signal \c0.n12131_cascade_\ : std_logic;
signal \c0.n12131\ : std_logic;
signal \c0.n19415\ : std_logic;
signal \c0.n19415_cascade_\ : std_logic;
signal \c0.n54_adj_3502\ : std_logic;
signal \c0.n39_adj_3398\ : std_logic;
signal \c0.n14_adj_3371\ : std_logic;
signal \c0.data_in_frame_3_6\ : std_logic;
signal \c0.n10_adj_3538_cascade_\ : std_logic;
signal \c0.data_in_frame_2_5\ : std_logic;
signal \c0.n22_adj_3356_cascade_\ : std_logic;
signal \c0.n13_adj_3513\ : std_logic;
signal \c0.n23_adj_3021\ : std_logic;
signal \c0.n23_adj_3021_cascade_\ : std_logic;
signal \c0.n26_adj_3114_cascade_\ : std_logic;
signal \c0.n24_adj_3011\ : std_logic;
signal \c0.n22\ : std_logic;
signal \c0.n22_adj_3356\ : std_logic;
signal \c0.n22_adj_3022\ : std_logic;
signal \c0.data_in_frame_12_4\ : std_logic;
signal \c0.n18_adj_3372\ : std_logic;
signal \c0.n88\ : std_logic;
signal \c0.n33\ : std_logic;
signal \c0.n20029\ : std_logic;
signal \c0.n26_adj_3114\ : std_logic;
signal \c0.n30\ : std_logic;
signal \c0.n18422\ : std_logic;
signal \c0.n18422_cascade_\ : std_logic;
signal \c0.n19433_cascade_\ : std_logic;
signal \c0.data_in_frame_10_3\ : std_logic;
signal \c0.n11891_cascade_\ : std_logic;
signal \c0.n44_adj_3117\ : std_logic;
signal \c0.n43_adj_3116\ : std_logic;
signal \c0.n27_adj_3118_cascade_\ : std_logic;
signal \c0.n20052\ : std_logic;
signal \c0.data_in_frame_14_5\ : std_logic;
signal \c0.n11_adj_3340\ : std_logic;
signal \c0.n19916_cascade_\ : std_logic;
signal \c0.n18_adj_3369\ : std_logic;
signal \c0.n19477_cascade_\ : std_logic;
signal \c0.n12_adj_3348_cascade_\ : std_logic;
signal \c0.n21045_cascade_\ : std_logic;
signal \c0.n27_adj_3118\ : std_logic;
signal \c0.n19_adj_3303\ : std_logic;
signal \c0.n12\ : std_logic;
signal \c0.n12_adj_3477\ : std_logic;
signal \c0.data_in_frame_14_4\ : std_logic;
signal \c0.n21110_cascade_\ : std_logic;
signal \c0.n20246\ : std_logic;
signal \c0.data_in_frame_14_3\ : std_logic;
signal \c0.n67_adj_3063\ : std_logic;
signal \c0.n20490\ : std_logic;
signal \c0.n19433\ : std_logic;
signal \c0.n42_adj_3064\ : std_logic;
signal \c0.n12_adj_3518\ : std_logic;
signal \c0.n12_adj_3517_cascade_\ : std_logic;
signal data_in_frame_18_5 : std_logic;
signal \c0.n21_adj_3337\ : std_logic;
signal \c0.n20_adj_3487\ : std_logic;
signal \c0.n20451_cascade_\ : std_logic;
signal \c0.n5_adj_3220\ : std_logic;
signal data_in_frame_18_1 : std_logic;
signal \c0.n27_adj_3529_cascade_\ : std_logic;
signal \c0.n32_adj_3530_cascade_\ : std_logic;
signal \c0.n19244_cascade_\ : std_logic;
signal \c0.n85_adj_3074\ : std_logic;
signal \c0.n85_adj_3074_cascade_\ : std_logic;
signal \c0.n10_adj_3474\ : std_logic;
signal \c0.n20801\ : std_logic;
signal \c0.n49\ : std_logic;
signal \c0.n48_adj_3409\ : std_logic;
signal \c0.n22_adj_3287_cascade_\ : std_logic;
signal \c0.n39_adj_3050\ : std_logic;
signal \c0.n19384\ : std_logic;
signal \c0.n13_adj_3463\ : std_logic;
signal \c0.n10\ : std_logic;
signal \c0.n19384_cascade_\ : std_logic;
signal data_in_frame_16_5 : std_logic;
signal data_in_frame_19_0 : std_logic;
signal \c0.n9_adj_3430_cascade_\ : std_logic;
signal \c0.n10_adj_3445\ : std_logic;
signal \c0.n9_adj_3430\ : std_logic;
signal \c0.n14_adj_3421\ : std_logic;
signal \c0.n18433_cascade_\ : std_logic;
signal \c0.n19511\ : std_logic;
signal \c0.n19511_cascade_\ : std_logic;
signal \c0.n21110\ : std_logic;
signal \c0.n20_adj_3448\ : std_logic;
signal \c0.n20431\ : std_logic;
signal \c0.n64_adj_3512\ : std_logic;
signal data_in_frame_16_4 : std_logic;
signal \c0.n7_adj_3440\ : std_logic;
signal \c0.data_in_frame_13_0\ : std_logic;
signal \c0.n11_adj_3219\ : std_logic;
signal \c0.n13_adj_3221\ : std_logic;
signal data_in_frame_23_3 : std_logic;
signal \c0.n25_adj_3524\ : std_logic;
signal \c0.n21044_cascade_\ : std_logic;
signal \c0.data_in_frame_26_7\ : std_logic;
signal \c0.n16_adj_3109_cascade_\ : std_logic;
signal \c0.n21071\ : std_logic;
signal \c0.n20479\ : std_logic;
signal \c0.n77\ : std_logic;
signal \c0.n34_adj_3096\ : std_logic;
signal \c0.n32_adj_3095\ : std_logic;
signal \c0.n18457_cascade_\ : std_logic;
signal \c0.n23_adj_3222\ : std_logic;
signal \c0.n43_adj_3280_cascade_\ : std_logic;
signal \c0.n41_adj_3281\ : std_logic;
signal \c0.n50_adj_3283\ : std_logic;
signal \c0.n18457\ : std_logic;
signal \c0.n21076\ : std_logic;
signal \c0.n33_adj_3308\ : std_logic;
signal \c0.n18417\ : std_logic;
signal \c0.n18417_cascade_\ : std_logic;
signal \c0.n19_adj_3292\ : std_logic;
signal \c0.data_in_frame_29_4\ : std_logic;
signal \c0.data_in_frame_29_2\ : std_logic;
signal \c0.data_in_frame_29_1\ : std_logic;
signal \c0.data_in_frame_28_1\ : std_logic;
signal \c0.data_in_frame_28_0\ : std_logic;
signal \c0.n20324\ : std_logic;
signal \c0.n14_adj_3349\ : std_logic;
signal \c0.n7_adj_3078\ : std_logic;
signal \c0.n17880\ : std_logic;
signal \c0.n26_adj_3523\ : std_logic;
signal data_in_0_4 : std_logic;
signal n20896 : std_logic;
signal \c0.n12085\ : std_logic;
signal \c0.n11865\ : std_logic;
signal \c0.n12085_cascade_\ : std_logic;
signal \c0.n6495\ : std_logic;
signal data_in_2_4 : std_logic;
signal data_in_1_4 : std_logic;
signal \c0.n6_adj_3343\ : std_logic;
signal \c0.data_out_frame_28_7\ : std_logic;
signal n8112 : std_logic;
signal \c0.data_in_frame_4_3\ : std_logic;
signal \c0.data_in_frame_4_2\ : std_logic;
signal \c0.data_in_frame_6_4\ : std_logic;
signal \c0.n13_adj_3496_cascade_\ : std_logic;
signal \c0.data_in_frame_2_2\ : std_logic;
signal data_in_frame_0_0 : std_logic;
signal \c0.n19277\ : std_logic;
signal \c0.data_in_frame_2_0\ : std_logic;
signal \c0.n8_adj_3397\ : std_logic;
signal \c0.n11833_cascade_\ : std_logic;
signal \c0.n92_cascade_\ : std_logic;
signal \c0.n80\ : std_logic;
signal \c0.n19196\ : std_logic;
signal \c0.data_in_frame_4_5\ : std_logic;
signal \c0.n54\ : std_logic;
signal \c0.n90\ : std_logic;
signal \c0.n98\ : std_logic;
signal \c0.n21277\ : std_logic;
signal \c0.n4_adj_3406\ : std_logic;
signal \c0.n14_adj_3476_cascade_\ : std_logic;
signal \c0.data_in_frame_7_3\ : std_logic;
signal \c0.n19508\ : std_logic;
signal \c0.n10_adj_3538\ : std_logic;
signal \c0.n85\ : std_logic;
signal \c0.n37\ : std_logic;
signal \c0.n67_cascade_\ : std_logic;
signal \c0.n96\ : std_logic;
signal \c0.n83\ : std_logic;
signal \c0.n40_adj_3032\ : std_logic;
signal \c0.n100_cascade_\ : std_logic;
signal \c0.n102\ : std_logic;
signal \c0.n4_adj_3009\ : std_logic;
signal \c0.n21_adj_3010\ : std_logic;
signal \c0.n28_adj_3023\ : std_logic;
signal \c0.n17_adj_3508\ : std_logic;
signal \c0.n19966\ : std_logic;
signal \c0.n30_adj_3075\ : std_logic;
signal \c0.n32_adj_3077_cascade_\ : std_logic;
signal \c0.n19372\ : std_logic;
signal \c0.n21047_cascade_\ : std_logic;
signal \c0.n42_adj_3111\ : std_logic;
signal \c0.data_in_frame_3_0\ : std_logic;
signal \c0.data_in_frame_2_6\ : std_logic;
signal \c0.n10_adj_3014_cascade_\ : std_logic;
signal \c0.n40\ : std_logic;
signal \c0.n16_adj_3218_cascade_\ : std_logic;
signal \c0.data_in_frame_12_2\ : std_logic;
signal \c0.n7_adj_3491\ : std_logic;
signal \c0.n30_adj_3531\ : std_logic;
signal \c0.n12_adj_3034\ : std_logic;
signal \c0.n31_adj_3532\ : std_logic;
signal \c0.n11537\ : std_logic;
signal \c0.data_in_frame_15_6\ : std_logic;
signal \c0.n16_adj_3481_cascade_\ : std_logic;
signal \c0.n11815_cascade_\ : std_logic;
signal \c0.n19291\ : std_logic;
signal data_in_frame_16_1 : std_logic;
signal \c0.n12056_cascade_\ : std_logic;
signal \c0.n12_adj_3249\ : std_logic;
signal \c0.n12_adj_3249_cascade_\ : std_logic;
signal \c0.n12056\ : std_logic;
signal \c0.n19301\ : std_logic;
signal \c0.n19301_cascade_\ : std_logic;
signal \c0.n31_adj_3126_cascade_\ : std_logic;
signal \c0.n19427\ : std_logic;
signal \c0.n19551\ : std_logic;
signal \c0.n27_adj_3455\ : std_logic;
signal \c0.n46_cascade_\ : std_logic;
signal \c0.n46\ : std_logic;
signal \c0.n8\ : std_logic;
signal \c0.n84\ : std_logic;
signal \c0.n19824_cascade_\ : std_logic;
signal \c0.n29\ : std_logic;
signal \c0.n18_adj_3360_cascade_\ : std_logic;
signal \c0.n32_adj_3362_cascade_\ : std_logic;
signal \c0.n20112_cascade_\ : std_logic;
signal \c0.data_in_frame_13_1\ : std_logic;
signal \c0.n18398_cascade_\ : std_logic;
signal \c0.n37_adj_3390_cascade_\ : std_logic;
signal \c0.n37_adj_3390\ : std_logic;
signal \c0.n60_adj_3368_cascade_\ : std_logic;
signal \c0.n51_adj_3376\ : std_logic;
signal \c0.n19916\ : std_logic;
signal \c0.n18443\ : std_logic;
signal \c0.n39_adj_3334\ : std_logic;
signal \c0.n19_adj_3336\ : std_logic;
signal \c0.n39_adj_3334_cascade_\ : std_logic;
signal \c0.n25_adj_3431\ : std_logic;
signal \c0.n42_adj_3367\ : std_logic;
signal \c0.n43_adj_3386\ : std_logic;
signal \c0.n40_adj_3366\ : std_logic;
signal \c0.n30_adj_3429\ : std_logic;
signal \c0.n35_adj_3274_cascade_\ : std_logic;
signal \c0.n59\ : std_logic;
signal \c0.n30_adj_3392\ : std_logic;
signal \c0.n21047\ : std_logic;
signal \c0.n12_adj_3049\ : std_logic;
signal \c0.n91\ : std_logic;
signal \c0.n35_adj_3274\ : std_logic;
signal \c0.n17_adj_3451\ : std_logic;
signal \c0.n20403\ : std_logic;
signal \c0.n22_adj_3450\ : std_logic;
signal \c0.n24_adj_3427_cascade_\ : std_logic;
signal \c0.data_in_frame_17_0\ : std_logic;
signal \c0.n32_adj_3057_cascade_\ : std_logic;
signal \c0.n33_adj_3289\ : std_logic;
signal \c0.n10_adj_3555\ : std_logic;
signal \c0.n4_adj_3522\ : std_logic;
signal \c0.n55_adj_3273\ : std_logic;
signal \c0.n19514\ : std_logic;
signal \c0.n20965_cascade_\ : std_logic;
signal \c0.n40_adj_3323\ : std_logic;
signal \c0.data_in_frame_27_3\ : std_logic;
signal \c0.n20336_cascade_\ : std_logic;
signal \c0.n61_adj_3387\ : std_logic;
signal \c0.n63_adj_3391\ : std_logic;
signal \c0.n21034_cascade_\ : std_logic;
signal \c0.n12134\ : std_logic;
signal \c0.n58_adj_3381\ : std_logic;
signal \c0.n43_adj_3330\ : std_logic;
signal \c0.n50_adj_3331\ : std_logic;
signal \c0.n35_adj_3266\ : std_logic;
signal \c0.n33_adj_3097\ : std_logic;
signal \c0.n9_adj_3240\ : std_logic;
signal \c0.n20112\ : std_logic;
signal \c0.n32_adj_3236\ : std_logic;
signal \c0.n28_adj_3245\ : std_logic;
signal \c0.n27_adj_3241_cascade_\ : std_logic;
signal \c0.n13_adj_3244\ : std_logic;
signal \c0.n19_adj_3135\ : std_logic;
signal \c0.n19_adj_3135_cascade_\ : std_logic;
signal \c0.n24_adj_3134\ : std_logic;
signal \c0.n86\ : std_logic;
signal \c0.n22_adj_3136_cascade_\ : std_logic;
signal \c0.n11936_cascade_\ : std_logic;
signal \c0.data_in_frame_27_4\ : std_logic;
signal \c0.data_in_frame_27_5\ : std_logic;
signal \c0.n17_adj_3318\ : std_logic;
signal \c0.n11936\ : std_logic;
signal \c0.n12_adj_3141\ : std_logic;
signal data_in_frame_24_6 : std_logic;
signal data_in_frame_24_4 : std_logic;
signal \c0.n19465_cascade_\ : std_logic;
signal \c0.n17\ : std_logic;
signal \c0.n21044\ : std_logic;
signal \c0.n19703\ : std_logic;
signal \c0.n19703_cascade_\ : std_logic;
signal \c0.n44_adj_3278\ : std_logic;
signal \c0.data_in_frame_25_1\ : std_logic;
signal \c0.n18377\ : std_logic;
signal \c0.data_in_frame_25_2\ : std_logic;
signal \c0.data_in_frame_25_3\ : std_logic;
signal \c0.n19400\ : std_logic;
signal \c0.data_in_frame_26_5\ : std_logic;
signal \c0.n17840\ : std_logic;
signal data_in_3_0 : std_logic;
signal \c0.n12_adj_3498\ : std_logic;
signal \c0.FRAME_MATCHER_i_5\ : std_logic;
signal \c0.n6_adj_3149\ : std_logic;
signal \c0.data_in_frame_8_6\ : std_logic;
signal \c0.data_in_frame_4_0\ : std_logic;
signal \c0.n17_adj_3113\ : std_logic;
signal \c0.n5_adj_3030\ : std_logic;
signal \c0.n60_cascade_\ : std_logic;
signal \c0.n93\ : std_logic;
signal \c0.data_in_frame_6_1\ : std_logic;
signal \c0.n5_adj_3028\ : std_logic;
signal \c0.n19443\ : std_logic;
signal \c0.n11687\ : std_logic;
signal \c0.n20313\ : std_logic;
signal \c0.n8_adj_3066_cascade_\ : std_logic;
signal \c0.n19170\ : std_logic;
signal \c0.n19170_cascade_\ : std_logic;
signal \c0.data_in_frame_8_2\ : std_logic;
signal \c0.n21_adj_3053\ : std_logic;
signal \c0.n21\ : std_logic;
signal \c0.data_in_frame_5_4\ : std_logic;
signal \c0.n25\ : std_logic;
signal \c0.n89\ : std_logic;
signal \c0.data_in_frame_3_1\ : std_logic;
signal data_in_frame_0_5 : std_logic;
signal \c0.n33_adj_3088\ : std_logic;
signal \c0.n15_adj_3545\ : std_logic;
signal \c0.n24_adj_3013\ : std_logic;
signal \c0.data_in_frame_3_3\ : std_logic;
signal \c0.data_in_frame_3_2\ : std_logic;
signal \data_out_frame_29__3__N_647\ : std_logic;
signal \c0.n29_adj_3216\ : std_logic;
signal \c0.n78\ : std_logic;
signal \c0.n37_adj_3215\ : std_logic;
signal \c0.n29_adj_3216_cascade_\ : std_logic;
signal \c0.n44_adj_3217\ : std_logic;
signal \c0.n36_adj_3212_cascade_\ : std_logic;
signal \c0.n41_adj_3213\ : std_logic;
signal \c0.n20340\ : std_logic;
signal \c0.n11651_cascade_\ : std_logic;
signal \c0.n27_adj_3082\ : std_logic;
signal \c0.n11800\ : std_logic;
signal \c0.n31\ : std_logic;
signal \c0.n37_adj_3153\ : std_logic;
signal \c0.n35_adj_3233\ : std_logic;
signal \c0.n60\ : std_logic;
signal \c0.n52_adj_3223_cascade_\ : std_logic;
signal \c0.n60_adj_3503\ : std_logic;
signal \c0.n52_adj_3402\ : std_logic;
signal \c0.data_in_frame_7_4\ : std_logic;
signal \c0.n20391\ : std_logic;
signal \c0.n4\ : std_logic;
signal \c0.n12026\ : std_logic;
signal \c0.n5\ : std_logic;
signal \c0.n4_cascade_\ : std_logic;
signal \c0.data_in_frame_11_4\ : std_logic;
signal \c0.data_in_frame_10_0\ : std_logic;
signal \c0.data_in_frame_21_0\ : std_logic;
signal \c0.n16_adj_3218\ : std_logic;
signal \c0.n48\ : std_logic;
signal \c0.data_in_frame_5_1\ : std_logic;
signal \c0.n20224\ : std_logic;
signal \c0.n5_adj_3549\ : std_logic;
signal \c0.data_in_frame_4_7\ : std_logic;
signal \c0.n11613\ : std_logic;
signal \c0.data_in_frame_17_6\ : std_logic;
signal data_in_frame_18_0 : std_logic;
signal \c0.n11613_cascade_\ : std_logic;
signal \c0.n19477\ : std_logic;
signal \c0.n17_adj_3482\ : std_logic;
signal \c0.data_in_frame_13_6\ : std_logic;
signal \c0.data_in_frame_13_5\ : std_logic;
signal \c0.n20826\ : std_logic;
signal \c0.n54_adj_3234\ : std_logic;
signal \c0.n43_adj_3232_cascade_\ : std_logic;
signal \c0.n17849\ : std_logic;
signal \c0.n49_adj_3237\ : std_logic;
signal \c0.n7_adj_3225_cascade_\ : std_logic;
signal \c0.data_in_frame_15_4\ : std_logic;
signal \c0.n7_adj_3225\ : std_logic;
signal \c0.n44_adj_3226\ : std_logic;
signal \c0.data_in_frame_10_4\ : std_logic;
signal \c0.data_in_frame_8_1\ : std_logic;
signal \c0.n41_adj_3365\ : std_logic;
signal \c0.n22_adj_3287\ : std_logic;
signal \c0.n47_adj_3286_cascade_\ : std_logic;
signal \c0.n51_adj_3290\ : std_logic;
signal \c0.n52_adj_3288_cascade_\ : std_logic;
signal \c0.n6_adj_3291\ : std_logic;
signal \c0.data_in_frame_11_6\ : std_logic;
signal \c0.n19909_cascade_\ : std_logic;
signal \c0.n87\ : std_logic;
signal \c0.n6_adj_3137\ : std_logic;
signal \c0.n35_adj_3098\ : std_logic;
signal \c0.n19909\ : std_logic;
signal \c0.n19223\ : std_logic;
signal \c0.n12218\ : std_logic;
signal \c0.n7_adj_3047_cascade_\ : std_logic;
signal \c0.n28_adj_3059_cascade_\ : std_logic;
signal \c0.n36_adj_3452\ : std_logic;
signal \c0.n47\ : std_logic;
signal \c0.n17819\ : std_logic;
signal \c0.n20321\ : std_logic;
signal \c0.n19824\ : std_logic;
signal \c0.n12_adj_3469\ : std_logic;
signal \c0.n29_adj_3461_cascade_\ : std_logic;
signal \c0.n25_adj_3035\ : std_logic;
signal \c0.n23_adj_3364\ : std_logic;
signal \c0.n24_adj_3335\ : std_logic;
signal \c0.n36_adj_3470_cascade_\ : std_logic;
signal \c0.n22_adj_3341\ : std_logic;
signal \c0.n11_adj_3124_cascade_\ : std_logic;
signal \c0.n32_adj_3465\ : std_logic;
signal \c0.n33_adj_3315\ : std_logic;
signal \c0.n49_adj_3316\ : std_logic;
signal \c0.n35_adj_3317\ : std_logic;
signal \c0.data_in_frame_17_1\ : std_logic;
signal \c0.n17871\ : std_logic;
signal \c0.n22_adj_3363\ : std_logic;
signal \c0.n22_adj_3363_cascade_\ : std_logic;
signal \c0.n30_adj_3468\ : std_logic;
signal \c0.n65\ : std_logic;
signal \c0.n70_adj_3087_cascade_\ : std_logic;
signal \c0.n20339\ : std_logic;
signal \c0.n27_adj_3311\ : std_logic;
signal \c0.n7_adj_3094\ : std_logic;
signal \c0.n20_adj_3293\ : std_logic;
signal \c0.n33_adj_3279\ : std_logic;
signal \c0.n30_adj_3295\ : std_logic;
signal \c0.n32_adj_3294_cascade_\ : std_logic;
signal \c0.n21075\ : std_logic;
signal \c0.n7_adj_3079\ : std_logic;
signal \c0.n29_adj_3299\ : std_logic;
signal \c0.n19_adj_3320\ : std_logic;
signal \c0.n20336\ : std_logic;
signal \c0.n18379\ : std_logic;
signal \c0.n21034\ : std_logic;
signal \c0.n57\ : std_logic;
signal \c0.n24_adj_3427\ : std_logic;
signal \c0.n11714\ : std_logic;
signal \c0.n22_adj_3296\ : std_logic;
signal \c0.n19159_cascade_\ : std_logic;
signal \c0.n11632\ : std_logic;
signal \c0.n19159\ : std_logic;
signal \c0.data_in_frame_28_7\ : std_logic;
signal \c0.n79\ : std_logic;
signal \c0.n10_adj_3207\ : std_logic;
signal \c0.n11_adj_3206\ : std_logic;
signal \c0.n11776_cascade_\ : std_logic;
signal \c0.n6_adj_3319\ : std_logic;
signal data_in_frame_24_7 : std_logic;
signal \c0.n12206\ : std_logic;
signal \c0.n19268\ : std_logic;
signal \c0.n19268_cascade_\ : std_logic;
signal \c0.n20_adj_3301\ : std_logic;
signal \c0.n7_adj_3054\ : std_logic;
signal \c0.n11601\ : std_logic;
signal \c0.n19764\ : std_logic;
signal \c0.n42_adj_3055\ : std_logic;
signal \c0.n11815\ : std_logic;
signal \c0.n4_adj_3100\ : std_logic;
signal \c0.data_in_frame_25_0\ : std_logic;
signal \c0.n19436\ : std_logic;
signal data_in_frame_22_4 : std_logic;
signal \c0.n19436_cascade_\ : std_logic;
signal \c0.n11776\ : std_logic;
signal \c0.n6_adj_3112\ : std_logic;
signal \c0.n19151\ : std_logic;
signal \c0.n20933\ : std_logic;
signal rx_data_ready : std_logic;
signal data_in_3_6 : std_logic;
signal data_in_2_6 : std_logic;
signal \c0.n25_adj_3048\ : std_logic;
signal \c0.n19312\ : std_logic;
signal \c0.n20512\ : std_logic;
signal \c0.n19202\ : std_logic;
signal \c0.n12_adj_3210_cascade_\ : std_logic;
signal \c0.n18433\ : std_logic;
signal \c0.n17834\ : std_logic;
signal \c0.n21767\ : std_logic;
signal data_in_frame_22_6 : std_logic;
signal data_in_frame_23_0 : std_logic;
signal data_in_frame_23_4 : std_logic;
signal n19126 : std_logic;
signal \c0.data_in_frame_11_0\ : std_logic;
signal \c0.data_in_frame_2_1\ : std_logic;
signal \c0.n34_adj_3326\ : std_logic;
signal \c0.n13_adj_3344\ : std_logic;
signal \c0.n23_adj_3076\ : std_logic;
signal \c0.n19424\ : std_logic;
signal \c0.n7_adj_3029\ : std_logic;
signal data_in_frame_0_4 : std_logic;
signal \c0.data_in_frame_2_3\ : std_logic;
signal \c0.data_in_frame_4_4\ : std_logic;
signal \c0.n8_adj_3345\ : std_logic;
signal \c0.n7_adj_3520\ : std_logic;
signal \c0.n9_adj_3346\ : std_logic;
signal \c0.n8_adj_3345_cascade_\ : std_logic;
signal \c0.n11626_cascade_\ : std_logic;
signal \c0.data_in_frame_8_7\ : std_logic;
signal data_in_frame_1_1 : std_logic;
signal \c0.n19970\ : std_logic;
signal \c0.n6_adj_3501\ : std_logic;
signal \c0.data_in_frame_6_3\ : std_logic;
signal \c0.n11478_cascade_\ : std_logic;
signal \c0.n81\ : std_logic;
signal data_in_frame_1_6 : std_logic;
signal \c0.n11526\ : std_logic;
signal \c0.data_in_frame_6_5\ : std_logic;
signal \c0.n11549\ : std_logic;
signal \c0.n11651\ : std_logic;
signal \c0.n27_adj_3457\ : std_logic;
signal data_in_frame_1_7 : std_logic;
signal \c0.n12_adj_3378\ : std_logic;
signal \c0.n11626\ : std_logic;
signal \c0.n21_adj_3205\ : std_logic;
signal \c0.n28_adj_3428\ : std_logic;
signal data_in_frame_1_5 : std_logic;
signal \c0.n7_adj_3509\ : std_logic;
signal \c0.n7_adj_3509_cascade_\ : std_logic;
signal \c0.n10_adj_3012\ : std_logic;
signal \c0.n45\ : std_logic;
signal \c0.data_in_frame_4_1\ : std_logic;
signal data_in_frame_0_6 : std_logic;
signal data_in_frame_1_0 : std_logic;
signal \c0.n20341\ : std_logic;
signal \c0.n58_adj_3497\ : std_logic;
signal \c0.n56_adj_3505\ : std_logic;
signal \c0.n64_adj_3506\ : std_logic;
signal \c0.n19217\ : std_logic;
signal \c0.n4_adj_3036_cascade_\ : std_logic;
signal \c0.n57_adj_3499\ : std_logic;
signal \c0.n6_adj_3019\ : std_logic;
signal \c0.data_in_frame_7_5\ : std_logic;
signal \c0.n6_adj_3019_cascade_\ : std_logic;
signal \c0.n20386\ : std_logic;
signal \c0.data_in_frame_9_6\ : std_logic;
signal \c0.data_in_frame_3_7\ : std_logic;
signal \c0.data_in_frame_5_5\ : std_logic;
signal \c0.data_in_frame_5_3\ : std_logic;
signal n11461 : std_logic;
signal \c0.n23\ : std_logic;
signal \c0.n51_adj_3426\ : std_logic;
signal n15645 : std_logic;
signal \r_Rx_Data\ : std_logic;
signal n11466 : std_logic;
signal \c0.data_in_frame_13_7\ : std_logic;
signal \c0.n13_adj_3541\ : std_logic;
signal \c0.data_in_frame_13_2\ : std_logic;
signal \c0.data_in_frame_9_5\ : std_logic;
signal \c0.n9_adj_3211\ : std_logic;
signal data_in_frame_0_1 : std_logic;
signal \c0.n17_adj_3544\ : std_logic;
signal \c0.data_in_frame_9_1\ : std_logic;
signal \c0.n11858_cascade_\ : std_logic;
signal \c0.n19446\ : std_logic;
signal \c0.n19446_cascade_\ : std_logic;
signal \c0.data_out_frame_0__7__N_1537\ : std_logic;
signal \c0.n11982\ : std_logic;
signal \c0.n33_adj_3209_cascade_\ : std_logic;
signal \c0.n5598\ : std_logic;
signal \c0.data_in_frame_17_7\ : std_logic;
signal \c0.n9_adj_3350\ : std_logic;
signal \c0.n29_adj_3533\ : std_logic;
signal \c0.n33_adj_3209\ : std_logic;
signal \c0.n12209\ : std_logic;
signal \c0.n9_adj_3027\ : std_logic;
signal \c0.n45_adj_3224\ : std_logic;
signal \c0.data_in_frame_7_6\ : std_logic;
signal \c0.n15\ : std_logic;
signal \c0.n5753\ : std_logic;
signal \c0.data_in_frame_14_0\ : std_logic;
signal \c0.data_in_frame_12_0\ : std_logic;
signal \c0.n20055\ : std_logic;
signal \c0.n20_adj_3536_cascade_\ : std_logic;
signal \c0.n12_adj_3558_cascade_\ : std_logic;
signal \c0.data_in_frame_8_5\ : std_logic;
signal \c0.data_in_frame_12_7\ : std_logic;
signal \c0.n5_adj_3031\ : std_logic;
signal \c0.n19359_cascade_\ : std_logic;
signal \c0.data_in_frame_8_4\ : std_logic;
signal \c0.n11478\ : std_logic;
signal \c0.n19199\ : std_logic;
signal \c0.data_in_frame_10_5\ : std_logic;
signal \c0.n19199_cascade_\ : std_logic;
signal \c0.n19_adj_3540\ : std_logic;
signal \c0.data_in_frame_14_1\ : std_logic;
signal \c0.data_in_frame_15_7\ : std_logic;
signal \c0.data_in_frame_14_2\ : std_logic;
signal \c0.data_in_frame_7_2\ : std_logic;
signal \c0.n20981\ : std_logic;
signal \c0.n25_adj_3157\ : std_logic;
signal \c0.n69\ : std_logic;
signal \c0.n28_adj_3059\ : std_logic;
signal \c0.n38_adj_3058_cascade_\ : std_logic;
signal \c0.n32_adj_3060\ : std_logic;
signal \c0.n8_adj_3061_cascade_\ : std_logic;
signal \c0.n52\ : std_logic;
signal \c0.n8_adj_3061\ : std_logic;
signal \c0.n43_adj_3285_cascade_\ : std_logic;
signal \c0.n53\ : std_logic;
signal \c0.n4_adj_3123\ : std_logic;
signal data_in_frame_16_7 : std_logic;
signal \c0.data_in_frame_12_5\ : std_logic;
signal \c0.n12_adj_3554_cascade_\ : std_logic;
signal \c0.n20151\ : std_logic;
signal \c0.n20542\ : std_logic;
signal \c0.n20542_cascade_\ : std_logic;
signal \c0.n45_adj_3423\ : std_logic;
signal \c0.n25_adj_3510_cascade_\ : std_logic;
signal \c0.n58_adj_3511\ : std_logic;
signal \c0.n20085\ : std_logic;
signal \c0.n19244\ : std_logic;
signal \c0.n88_adj_3422\ : std_logic;
signal \c0.n25_adj_3510\ : std_logic;
signal \c0.n56\ : std_logic;
signal \c0.n44_adj_3125\ : std_logic;
signal \c0.n11_adj_3124\ : std_logic;
signal \c0.n48_adj_3313\ : std_logic;
signal \c0.n35_cascade_\ : std_logic;
signal \c0.n67_adj_3092\ : std_logic;
signal \c0.n43_adj_3089\ : std_logic;
signal \c0.n41_adj_3085\ : std_logic;
signal \c0.n42_adj_3086\ : std_logic;
signal \c0.n60_adj_3127\ : std_logic;
signal \c0.n55_adj_3128_cascade_\ : std_logic;
signal \c0.n19749\ : std_logic;
signal \c0.n58\ : std_logic;
signal \c0.n16_adj_3489\ : std_logic;
signal \c0.n31_adj_3126\ : std_logic;
signal \c0.n10_adj_3425_cascade_\ : std_logic;
signal \c0.n42_adj_3130\ : std_logic;
signal \c0.n92_adj_3272\ : std_logic;
signal \c0.n39_adj_3269\ : std_logic;
signal \c0.n36_adj_3275\ : std_logic;
signal \c0.n38_adj_3270\ : std_logic;
signal \c0.n39_adj_3269_cascade_\ : std_logic;
signal \c0.n37_adj_3268\ : std_logic;
signal \c0.n94_adj_3375\ : std_logic;
signal \c0.n92_adj_3377_cascade_\ : std_logic;
signal \c0.n91_adj_3389\ : std_logic;
signal \c0.n100_adj_3420\ : std_logic;
signal \c0.n11942\ : std_logic;
signal \c0.n12_adj_3208\ : std_logic;
signal \c0.n10_adj_3425\ : std_logic;
signal \c0.n82\ : std_logic;
signal \c0.n93_adj_3385\ : std_logic;
signal \c0.n32_adj_3057\ : std_logic;
signal \c0.n62\ : std_logic;
signal \c0.n68\ : std_logic;
signal \c0.n19502\ : std_logic;
signal \c0.n20_adj_3536\ : std_logic;
signal \c0.n23_adj_3534\ : std_logic;
signal \c0.n40_adj_3374\ : std_logic;
signal \c0.n38_adj_3062_cascade_\ : std_logic;
signal \c0.n39_adj_3384\ : std_logic;
signal \c0.n93_adj_3329\ : std_logic;
signal \c0.data_in_frame_8_3\ : std_logic;
signal \c0.n19505\ : std_logic;
signal \c0.n26_adj_3537\ : std_logic;
signal \c0.n20917_cascade_\ : std_logic;
signal \c0.n19524\ : std_logic;
signal \c0.n6_adj_3433_cascade_\ : std_logic;
signal \c0.n18375_cascade_\ : std_logic;
signal \c0.n38_adj_3062\ : std_logic;
signal \c0.n83_adj_3442\ : std_logic;
signal data_in_frame_18_7 : std_logic;
signal \c0.n12052\ : std_logic;
signal \c0.n19_adj_3056\ : std_logic;
signal \c0.n19_adj_3056_cascade_\ : std_logic;
signal \c0.n21045\ : std_logic;
signal \c0.n29_adj_3454\ : std_logic;
signal \c0.n18398\ : std_logic;
signal \c0.n6_adj_3239\ : std_logic;
signal data_in_frame_22_2 : std_logic;
signal \c0.n19354\ : std_logic;
signal data_in_frame_22_7 : std_logic;
signal data_in_frame_22_3 : std_logic;
signal data_in_frame_24_0 : std_logic;
signal \c0.data_in_frame_26_2\ : std_logic;
signal \c0.n18431\ : std_logic;
signal \c0.n15701\ : std_logic;
signal \c0.n7_adj_3047\ : std_logic;
signal \c0.n20965\ : std_logic;
signal \c0.data_in_frame_26_0\ : std_logic;
signal \c0.data_in_frame_27_1\ : std_logic;
signal \c0.data_in_frame_27_2\ : std_logic;
signal \c0.data_in_frame_28_2\ : std_logic;
signal \c0.n20709\ : std_logic;
signal \c0.n17942\ : std_logic;
signal \c0.n77_adj_3396_cascade_\ : std_logic;
signal \c0.n90_adj_3400\ : std_logic;
signal \c0.data_in_frame_25_7\ : std_logic;
signal \c0.data_in_frame_25_5\ : std_logic;
signal \c0.data_in_frame_25_4\ : std_logic;
signal \c0.n19214_cascade_\ : std_logic;
signal data_in_frame_24_5 : std_logic;
signal \c0.n12_adj_3214\ : std_logic;
signal \c0.data_in_frame_25_6\ : std_logic;
signal \c0.n5784\ : std_logic;
signal \c0.n11833\ : std_logic;
signal \c0.n19456\ : std_logic;
signal \c0.n5595\ : std_logic;
signal n2108 : std_logic;
signal \c0.n6_adj_3140\ : std_logic;
signal \c0.data_in_frame_6_0\ : std_logic;
signal \c0.data_in_frame_6_2\ : std_logic;
signal data_in_frame_1_2 : std_logic;
signal \c0.n9_adj_3101\ : std_logic;
signal \FRAME_MATCHER_i_0\ : std_logic;
signal \c0.FRAME_MATCHER_i_1\ : std_logic;
signal \c0.FRAME_MATCHER_i_2\ : std_logic;
signal n19100 : std_logic;
signal \c0.n20095\ : std_logic;
signal data_in_frame_0_3 : std_logic;
signal \c0.n5240\ : std_logic;
signal \c0.n7_cascade_\ : std_logic;
signal \c0.n9_adj_3038\ : std_logic;
signal \c0.data_in_frame_6_7\ : std_logic;
signal \c0.n19098\ : std_logic;
signal \c0.n9_adj_3251\ : std_logic;
signal \c0.data_in_frame_3_4\ : std_logic;
signal \c0.n12_adj_2998\ : std_logic;
signal \c0.n19176\ : std_logic;
signal \c0.n11953\ : std_logic;
signal \c0.data_in_frame_5_2\ : std_logic;
signal data_in_frame_1_3 : std_logic;
signal \c0.n55_adj_3500\ : std_logic;
signal data_in_frame_0_2 : std_logic;
signal \c0.n7\ : std_logic;
signal \c0.n19241\ : std_logic;
signal \c0.data_in_frame_2_4\ : std_logic;
signal data_in_frame_1_4 : std_logic;
signal \c0.n6_adj_3037\ : std_logic;
signal \c0.data_in_frame_5_7\ : std_logic;
signal \c0.n4_adj_3036\ : std_logic;
signal \c0.n6_adj_3037_cascade_\ : std_logic;
signal \c0.data_in_frame_3_5\ : std_logic;
signal \c0.n19560\ : std_logic;
signal \c0.data_out_frame_0__7__N_1540\ : std_logic;
signal \c0.data_in_frame_6_6\ : std_logic;
signal \c0.n19258\ : std_logic;
signal \c0.data_in_frame_8_0\ : std_logic;
signal \c0.data_in_frame_7_7\ : std_logic;
signal \c0.data_in_frame_5_6\ : std_logic;
signal \c0.n8_adj_3020\ : std_logic;
signal \c0.data_in_frame_13_3\ : std_logic;
signal \c0.data_in_frame_9_2\ : std_logic;
signal \c0.n19115\ : std_logic;
signal \c0.data_in_frame_9_3\ : std_logic;
signal \c0.data_in_frame_11_5\ : std_logic;
signal \c0.n5_adj_3043\ : std_logic;
signal \c0.data_in_frame_7_1\ : std_logic;
signal \c0.data_in_frame_9_0\ : std_logic;
signal \c0.data_in_frame_11_3\ : std_logic;
signal \c0.data_in_frame_13_4\ : std_logic;
signal \c0.n11_adj_3492\ : std_logic;
signal \c0.n11_adj_3492_cascade_\ : std_logic;
signal data_in_frame_16_0 : std_logic;
signal \c0.n20_adj_3527\ : std_logic;
signal \c0.data_in_frame_11_1\ : std_logic;
signal \c0.n19229\ : std_logic;
signal \c0.data_in_frame_11_2\ : std_logic;
signal \c0.n19134\ : std_logic;
signal \c0.data_in_frame_10_7\ : std_logic;
signal \c0.n19131\ : std_logic;
signal \c0.data_in_frame_11_7\ : std_logic;
signal \c0.n15489\ : std_logic;
signal \c0.n19140\ : std_logic;
signal \c0.data_in_frame_15_5\ : std_logic;
signal \c0.n9_adj_3552_cascade_\ : std_logic;
signal data_in_frame_18_3 : std_logic;
signal n19129 : std_logic;
signal data_in_frame_18_4 : std_logic;
signal \c0.data_in_frame_12_1\ : std_logic;
signal \c0.n7_adj_3000\ : std_logic;
signal \c0.n19430\ : std_logic;
signal \c0.n7_adj_3000_cascade_\ : std_logic;
signal data_in_frame_16_3 : std_logic;
signal \c0.n6\ : std_logic;
signal \c0.n19187\ : std_logic;
signal \c0.n46_adj_3443\ : std_logic;
signal \c0.data_in_frame_15_0\ : std_logic;
signal \c0.n40_adj_3413\ : std_logic;
signal \c0.n45_adj_3138\ : std_logic;
signal \c0.n19381\ : std_logic;
signal \c0.data_in_frame_7_0\ : std_logic;
signal \c0.n7_adj_3355\ : std_logic;
signal \c0.data_in_frame_17_5\ : std_logic;
signal \c0.n11590\ : std_logic;
signal \c0.n14_adj_3449\ : std_logic;
signal rx_data_0 : std_logic;
signal \c0.data_in_frame_15_1\ : std_logic;
signal \c0.data_in_frame_14_7\ : std_logic;
signal \c0.data_in_frame_14_6\ : std_logic;
signal \c0.n19554\ : std_logic;
signal \c0.data_in_frame_17_4\ : std_logic;
signal \c0.n18_adj_3235\ : std_logic;
signal \c0.data_in_frame_15_3\ : std_logic;
signal \c0.n10_adj_3483\ : std_logic;
signal \c0.n18420\ : std_logic;
signal \c0.n19251\ : std_logic;
signal \c0.n7_adj_3347\ : std_logic;
signal \c0.data_in_frame_10_6\ : std_logic;
signal \c0.n19359\ : std_logic;
signal \c0.data_in_frame_12_6\ : std_logic;
signal \c0.n22_adj_3535\ : std_logic;
signal \c0.data_in_frame_20_1\ : std_logic;
signal \c0.n12_adj_3265\ : std_logic;
signal \c0.data_in_frame_12_3\ : std_logic;
signal data_in_frame_19_2 : std_logic;
signal data_in_frame_19_5 : std_logic;
signal data_in_frame_19_1 : std_logic;
signal \c0.n6166\ : std_logic;
signal n19130 : std_logic;
signal data_in_frame_16_2 : std_logic;
signal \c0.data_in_frame_28_5\ : std_logic;
signal \c0.n19111\ : std_logic;
signal \c0.data_in_frame_29_3\ : std_logic;
signal \c0.n12_adj_3006\ : std_logic;
signal \c0.data_in_frame_29_5\ : std_logic;
signal \c0.n15_adj_3432\ : std_logic;
signal \c0.n20503\ : std_logic;
signal data_in_frame_23_1 : std_logic;
signal \c0.n20503_cascade_\ : std_logic;
signal \c0.n12_adj_3494\ : std_logic;
signal \c0.n27_adj_3399\ : std_logic;
signal \c0.data_in_frame_28_3\ : std_logic;
signal \c0.n27_adj_3399_cascade_\ : std_logic;
signal \c0.data_in_frame_26_1\ : std_logic;
signal \c0.n78_adj_3414\ : std_logic;
signal data_in_frame_23_6 : std_logic;
signal data_in_frame_23_5 : std_logic;
signal \c0.n19487\ : std_logic;
signal data_in_frame_23_7 : std_logic;
signal \c0.n11971\ : std_logic;
signal \c0.n19484\ : std_logic;
signal \c0.n7_adj_3072_cascade_\ : std_logic;
signal \c0.n18413_cascade_\ : std_logic;
signal \c0.data_in_frame_26_3\ : std_logic;
signal n19127 : std_logic;
signal data_in_frame_22_5 : std_logic;
signal \c0.n9_adj_3069\ : std_logic;
signal \c0.n20451\ : std_logic;
signal \c0.n8_adj_3070\ : std_logic;
signal \c0.n19315\ : std_logic;
signal \c0.n26_adj_3550\ : std_logic;
signal \c0.n27_adj_3551\ : std_logic;
signal \c0.n25_adj_3553\ : std_logic;
signal \c0.n49_adj_3358\ : std_logic;
signal \c0.n17832\ : std_logic;
signal \c0.n40_adj_3271\ : std_logic;
signal rx_data_6 : std_logic;
signal rx_data_2 : std_logic;
signal \c0.n19474\ : std_logic;
signal \c0.data_in_frame_17_2\ : std_logic;
signal \c0.data_in_frame_17_3\ : std_logic;
signal \c0.n14_adj_3436\ : std_logic;
signal \c0.data_in_frame_20_4\ : std_logic;
signal \c0.n19274\ : std_logic;
signal \c0.data_in_frame_20_3\ : std_logic;
signal \c0.n54_adj_3388\ : std_logic;
signal \c0.n32_adj_3310\ : std_logic;
signal \c0.n43_adj_3131\ : std_logic;
signal rx_data_5 : std_logic;
signal \c0.data_in_frame_20_2\ : std_logic;
signal \c0.n20840\ : std_logic;
signal \c0.n22_adj_3322\ : std_logic;
signal \c0.n22_adj_3322_cascade_\ : std_logic;
signal \c0.n36_adj_3090\ : std_logic;
signal \c0.data_in_frame_21_2\ : std_logic;
signal \c0.n29_adj_3383\ : std_logic;
signal \c0.n20917\ : std_logic;
signal \c0.data_in_frame_20_0\ : std_logic;
signal \c0.n4_adj_3435\ : std_logic;
signal \c0.n6_adj_3091\ : std_logic;
signal \c0.n18375\ : std_logic;
signal \c0.n6_adj_3091_cascade_\ : std_logic;
signal \c0.n17900\ : std_logic;
signal \c0.data_in_frame_21_3\ : std_logic;
signal \c0.data_in_frame_21_5\ : std_logic;
signal \c0.n19321\ : std_logic;
signal \c0.n12037\ : std_logic;
signal data_in_frame_19_7 : std_logic;
signal rx_data_3 : std_logic;
signal n19128 : std_logic;
signal data_in_frame_19_3 : std_logic;
signal \c0.n19162\ : std_logic;
signal data_in_frame_22_1 : std_logic;
signal \c0.n20332\ : std_logic;
signal data_in_frame_24_1 : std_logic;
signal data_in_frame_24_3 : std_logic;
signal \c0.n20332_cascade_\ : std_logic;
signal \c0.n18413\ : std_logic;
signal \c0.n36\ : std_logic;
signal \c0.n20642\ : std_logic;
signal \c0.n18525\ : std_logic;
signal data_in_frame_24_2 : std_logic;
signal \c0.n18498\ : std_logic;
signal \c0.n10_adj_3410\ : std_logic;
signal \c0.data_in_frame_20_7\ : std_logic;
signal \c0.data_in_frame_20_6\ : std_logic;
signal \c0.n20576\ : std_logic;
signal \c0.n12_adj_3439\ : std_logic;
signal data_in_frame_22_0 : std_logic;
signal \c0.n18415\ : std_logic;
signal \c0.n4_adj_3067_cascade_\ : std_logic;
signal \c0.n6009\ : std_logic;
signal \c0.n19369\ : std_logic;
signal data_in_frame_19_4 : std_logic;
signal \c0.n11669\ : std_logic;
signal rx_data_4 : std_logic;
signal \c0.data_in_frame_21_6\ : std_logic;
signal \c0.data_in_frame_20_5\ : std_logic;
signal \c0.data_in_frame_21_4\ : std_logic;
signal \c0.n11939_cascade_\ : std_logic;
signal data_in_frame_19_6 : std_logic;
signal \c0.n13_adj_3485\ : std_logic;
signal rx_data_7 : std_logic;
signal \c0.data_in_frame_21_7\ : std_logic;
signal \c0.n19107\ : std_logic;
signal \c0.n12_adj_3361\ : std_logic;
signal rx_data_1 : std_logic;
signal \c0.data_in_frame_21_1\ : std_logic;
signal \CLK_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \LED_wire\ : std_logic;
signal \PIN_12_wire\ : std_logic;
signal \PIN_13_wire\ : std_logic;
signal \PIN_1_wire\ : std_logic;
signal \PIN_22_wire\ : std_logic;
signal \PIN_23_wire\ : std_logic;
signal \PIN_24_wire\ : std_logic;
signal \PIN_2_wire\ : std_logic;
signal \PIN_3_wire\ : std_logic;
signal \PIN_7_wire\ : std_logic;
signal \PIN_8_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    LED <= \LED_wire\;
    \PIN_12_wire\ <= PIN_12;
    \PIN_13_wire\ <= PIN_13;
    PIN_1 <= \PIN_1_wire\;
    PIN_22 <= \PIN_22_wire\;
    PIN_23 <= \PIN_23_wire\;
    PIN_24 <= \PIN_24_wire\;
    PIN_2 <= \PIN_2_wire\;
    PIN_3 <= \PIN_3_wire\;
    \PIN_7_wire\ <= PIN_7;
    \PIN_8_wire\ <= PIN_8;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__73031\,
            DIN => \N__73030\,
            DOUT => \N__73029\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__73031\,
            PADOUT => \N__73030\,
            PADIN => \N__73029\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__24736\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_12_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__73022\,
            DIN => \N__73021\,
            DOUT => \N__73020\,
            PACKAGEPIN => \PIN_12_wire\
        );

    \PIN_12_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__73022\,
            PADOUT => \N__73021\,
            PADIN => \N__73020\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_12_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_13_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__73013\,
            DIN => \N__73012\,
            DOUT => \N__73011\,
            PACKAGEPIN => \PIN_13_wire\
        );

    \PIN_13_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__73013\,
            PADOUT => \N__73012\,
            PADIN => \N__73011\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_13_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__73004\,
            DIN => \N__73003\,
            DOUT => \N__73002\,
            PACKAGEPIN => \PIN_1_wire\
        );

    \PIN_1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__73004\,
            PADOUT => \N__73003\,
            PADIN => \N__73002\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_22_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__72995\,
            DIN => \N__72994\,
            DOUT => \N__72993\,
            PACKAGEPIN => \PIN_22_wire\
        );

    \PIN_22_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__72995\,
            PADOUT => \N__72994\,
            PADIN => \N__72993\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_23_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__72986\,
            DIN => \N__72985\,
            DOUT => \N__72984\,
            PACKAGEPIN => \PIN_23_wire\
        );

    \PIN_23_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__72986\,
            PADOUT => \N__72985\,
            PADIN => \N__72984\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_24_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__72977\,
            DIN => \N__72976\,
            DOUT => \N__72975\,
            PACKAGEPIN => \PIN_24_wire\
        );

    \PIN_24_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__72977\,
            PADOUT => \N__72976\,
            PADIN => \N__72975\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__72968\,
            DIN => \N__72967\,
            DOUT => \N__72966\,
            PACKAGEPIN => \PIN_2_wire\
        );

    \PIN_2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__72968\,
            PADOUT => \N__72967\,
            PADIN => \N__72966\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__72959\,
            DIN => \N__72958\,
            DOUT => \N__72957\,
            PACKAGEPIN => \PIN_3_wire\
        );

    \PIN_3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__72959\,
            PADOUT => \N__72958\,
            PADIN => \N__72957\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_7_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__72950\,
            DIN => \N__72949\,
            DOUT => \N__72948\,
            PACKAGEPIN => \PIN_7_wire\
        );

    \PIN_7_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__72950\,
            PADOUT => \N__72949\,
            PADIN => \N__72948\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_7_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_8_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__72941\,
            DIN => \N__72940\,
            DOUT => \N__72939\,
            PACKAGEPIN => \PIN_8_wire\
        );

    \PIN_8_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__72941\,
            PADOUT => \N__72940\,
            PADIN => \N__72939\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_8_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__72932\,
            DIN => \N__72931\,
            DOUT => \N__72930\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__72932\,
            PADOUT => \N__72931\,
            PADIN => \N__72930\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall1_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__72923\,
            DIN => \N__72922\,
            DOUT => \N__72921\,
            PACKAGEPIN => PIN_4
        );

    \hall1_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__72923\,
            PADOUT => \N__72922\,
            PADIN => \N__72921\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall2_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__72914\,
            DIN => \N__72913\,
            DOUT => \N__72912\,
            PACKAGEPIN => PIN_5
        );

    \hall2_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__72914\,
            PADOUT => \N__72913\,
            PADIN => \N__72912\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall3_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__72905\,
            DIN => \N__72904\,
            DOUT => \N__72903\,
            PACKAGEPIN => PIN_6
        );

    \hall3_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__72905\,
            PADOUT => \N__72904\,
            PADIN => \N__72903\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rx_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__72896\,
            DIN => \N__72895\,
            DOUT => \N__72894\,
            PACKAGEPIN => PIN_11
        );

    \rx_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__72896\,
            PADOUT => \N__72895\,
            PADIN => \N__72894\,
            CLOCKENABLE => 'H',
            DIN0 => \LED_c\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \tx_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__72887\,
            DIN => \N__72886\,
            DOUT => \N__72885\,
            PACKAGEPIN => PIN_10
        );

    \tx_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__72887\,
            PADOUT => \N__72886\,
            PADIN => \N__72885\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__34183\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__24745\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__72878\,
            DIN => \N__72877\,
            DOUT => \N__72876\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__72878\,
            PADOUT => \N__72877\,
            PADIN => \N__72876\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__18132\ : InMux
    port map (
            O => \N__72859\,
            I => \N__72855\
        );

    \I__18131\ : InMux
    port map (
            O => \N__72858\,
            I => \N__72852\
        );

    \I__18130\ : LocalMux
    port map (
            O => \N__72855\,
            I => \N__72848\
        );

    \I__18129\ : LocalMux
    port map (
            O => \N__72852\,
            I => \N__72845\
        );

    \I__18128\ : CascadeMux
    port map (
            O => \N__72851\,
            I => \N__72841\
        );

    \I__18127\ : Span4Mux_h
    port map (
            O => \N__72848\,
            I => \N__72838\
        );

    \I__18126\ : Span4Mux_v
    port map (
            O => \N__72845\,
            I => \N__72835\
        );

    \I__18125\ : CascadeMux
    port map (
            O => \N__72844\,
            I => \N__72828\
        );

    \I__18124\ : InMux
    port map (
            O => \N__72841\,
            I => \N__72824\
        );

    \I__18123\ : Span4Mux_v
    port map (
            O => \N__72838\,
            I => \N__72819\
        );

    \I__18122\ : Span4Mux_h
    port map (
            O => \N__72835\,
            I => \N__72819\
        );

    \I__18121\ : InMux
    port map (
            O => \N__72834\,
            I => \N__72812\
        );

    \I__18120\ : InMux
    port map (
            O => \N__72833\,
            I => \N__72812\
        );

    \I__18119\ : InMux
    port map (
            O => \N__72832\,
            I => \N__72812\
        );

    \I__18118\ : InMux
    port map (
            O => \N__72831\,
            I => \N__72809\
        );

    \I__18117\ : InMux
    port map (
            O => \N__72828\,
            I => \N__72806\
        );

    \I__18116\ : InMux
    port map (
            O => \N__72827\,
            I => \N__72803\
        );

    \I__18115\ : LocalMux
    port map (
            O => \N__72824\,
            I => \N__72800\
        );

    \I__18114\ : Sp12to4
    port map (
            O => \N__72819\,
            I => \N__72795\
        );

    \I__18113\ : LocalMux
    port map (
            O => \N__72812\,
            I => \N__72795\
        );

    \I__18112\ : LocalMux
    port map (
            O => \N__72809\,
            I => \N__72790\
        );

    \I__18111\ : LocalMux
    port map (
            O => \N__72806\,
            I => \N__72790\
        );

    \I__18110\ : LocalMux
    port map (
            O => \N__72803\,
            I => data_in_frame_19_4
        );

    \I__18109\ : Odrv4
    port map (
            O => \N__72800\,
            I => data_in_frame_19_4
        );

    \I__18108\ : Odrv12
    port map (
            O => \N__72795\,
            I => data_in_frame_19_4
        );

    \I__18107\ : Odrv4
    port map (
            O => \N__72790\,
            I => data_in_frame_19_4
        );

    \I__18106\ : InMux
    port map (
            O => \N__72781\,
            I => \N__72778\
        );

    \I__18105\ : LocalMux
    port map (
            O => \N__72778\,
            I => \c0.n11669\
        );

    \I__18104\ : InMux
    port map (
            O => \N__72775\,
            I => \N__72771\
        );

    \I__18103\ : InMux
    port map (
            O => \N__72774\,
            I => \N__72768\
        );

    \I__18102\ : LocalMux
    port map (
            O => \N__72771\,
            I => \N__72761\
        );

    \I__18101\ : LocalMux
    port map (
            O => \N__72768\,
            I => \N__72761\
        );

    \I__18100\ : InMux
    port map (
            O => \N__72767\,
            I => \N__72756\
        );

    \I__18099\ : InMux
    port map (
            O => \N__72766\,
            I => \N__72756\
        );

    \I__18098\ : Span4Mux_h
    port map (
            O => \N__72761\,
            I => \N__72749\
        );

    \I__18097\ : LocalMux
    port map (
            O => \N__72756\,
            I => \N__72749\
        );

    \I__18096\ : CascadeMux
    port map (
            O => \N__72755\,
            I => \N__72745\
        );

    \I__18095\ : InMux
    port map (
            O => \N__72754\,
            I => \N__72741\
        );

    \I__18094\ : Span4Mux_v
    port map (
            O => \N__72749\,
            I => \N__72734\
        );

    \I__18093\ : InMux
    port map (
            O => \N__72748\,
            I => \N__72730\
        );

    \I__18092\ : InMux
    port map (
            O => \N__72745\,
            I => \N__72726\
        );

    \I__18091\ : InMux
    port map (
            O => \N__72744\,
            I => \N__72723\
        );

    \I__18090\ : LocalMux
    port map (
            O => \N__72741\,
            I => \N__72720\
        );

    \I__18089\ : InMux
    port map (
            O => \N__72740\,
            I => \N__72717\
        );

    \I__18088\ : InMux
    port map (
            O => \N__72739\,
            I => \N__72712\
        );

    \I__18087\ : InMux
    port map (
            O => \N__72738\,
            I => \N__72712\
        );

    \I__18086\ : InMux
    port map (
            O => \N__72737\,
            I => \N__72707\
        );

    \I__18085\ : Span4Mux_h
    port map (
            O => \N__72734\,
            I => \N__72704\
        );

    \I__18084\ : InMux
    port map (
            O => \N__72733\,
            I => \N__72701\
        );

    \I__18083\ : LocalMux
    port map (
            O => \N__72730\,
            I => \N__72694\
        );

    \I__18082\ : InMux
    port map (
            O => \N__72729\,
            I => \N__72691\
        );

    \I__18081\ : LocalMux
    port map (
            O => \N__72726\,
            I => \N__72686\
        );

    \I__18080\ : LocalMux
    port map (
            O => \N__72723\,
            I => \N__72686\
        );

    \I__18079\ : Span4Mux_v
    port map (
            O => \N__72720\,
            I => \N__72681\
        );

    \I__18078\ : LocalMux
    port map (
            O => \N__72717\,
            I => \N__72681\
        );

    \I__18077\ : LocalMux
    port map (
            O => \N__72712\,
            I => \N__72678\
        );

    \I__18076\ : InMux
    port map (
            O => \N__72711\,
            I => \N__72674\
        );

    \I__18075\ : InMux
    port map (
            O => \N__72710\,
            I => \N__72669\
        );

    \I__18074\ : LocalMux
    port map (
            O => \N__72707\,
            I => \N__72666\
        );

    \I__18073\ : Span4Mux_h
    port map (
            O => \N__72704\,
            I => \N__72661\
        );

    \I__18072\ : LocalMux
    port map (
            O => \N__72701\,
            I => \N__72661\
        );

    \I__18071\ : InMux
    port map (
            O => \N__72700\,
            I => \N__72656\
        );

    \I__18070\ : InMux
    port map (
            O => \N__72699\,
            I => \N__72653\
        );

    \I__18069\ : InMux
    port map (
            O => \N__72698\,
            I => \N__72650\
        );

    \I__18068\ : InMux
    port map (
            O => \N__72697\,
            I => \N__72646\
        );

    \I__18067\ : Span4Mux_v
    port map (
            O => \N__72694\,
            I => \N__72641\
        );

    \I__18066\ : LocalMux
    port map (
            O => \N__72691\,
            I => \N__72641\
        );

    \I__18065\ : Span4Mux_v
    port map (
            O => \N__72686\,
            I => \N__72636\
        );

    \I__18064\ : Span4Mux_h
    port map (
            O => \N__72681\,
            I => \N__72636\
        );

    \I__18063\ : Span4Mux_h
    port map (
            O => \N__72678\,
            I => \N__72633\
        );

    \I__18062\ : InMux
    port map (
            O => \N__72677\,
            I => \N__72630\
        );

    \I__18061\ : LocalMux
    port map (
            O => \N__72674\,
            I => \N__72627\
        );

    \I__18060\ : InMux
    port map (
            O => \N__72673\,
            I => \N__72622\
        );

    \I__18059\ : InMux
    port map (
            O => \N__72672\,
            I => \N__72622\
        );

    \I__18058\ : LocalMux
    port map (
            O => \N__72669\,
            I => \N__72615\
        );

    \I__18057\ : Span4Mux_v
    port map (
            O => \N__72666\,
            I => \N__72615\
        );

    \I__18056\ : Span4Mux_v
    port map (
            O => \N__72661\,
            I => \N__72615\
        );

    \I__18055\ : InMux
    port map (
            O => \N__72660\,
            I => \N__72607\
        );

    \I__18054\ : InMux
    port map (
            O => \N__72659\,
            I => \N__72604\
        );

    \I__18053\ : LocalMux
    port map (
            O => \N__72656\,
            I => \N__72601\
        );

    \I__18052\ : LocalMux
    port map (
            O => \N__72653\,
            I => \N__72598\
        );

    \I__18051\ : LocalMux
    port map (
            O => \N__72650\,
            I => \N__72595\
        );

    \I__18050\ : InMux
    port map (
            O => \N__72649\,
            I => \N__72592\
        );

    \I__18049\ : LocalMux
    port map (
            O => \N__72646\,
            I => \N__72589\
        );

    \I__18048\ : Span4Mux_v
    port map (
            O => \N__72641\,
            I => \N__72584\
        );

    \I__18047\ : Span4Mux_h
    port map (
            O => \N__72636\,
            I => \N__72584\
        );

    \I__18046\ : Span4Mux_h
    port map (
            O => \N__72633\,
            I => \N__72575\
        );

    \I__18045\ : LocalMux
    port map (
            O => \N__72630\,
            I => \N__72575\
        );

    \I__18044\ : Span4Mux_h
    port map (
            O => \N__72627\,
            I => \N__72575\
        );

    \I__18043\ : LocalMux
    port map (
            O => \N__72622\,
            I => \N__72575\
        );

    \I__18042\ : Sp12to4
    port map (
            O => \N__72615\,
            I => \N__72572\
        );

    \I__18041\ : InMux
    port map (
            O => \N__72614\,
            I => \N__72569\
        );

    \I__18040\ : InMux
    port map (
            O => \N__72613\,
            I => \N__72566\
        );

    \I__18039\ : InMux
    port map (
            O => \N__72612\,
            I => \N__72563\
        );

    \I__18038\ : InMux
    port map (
            O => \N__72611\,
            I => \N__72558\
        );

    \I__18037\ : InMux
    port map (
            O => \N__72610\,
            I => \N__72558\
        );

    \I__18036\ : LocalMux
    port map (
            O => \N__72607\,
            I => \N__72549\
        );

    \I__18035\ : LocalMux
    port map (
            O => \N__72604\,
            I => \N__72549\
        );

    \I__18034\ : Span4Mux_v
    port map (
            O => \N__72601\,
            I => \N__72549\
        );

    \I__18033\ : Span4Mux_v
    port map (
            O => \N__72598\,
            I => \N__72549\
        );

    \I__18032\ : Span4Mux_h
    port map (
            O => \N__72595\,
            I => \N__72546\
        );

    \I__18031\ : LocalMux
    port map (
            O => \N__72592\,
            I => \N__72541\
        );

    \I__18030\ : Span4Mux_v
    port map (
            O => \N__72589\,
            I => \N__72541\
        );

    \I__18029\ : Span4Mux_v
    port map (
            O => \N__72584\,
            I => \N__72538\
        );

    \I__18028\ : Span4Mux_v
    port map (
            O => \N__72575\,
            I => \N__72535\
        );

    \I__18027\ : Span12Mux_h
    port map (
            O => \N__72572\,
            I => \N__72532\
        );

    \I__18026\ : LocalMux
    port map (
            O => \N__72569\,
            I => \N__72528\
        );

    \I__18025\ : LocalMux
    port map (
            O => \N__72566\,
            I => \N__72525\
        );

    \I__18024\ : LocalMux
    port map (
            O => \N__72563\,
            I => \N__72522\
        );

    \I__18023\ : LocalMux
    port map (
            O => \N__72558\,
            I => \N__72517\
        );

    \I__18022\ : Span4Mux_h
    port map (
            O => \N__72549\,
            I => \N__72517\
        );

    \I__18021\ : Span4Mux_h
    port map (
            O => \N__72546\,
            I => \N__72510\
        );

    \I__18020\ : Span4Mux_h
    port map (
            O => \N__72541\,
            I => \N__72510\
        );

    \I__18019\ : Span4Mux_v
    port map (
            O => \N__72538\,
            I => \N__72510\
        );

    \I__18018\ : Sp12to4
    port map (
            O => \N__72535\,
            I => \N__72505\
        );

    \I__18017\ : Span12Mux_v
    port map (
            O => \N__72532\,
            I => \N__72505\
        );

    \I__18016\ : InMux
    port map (
            O => \N__72531\,
            I => \N__72502\
        );

    \I__18015\ : Span4Mux_h
    port map (
            O => \N__72528\,
            I => \N__72499\
        );

    \I__18014\ : Span4Mux_v
    port map (
            O => \N__72525\,
            I => \N__72496\
        );

    \I__18013\ : Span4Mux_h
    port map (
            O => \N__72522\,
            I => \N__72491\
        );

    \I__18012\ : Span4Mux_v
    port map (
            O => \N__72517\,
            I => \N__72491\
        );

    \I__18011\ : Sp12to4
    port map (
            O => \N__72510\,
            I => \N__72486\
        );

    \I__18010\ : Span12Mux_h
    port map (
            O => \N__72505\,
            I => \N__72486\
        );

    \I__18009\ : LocalMux
    port map (
            O => \N__72502\,
            I => rx_data_4
        );

    \I__18008\ : Odrv4
    port map (
            O => \N__72499\,
            I => rx_data_4
        );

    \I__18007\ : Odrv4
    port map (
            O => \N__72496\,
            I => rx_data_4
        );

    \I__18006\ : Odrv4
    port map (
            O => \N__72491\,
            I => rx_data_4
        );

    \I__18005\ : Odrv12
    port map (
            O => \N__72486\,
            I => rx_data_4
        );

    \I__18004\ : InMux
    port map (
            O => \N__72475\,
            I => \N__72468\
        );

    \I__18003\ : InMux
    port map (
            O => \N__72474\,
            I => \N__72468\
        );

    \I__18002\ : CascadeMux
    port map (
            O => \N__72473\,
            I => \N__72463\
        );

    \I__18001\ : LocalMux
    port map (
            O => \N__72468\,
            I => \N__72460\
        );

    \I__18000\ : InMux
    port map (
            O => \N__72467\,
            I => \N__72455\
        );

    \I__17999\ : InMux
    port map (
            O => \N__72466\,
            I => \N__72455\
        );

    \I__17998\ : InMux
    port map (
            O => \N__72463\,
            I => \N__72452\
        );

    \I__17997\ : Span4Mux_v
    port map (
            O => \N__72460\,
            I => \N__72449\
        );

    \I__17996\ : LocalMux
    port map (
            O => \N__72455\,
            I => \N__72446\
        );

    \I__17995\ : LocalMux
    port map (
            O => \N__72452\,
            I => \c0.data_in_frame_21_6\
        );

    \I__17994\ : Odrv4
    port map (
            O => \N__72449\,
            I => \c0.data_in_frame_21_6\
        );

    \I__17993\ : Odrv4
    port map (
            O => \N__72446\,
            I => \c0.data_in_frame_21_6\
        );

    \I__17992\ : InMux
    port map (
            O => \N__72439\,
            I => \N__72434\
        );

    \I__17991\ : InMux
    port map (
            O => \N__72438\,
            I => \N__72429\
        );

    \I__17990\ : InMux
    port map (
            O => \N__72437\,
            I => \N__72429\
        );

    \I__17989\ : LocalMux
    port map (
            O => \N__72434\,
            I => \N__72426\
        );

    \I__17988\ : LocalMux
    port map (
            O => \N__72429\,
            I => \N__72421\
        );

    \I__17987\ : Span4Mux_v
    port map (
            O => \N__72426\,
            I => \N__72418\
        );

    \I__17986\ : InMux
    port map (
            O => \N__72425\,
            I => \N__72415\
        );

    \I__17985\ : InMux
    port map (
            O => \N__72424\,
            I => \N__72412\
        );

    \I__17984\ : Span12Mux_s11_v
    port map (
            O => \N__72421\,
            I => \N__72409\
        );

    \I__17983\ : Span4Mux_v
    port map (
            O => \N__72418\,
            I => \N__72404\
        );

    \I__17982\ : LocalMux
    port map (
            O => \N__72415\,
            I => \N__72404\
        );

    \I__17981\ : LocalMux
    port map (
            O => \N__72412\,
            I => \c0.data_in_frame_20_5\
        );

    \I__17980\ : Odrv12
    port map (
            O => \N__72409\,
            I => \c0.data_in_frame_20_5\
        );

    \I__17979\ : Odrv4
    port map (
            O => \N__72404\,
            I => \c0.data_in_frame_20_5\
        );

    \I__17978\ : CascadeMux
    port map (
            O => \N__72397\,
            I => \N__72394\
        );

    \I__17977\ : InMux
    port map (
            O => \N__72394\,
            I => \N__72389\
        );

    \I__17976\ : CascadeMux
    port map (
            O => \N__72393\,
            I => \N__72386\
        );

    \I__17975\ : InMux
    port map (
            O => \N__72392\,
            I => \N__72382\
        );

    \I__17974\ : LocalMux
    port map (
            O => \N__72389\,
            I => \N__72379\
        );

    \I__17973\ : InMux
    port map (
            O => \N__72386\,
            I => \N__72376\
        );

    \I__17972\ : InMux
    port map (
            O => \N__72385\,
            I => \N__72373\
        );

    \I__17971\ : LocalMux
    port map (
            O => \N__72382\,
            I => \N__72370\
        );

    \I__17970\ : Span4Mux_v
    port map (
            O => \N__72379\,
            I => \N__72366\
        );

    \I__17969\ : LocalMux
    port map (
            O => \N__72376\,
            I => \N__72359\
        );

    \I__17968\ : LocalMux
    port map (
            O => \N__72373\,
            I => \N__72359\
        );

    \I__17967\ : Span4Mux_v
    port map (
            O => \N__72370\,
            I => \N__72359\
        );

    \I__17966\ : InMux
    port map (
            O => \N__72369\,
            I => \N__72356\
        );

    \I__17965\ : Odrv4
    port map (
            O => \N__72366\,
            I => \c0.data_in_frame_21_4\
        );

    \I__17964\ : Odrv4
    port map (
            O => \N__72359\,
            I => \c0.data_in_frame_21_4\
        );

    \I__17963\ : LocalMux
    port map (
            O => \N__72356\,
            I => \c0.data_in_frame_21_4\
        );

    \I__17962\ : CascadeMux
    port map (
            O => \N__72349\,
            I => \c0.n11939_cascade_\
        );

    \I__17961\ : InMux
    port map (
            O => \N__72346\,
            I => \N__72343\
        );

    \I__17960\ : LocalMux
    port map (
            O => \N__72343\,
            I => \N__72339\
        );

    \I__17959\ : CascadeMux
    port map (
            O => \N__72342\,
            I => \N__72332\
        );

    \I__17958\ : Span4Mux_v
    port map (
            O => \N__72339\,
            I => \N__72329\
        );

    \I__17957\ : InMux
    port map (
            O => \N__72338\,
            I => \N__72324\
        );

    \I__17956\ : InMux
    port map (
            O => \N__72337\,
            I => \N__72324\
        );

    \I__17955\ : InMux
    port map (
            O => \N__72336\,
            I => \N__72319\
        );

    \I__17954\ : InMux
    port map (
            O => \N__72335\,
            I => \N__72319\
        );

    \I__17953\ : InMux
    port map (
            O => \N__72332\,
            I => \N__72316\
        );

    \I__17952\ : Sp12to4
    port map (
            O => \N__72329\,
            I => \N__72309\
        );

    \I__17951\ : LocalMux
    port map (
            O => \N__72324\,
            I => \N__72309\
        );

    \I__17950\ : LocalMux
    port map (
            O => \N__72319\,
            I => \N__72309\
        );

    \I__17949\ : LocalMux
    port map (
            O => \N__72316\,
            I => data_in_frame_19_6
        );

    \I__17948\ : Odrv12
    port map (
            O => \N__72309\,
            I => data_in_frame_19_6
        );

    \I__17947\ : InMux
    port map (
            O => \N__72304\,
            I => \N__72301\
        );

    \I__17946\ : LocalMux
    port map (
            O => \N__72301\,
            I => \N__72298\
        );

    \I__17945\ : Odrv4
    port map (
            O => \N__72298\,
            I => \c0.n13_adj_3485\
        );

    \I__17944\ : InMux
    port map (
            O => \N__72295\,
            I => \N__72288\
        );

    \I__17943\ : InMux
    port map (
            O => \N__72294\,
            I => \N__72280\
        );

    \I__17942\ : InMux
    port map (
            O => \N__72293\,
            I => \N__72277\
        );

    \I__17941\ : InMux
    port map (
            O => \N__72292\,
            I => \N__72274\
        );

    \I__17940\ : InMux
    port map (
            O => \N__72291\,
            I => \N__72271\
        );

    \I__17939\ : LocalMux
    port map (
            O => \N__72288\,
            I => \N__72267\
        );

    \I__17938\ : InMux
    port map (
            O => \N__72287\,
            I => \N__72262\
        );

    \I__17937\ : InMux
    port map (
            O => \N__72286\,
            I => \N__72262\
        );

    \I__17936\ : InMux
    port map (
            O => \N__72285\,
            I => \N__72257\
        );

    \I__17935\ : InMux
    port map (
            O => \N__72284\,
            I => \N__72251\
        );

    \I__17934\ : InMux
    port map (
            O => \N__72283\,
            I => \N__72248\
        );

    \I__17933\ : LocalMux
    port map (
            O => \N__72280\,
            I => \N__72243\
        );

    \I__17932\ : LocalMux
    port map (
            O => \N__72277\,
            I => \N__72243\
        );

    \I__17931\ : LocalMux
    port map (
            O => \N__72274\,
            I => \N__72238\
        );

    \I__17930\ : LocalMux
    port map (
            O => \N__72271\,
            I => \N__72235\
        );

    \I__17929\ : CascadeMux
    port map (
            O => \N__72270\,
            I => \N__72232\
        );

    \I__17928\ : Span4Mux_h
    port map (
            O => \N__72267\,
            I => \N__72228\
        );

    \I__17927\ : LocalMux
    port map (
            O => \N__72262\,
            I => \N__72225\
        );

    \I__17926\ : InMux
    port map (
            O => \N__72261\,
            I => \N__72222\
        );

    \I__17925\ : InMux
    port map (
            O => \N__72260\,
            I => \N__72218\
        );

    \I__17924\ : LocalMux
    port map (
            O => \N__72257\,
            I => \N__72214\
        );

    \I__17923\ : InMux
    port map (
            O => \N__72256\,
            I => \N__72211\
        );

    \I__17922\ : InMux
    port map (
            O => \N__72255\,
            I => \N__72208\
        );

    \I__17921\ : InMux
    port map (
            O => \N__72254\,
            I => \N__72202\
        );

    \I__17920\ : LocalMux
    port map (
            O => \N__72251\,
            I => \N__72196\
        );

    \I__17919\ : LocalMux
    port map (
            O => \N__72248\,
            I => \N__72193\
        );

    \I__17918\ : Span4Mux_h
    port map (
            O => \N__72243\,
            I => \N__72190\
        );

    \I__17917\ : InMux
    port map (
            O => \N__72242\,
            I => \N__72187\
        );

    \I__17916\ : InMux
    port map (
            O => \N__72241\,
            I => \N__72184\
        );

    \I__17915\ : Span4Mux_v
    port map (
            O => \N__72238\,
            I => \N__72181\
        );

    \I__17914\ : Span4Mux_v
    port map (
            O => \N__72235\,
            I => \N__72178\
        );

    \I__17913\ : InMux
    port map (
            O => \N__72232\,
            I => \N__72175\
        );

    \I__17912\ : InMux
    port map (
            O => \N__72231\,
            I => \N__72172\
        );

    \I__17911\ : Span4Mux_v
    port map (
            O => \N__72228\,
            I => \N__72165\
        );

    \I__17910\ : Span4Mux_v
    port map (
            O => \N__72225\,
            I => \N__72165\
        );

    \I__17909\ : LocalMux
    port map (
            O => \N__72222\,
            I => \N__72165\
        );

    \I__17908\ : InMux
    port map (
            O => \N__72221\,
            I => \N__72162\
        );

    \I__17907\ : LocalMux
    port map (
            O => \N__72218\,
            I => \N__72159\
        );

    \I__17906\ : InMux
    port map (
            O => \N__72217\,
            I => \N__72156\
        );

    \I__17905\ : Span4Mux_v
    port map (
            O => \N__72214\,
            I => \N__72153\
        );

    \I__17904\ : LocalMux
    port map (
            O => \N__72211\,
            I => \N__72150\
        );

    \I__17903\ : LocalMux
    port map (
            O => \N__72208\,
            I => \N__72146\
        );

    \I__17902\ : InMux
    port map (
            O => \N__72207\,
            I => \N__72141\
        );

    \I__17901\ : InMux
    port map (
            O => \N__72206\,
            I => \N__72136\
        );

    \I__17900\ : InMux
    port map (
            O => \N__72205\,
            I => \N__72136\
        );

    \I__17899\ : LocalMux
    port map (
            O => \N__72202\,
            I => \N__72133\
        );

    \I__17898\ : CascadeMux
    port map (
            O => \N__72201\,
            I => \N__72129\
        );

    \I__17897\ : InMux
    port map (
            O => \N__72200\,
            I => \N__72125\
        );

    \I__17896\ : InMux
    port map (
            O => \N__72199\,
            I => \N__72122\
        );

    \I__17895\ : Span4Mux_v
    port map (
            O => \N__72196\,
            I => \N__72117\
        );

    \I__17894\ : Span4Mux_v
    port map (
            O => \N__72193\,
            I => \N__72117\
        );

    \I__17893\ : Span4Mux_h
    port map (
            O => \N__72190\,
            I => \N__72114\
        );

    \I__17892\ : LocalMux
    port map (
            O => \N__72187\,
            I => \N__72105\
        );

    \I__17891\ : LocalMux
    port map (
            O => \N__72184\,
            I => \N__72105\
        );

    \I__17890\ : Sp12to4
    port map (
            O => \N__72181\,
            I => \N__72105\
        );

    \I__17889\ : Sp12to4
    port map (
            O => \N__72178\,
            I => \N__72105\
        );

    \I__17888\ : LocalMux
    port map (
            O => \N__72175\,
            I => \N__72100\
        );

    \I__17887\ : LocalMux
    port map (
            O => \N__72172\,
            I => \N__72100\
        );

    \I__17886\ : Span4Mux_h
    port map (
            O => \N__72165\,
            I => \N__72097\
        );

    \I__17885\ : LocalMux
    port map (
            O => \N__72162\,
            I => \N__72092\
        );

    \I__17884\ : Span4Mux_h
    port map (
            O => \N__72159\,
            I => \N__72092\
        );

    \I__17883\ : LocalMux
    port map (
            O => \N__72156\,
            I => \N__72085\
        );

    \I__17882\ : Span4Mux_h
    port map (
            O => \N__72153\,
            I => \N__72085\
        );

    \I__17881\ : Span4Mux_h
    port map (
            O => \N__72150\,
            I => \N__72085\
        );

    \I__17880\ : InMux
    port map (
            O => \N__72149\,
            I => \N__72082\
        );

    \I__17879\ : Span4Mux_h
    port map (
            O => \N__72146\,
            I => \N__72079\
        );

    \I__17878\ : InMux
    port map (
            O => \N__72145\,
            I => \N__72074\
        );

    \I__17877\ : InMux
    port map (
            O => \N__72144\,
            I => \N__72074\
        );

    \I__17876\ : LocalMux
    port map (
            O => \N__72141\,
            I => \N__72071\
        );

    \I__17875\ : LocalMux
    port map (
            O => \N__72136\,
            I => \N__72066\
        );

    \I__17874\ : Span4Mux_v
    port map (
            O => \N__72133\,
            I => \N__72066\
        );

    \I__17873\ : InMux
    port map (
            O => \N__72132\,
            I => \N__72059\
        );

    \I__17872\ : InMux
    port map (
            O => \N__72129\,
            I => \N__72059\
        );

    \I__17871\ : InMux
    port map (
            O => \N__72128\,
            I => \N__72059\
        );

    \I__17870\ : LocalMux
    port map (
            O => \N__72125\,
            I => \N__72054\
        );

    \I__17869\ : LocalMux
    port map (
            O => \N__72122\,
            I => \N__72054\
        );

    \I__17868\ : Span4Mux_v
    port map (
            O => \N__72117\,
            I => \N__72051\
        );

    \I__17867\ : Sp12to4
    port map (
            O => \N__72114\,
            I => \N__72046\
        );

    \I__17866\ : Span12Mux_h
    port map (
            O => \N__72105\,
            I => \N__72046\
        );

    \I__17865\ : Span4Mux_v
    port map (
            O => \N__72100\,
            I => \N__72043\
        );

    \I__17864\ : Span4Mux_h
    port map (
            O => \N__72097\,
            I => \N__72036\
        );

    \I__17863\ : Span4Mux_h
    port map (
            O => \N__72092\,
            I => \N__72036\
        );

    \I__17862\ : Span4Mux_v
    port map (
            O => \N__72085\,
            I => \N__72036\
        );

    \I__17861\ : LocalMux
    port map (
            O => \N__72082\,
            I => \N__72031\
        );

    \I__17860\ : Sp12to4
    port map (
            O => \N__72079\,
            I => \N__72031\
        );

    \I__17859\ : LocalMux
    port map (
            O => \N__72074\,
            I => \N__72024\
        );

    \I__17858\ : Span4Mux_h
    port map (
            O => \N__72071\,
            I => \N__72024\
        );

    \I__17857\ : Span4Mux_v
    port map (
            O => \N__72066\,
            I => \N__72024\
        );

    \I__17856\ : LocalMux
    port map (
            O => \N__72059\,
            I => \N__72019\
        );

    \I__17855\ : Span12Mux_s11_v
    port map (
            O => \N__72054\,
            I => \N__72019\
        );

    \I__17854\ : Sp12to4
    port map (
            O => \N__72051\,
            I => \N__72014\
        );

    \I__17853\ : Span12Mux_v
    port map (
            O => \N__72046\,
            I => \N__72014\
        );

    \I__17852\ : Span4Mux_h
    port map (
            O => \N__72043\,
            I => \N__72009\
        );

    \I__17851\ : Span4Mux_v
    port map (
            O => \N__72036\,
            I => \N__72009\
        );

    \I__17850\ : Odrv12
    port map (
            O => \N__72031\,
            I => rx_data_7
        );

    \I__17849\ : Odrv4
    port map (
            O => \N__72024\,
            I => rx_data_7
        );

    \I__17848\ : Odrv12
    port map (
            O => \N__72019\,
            I => rx_data_7
        );

    \I__17847\ : Odrv12
    port map (
            O => \N__72014\,
            I => rx_data_7
        );

    \I__17846\ : Odrv4
    port map (
            O => \N__72009\,
            I => rx_data_7
        );

    \I__17845\ : InMux
    port map (
            O => \N__71998\,
            I => \N__71995\
        );

    \I__17844\ : LocalMux
    port map (
            O => \N__71995\,
            I => \N__71989\
        );

    \I__17843\ : InMux
    port map (
            O => \N__71994\,
            I => \N__71982\
        );

    \I__17842\ : InMux
    port map (
            O => \N__71993\,
            I => \N__71982\
        );

    \I__17841\ : InMux
    port map (
            O => \N__71992\,
            I => \N__71982\
        );

    \I__17840\ : Odrv4
    port map (
            O => \N__71989\,
            I => \c0.data_in_frame_21_7\
        );

    \I__17839\ : LocalMux
    port map (
            O => \N__71982\,
            I => \c0.data_in_frame_21_7\
        );

    \I__17838\ : InMux
    port map (
            O => \N__71977\,
            I => \N__71974\
        );

    \I__17837\ : LocalMux
    port map (
            O => \N__71974\,
            I => \N__71966\
        );

    \I__17836\ : CascadeMux
    port map (
            O => \N__71973\,
            I => \N__71955\
        );

    \I__17835\ : InMux
    port map (
            O => \N__71972\,
            I => \N__71952\
        );

    \I__17834\ : InMux
    port map (
            O => \N__71971\,
            I => \N__71949\
        );

    \I__17833\ : InMux
    port map (
            O => \N__71970\,
            I => \N__71942\
        );

    \I__17832\ : InMux
    port map (
            O => \N__71969\,
            I => \N__71942\
        );

    \I__17831\ : Span4Mux_h
    port map (
            O => \N__71966\,
            I => \N__71938\
        );

    \I__17830\ : InMux
    port map (
            O => \N__71965\,
            I => \N__71935\
        );

    \I__17829\ : InMux
    port map (
            O => \N__71964\,
            I => \N__71929\
        );

    \I__17828\ : InMux
    port map (
            O => \N__71963\,
            I => \N__71922\
        );

    \I__17827\ : InMux
    port map (
            O => \N__71962\,
            I => \N__71922\
        );

    \I__17826\ : InMux
    port map (
            O => \N__71961\,
            I => \N__71922\
        );

    \I__17825\ : InMux
    port map (
            O => \N__71960\,
            I => \N__71917\
        );

    \I__17824\ : InMux
    port map (
            O => \N__71959\,
            I => \N__71917\
        );

    \I__17823\ : InMux
    port map (
            O => \N__71958\,
            I => \N__71912\
        );

    \I__17822\ : InMux
    port map (
            O => \N__71955\,
            I => \N__71912\
        );

    \I__17821\ : LocalMux
    port map (
            O => \N__71952\,
            I => \N__71907\
        );

    \I__17820\ : LocalMux
    port map (
            O => \N__71949\,
            I => \N__71907\
        );

    \I__17819\ : InMux
    port map (
            O => \N__71948\,
            I => \N__71902\
        );

    \I__17818\ : InMux
    port map (
            O => \N__71947\,
            I => \N__71902\
        );

    \I__17817\ : LocalMux
    port map (
            O => \N__71942\,
            I => \N__71899\
        );

    \I__17816\ : InMux
    port map (
            O => \N__71941\,
            I => \N__71895\
        );

    \I__17815\ : Span4Mux_v
    port map (
            O => \N__71938\,
            I => \N__71890\
        );

    \I__17814\ : LocalMux
    port map (
            O => \N__71935\,
            I => \N__71890\
        );

    \I__17813\ : InMux
    port map (
            O => \N__71934\,
            I => \N__71883\
        );

    \I__17812\ : InMux
    port map (
            O => \N__71933\,
            I => \N__71883\
        );

    \I__17811\ : InMux
    port map (
            O => \N__71932\,
            I => \N__71883\
        );

    \I__17810\ : LocalMux
    port map (
            O => \N__71929\,
            I => \N__71876\
        );

    \I__17809\ : LocalMux
    port map (
            O => \N__71922\,
            I => \N__71876\
        );

    \I__17808\ : LocalMux
    port map (
            O => \N__71917\,
            I => \N__71876\
        );

    \I__17807\ : LocalMux
    port map (
            O => \N__71912\,
            I => \N__71871\
        );

    \I__17806\ : Span4Mux_v
    port map (
            O => \N__71907\,
            I => \N__71871\
        );

    \I__17805\ : LocalMux
    port map (
            O => \N__71902\,
            I => \N__71863\
        );

    \I__17804\ : Span4Mux_v
    port map (
            O => \N__71899\,
            I => \N__71863\
        );

    \I__17803\ : CascadeMux
    port map (
            O => \N__71898\,
            I => \N__71860\
        );

    \I__17802\ : LocalMux
    port map (
            O => \N__71895\,
            I => \N__71857\
        );

    \I__17801\ : Span4Mux_h
    port map (
            O => \N__71890\,
            I => \N__71854\
        );

    \I__17800\ : LocalMux
    port map (
            O => \N__71883\,
            I => \N__71851\
        );

    \I__17799\ : Span4Mux_v
    port map (
            O => \N__71876\,
            I => \N__71846\
        );

    \I__17798\ : Span4Mux_v
    port map (
            O => \N__71871\,
            I => \N__71846\
        );

    \I__17797\ : InMux
    port map (
            O => \N__71870\,
            I => \N__71839\
        );

    \I__17796\ : InMux
    port map (
            O => \N__71869\,
            I => \N__71839\
        );

    \I__17795\ : InMux
    port map (
            O => \N__71868\,
            I => \N__71839\
        );

    \I__17794\ : Span4Mux_v
    port map (
            O => \N__71863\,
            I => \N__71836\
        );

    \I__17793\ : InMux
    port map (
            O => \N__71860\,
            I => \N__71833\
        );

    \I__17792\ : Span4Mux_h
    port map (
            O => \N__71857\,
            I => \N__71830\
        );

    \I__17791\ : Sp12to4
    port map (
            O => \N__71854\,
            I => \N__71825\
        );

    \I__17790\ : Span12Mux_h
    port map (
            O => \N__71851\,
            I => \N__71825\
        );

    \I__17789\ : Span4Mux_h
    port map (
            O => \N__71846\,
            I => \N__71822\
        );

    \I__17788\ : LocalMux
    port map (
            O => \N__71839\,
            I => \N__71817\
        );

    \I__17787\ : Span4Mux_h
    port map (
            O => \N__71836\,
            I => \N__71817\
        );

    \I__17786\ : LocalMux
    port map (
            O => \N__71833\,
            I => \c0.n19107\
        );

    \I__17785\ : Odrv4
    port map (
            O => \N__71830\,
            I => \c0.n19107\
        );

    \I__17784\ : Odrv12
    port map (
            O => \N__71825\,
            I => \c0.n19107\
        );

    \I__17783\ : Odrv4
    port map (
            O => \N__71822\,
            I => \c0.n19107\
        );

    \I__17782\ : Odrv4
    port map (
            O => \N__71817\,
            I => \c0.n19107\
        );

    \I__17781\ : CascadeMux
    port map (
            O => \N__71806\,
            I => \N__71803\
        );

    \I__17780\ : InMux
    port map (
            O => \N__71803\,
            I => \N__71797\
        );

    \I__17779\ : InMux
    port map (
            O => \N__71802\,
            I => \N__71794\
        );

    \I__17778\ : InMux
    port map (
            O => \N__71801\,
            I => \N__71788\
        );

    \I__17777\ : InMux
    port map (
            O => \N__71800\,
            I => \N__71783\
        );

    \I__17776\ : LocalMux
    port map (
            O => \N__71797\,
            I => \N__71770\
        );

    \I__17775\ : LocalMux
    port map (
            O => \N__71794\,
            I => \N__71770\
        );

    \I__17774\ : InMux
    port map (
            O => \N__71793\,
            I => \N__71767\
        );

    \I__17773\ : CascadeMux
    port map (
            O => \N__71792\,
            I => \N__71763\
        );

    \I__17772\ : InMux
    port map (
            O => \N__71791\,
            I => \N__71759\
        );

    \I__17771\ : LocalMux
    port map (
            O => \N__71788\,
            I => \N__71756\
        );

    \I__17770\ : InMux
    port map (
            O => \N__71787\,
            I => \N__71749\
        );

    \I__17769\ : InMux
    port map (
            O => \N__71786\,
            I => \N__71749\
        );

    \I__17768\ : LocalMux
    port map (
            O => \N__71783\,
            I => \N__71746\
        );

    \I__17767\ : CascadeMux
    port map (
            O => \N__71782\,
            I => \N__71741\
        );

    \I__17766\ : CascadeMux
    port map (
            O => \N__71781\,
            I => \N__71735\
        );

    \I__17765\ : InMux
    port map (
            O => \N__71780\,
            I => \N__71729\
        );

    \I__17764\ : InMux
    port map (
            O => \N__71779\,
            I => \N__71729\
        );

    \I__17763\ : InMux
    port map (
            O => \N__71778\,
            I => \N__71726\
        );

    \I__17762\ : InMux
    port map (
            O => \N__71777\,
            I => \N__71723\
        );

    \I__17761\ : InMux
    port map (
            O => \N__71776\,
            I => \N__71718\
        );

    \I__17760\ : InMux
    port map (
            O => \N__71775\,
            I => \N__71718\
        );

    \I__17759\ : Span4Mux_v
    port map (
            O => \N__71770\,
            I => \N__71713\
        );

    \I__17758\ : LocalMux
    port map (
            O => \N__71767\,
            I => \N__71713\
        );

    \I__17757\ : InMux
    port map (
            O => \N__71766\,
            I => \N__71710\
        );

    \I__17756\ : InMux
    port map (
            O => \N__71763\,
            I => \N__71707\
        );

    \I__17755\ : InMux
    port map (
            O => \N__71762\,
            I => \N__71704\
        );

    \I__17754\ : LocalMux
    port map (
            O => \N__71759\,
            I => \N__71701\
        );

    \I__17753\ : Span4Mux_v
    port map (
            O => \N__71756\,
            I => \N__71698\
        );

    \I__17752\ : InMux
    port map (
            O => \N__71755\,
            I => \N__71693\
        );

    \I__17751\ : InMux
    port map (
            O => \N__71754\,
            I => \N__71693\
        );

    \I__17750\ : LocalMux
    port map (
            O => \N__71749\,
            I => \N__71688\
        );

    \I__17749\ : Span4Mux_h
    port map (
            O => \N__71746\,
            I => \N__71688\
        );

    \I__17748\ : InMux
    port map (
            O => \N__71745\,
            I => \N__71681\
        );

    \I__17747\ : InMux
    port map (
            O => \N__71744\,
            I => \N__71681\
        );

    \I__17746\ : InMux
    port map (
            O => \N__71741\,
            I => \N__71681\
        );

    \I__17745\ : InMux
    port map (
            O => \N__71740\,
            I => \N__71678\
        );

    \I__17744\ : InMux
    port map (
            O => \N__71739\,
            I => \N__71671\
        );

    \I__17743\ : InMux
    port map (
            O => \N__71738\,
            I => \N__71671\
        );

    \I__17742\ : InMux
    port map (
            O => \N__71735\,
            I => \N__71671\
        );

    \I__17741\ : InMux
    port map (
            O => \N__71734\,
            I => \N__71668\
        );

    \I__17740\ : LocalMux
    port map (
            O => \N__71729\,
            I => \N__71665\
        );

    \I__17739\ : LocalMux
    port map (
            O => \N__71726\,
            I => \N__71662\
        );

    \I__17738\ : LocalMux
    port map (
            O => \N__71723\,
            I => \N__71659\
        );

    \I__17737\ : LocalMux
    port map (
            O => \N__71718\,
            I => \N__71656\
        );

    \I__17736\ : Span4Mux_h
    port map (
            O => \N__71713\,
            I => \N__71653\
        );

    \I__17735\ : LocalMux
    port map (
            O => \N__71710\,
            I => \N__71650\
        );

    \I__17734\ : LocalMux
    port map (
            O => \N__71707\,
            I => \N__71647\
        );

    \I__17733\ : LocalMux
    port map (
            O => \N__71704\,
            I => \N__71644\
        );

    \I__17732\ : Span4Mux_v
    port map (
            O => \N__71701\,
            I => \N__71641\
        );

    \I__17731\ : Span4Mux_h
    port map (
            O => \N__71698\,
            I => \N__71636\
        );

    \I__17730\ : LocalMux
    port map (
            O => \N__71693\,
            I => \N__71636\
        );

    \I__17729\ : Span4Mux_h
    port map (
            O => \N__71688\,
            I => \N__71633\
        );

    \I__17728\ : LocalMux
    port map (
            O => \N__71681\,
            I => \N__71630\
        );

    \I__17727\ : LocalMux
    port map (
            O => \N__71678\,
            I => \N__71625\
        );

    \I__17726\ : LocalMux
    port map (
            O => \N__71671\,
            I => \N__71625\
        );

    \I__17725\ : LocalMux
    port map (
            O => \N__71668\,
            I => \N__71620\
        );

    \I__17724\ : Span4Mux_h
    port map (
            O => \N__71665\,
            I => \N__71615\
        );

    \I__17723\ : Span4Mux_v
    port map (
            O => \N__71662\,
            I => \N__71615\
        );

    \I__17722\ : Span4Mux_h
    port map (
            O => \N__71659\,
            I => \N__71612\
        );

    \I__17721\ : Span4Mux_h
    port map (
            O => \N__71656\,
            I => \N__71607\
        );

    \I__17720\ : Span4Mux_h
    port map (
            O => \N__71653\,
            I => \N__71607\
        );

    \I__17719\ : Span4Mux_h
    port map (
            O => \N__71650\,
            I => \N__71604\
        );

    \I__17718\ : Span4Mux_h
    port map (
            O => \N__71647\,
            I => \N__71601\
        );

    \I__17717\ : Span4Mux_v
    port map (
            O => \N__71644\,
            I => \N__71594\
        );

    \I__17716\ : Span4Mux_v
    port map (
            O => \N__71641\,
            I => \N__71594\
        );

    \I__17715\ : Span4Mux_h
    port map (
            O => \N__71636\,
            I => \N__71594\
        );

    \I__17714\ : Span4Mux_v
    port map (
            O => \N__71633\,
            I => \N__71591\
        );

    \I__17713\ : Span12Mux_v
    port map (
            O => \N__71630\,
            I => \N__71586\
        );

    \I__17712\ : Span12Mux_v
    port map (
            O => \N__71625\,
            I => \N__71586\
        );

    \I__17711\ : InMux
    port map (
            O => \N__71624\,
            I => \N__71583\
        );

    \I__17710\ : InMux
    port map (
            O => \N__71623\,
            I => \N__71580\
        );

    \I__17709\ : Span4Mux_v
    port map (
            O => \N__71620\,
            I => \N__71573\
        );

    \I__17708\ : Span4Mux_h
    port map (
            O => \N__71615\,
            I => \N__71573\
        );

    \I__17707\ : Span4Mux_v
    port map (
            O => \N__71612\,
            I => \N__71573\
        );

    \I__17706\ : Span4Mux_h
    port map (
            O => \N__71607\,
            I => \N__71570\
        );

    \I__17705\ : Span4Mux_h
    port map (
            O => \N__71604\,
            I => \N__71563\
        );

    \I__17704\ : Span4Mux_v
    port map (
            O => \N__71601\,
            I => \N__71563\
        );

    \I__17703\ : Span4Mux_h
    port map (
            O => \N__71594\,
            I => \N__71563\
        );

    \I__17702\ : Odrv4
    port map (
            O => \N__71591\,
            I => \c0.n12_adj_3361\
        );

    \I__17701\ : Odrv12
    port map (
            O => \N__71586\,
            I => \c0.n12_adj_3361\
        );

    \I__17700\ : LocalMux
    port map (
            O => \N__71583\,
            I => \c0.n12_adj_3361\
        );

    \I__17699\ : LocalMux
    port map (
            O => \N__71580\,
            I => \c0.n12_adj_3361\
        );

    \I__17698\ : Odrv4
    port map (
            O => \N__71573\,
            I => \c0.n12_adj_3361\
        );

    \I__17697\ : Odrv4
    port map (
            O => \N__71570\,
            I => \c0.n12_adj_3361\
        );

    \I__17696\ : Odrv4
    port map (
            O => \N__71563\,
            I => \c0.n12_adj_3361\
        );

    \I__17695\ : InMux
    port map (
            O => \N__71548\,
            I => \N__71544\
        );

    \I__17694\ : InMux
    port map (
            O => \N__71547\,
            I => \N__71540\
        );

    \I__17693\ : LocalMux
    port map (
            O => \N__71544\,
            I => \N__71537\
        );

    \I__17692\ : InMux
    port map (
            O => \N__71543\,
            I => \N__71531\
        );

    \I__17691\ : LocalMux
    port map (
            O => \N__71540\,
            I => \N__71528\
        );

    \I__17690\ : Span4Mux_v
    port map (
            O => \N__71537\,
            I => \N__71521\
        );

    \I__17689\ : InMux
    port map (
            O => \N__71536\,
            I => \N__71518\
        );

    \I__17688\ : InMux
    port map (
            O => \N__71535\,
            I => \N__71513\
        );

    \I__17687\ : InMux
    port map (
            O => \N__71534\,
            I => \N__71513\
        );

    \I__17686\ : LocalMux
    port map (
            O => \N__71531\,
            I => \N__71510\
        );

    \I__17685\ : Span4Mux_v
    port map (
            O => \N__71528\,
            I => \N__71507\
        );

    \I__17684\ : InMux
    port map (
            O => \N__71527\,
            I => \N__71500\
        );

    \I__17683\ : InMux
    port map (
            O => \N__71526\,
            I => \N__71497\
        );

    \I__17682\ : CascadeMux
    port map (
            O => \N__71525\,
            I => \N__71493\
        );

    \I__17681\ : InMux
    port map (
            O => \N__71524\,
            I => \N__71489\
        );

    \I__17680\ : Span4Mux_h
    port map (
            O => \N__71521\,
            I => \N__71480\
        );

    \I__17679\ : LocalMux
    port map (
            O => \N__71518\,
            I => \N__71480\
        );

    \I__17678\ : LocalMux
    port map (
            O => \N__71513\,
            I => \N__71473\
        );

    \I__17677\ : Span4Mux_v
    port map (
            O => \N__71510\,
            I => \N__71473\
        );

    \I__17676\ : Span4Mux_h
    port map (
            O => \N__71507\,
            I => \N__71473\
        );

    \I__17675\ : InMux
    port map (
            O => \N__71506\,
            I => \N__71470\
        );

    \I__17674\ : InMux
    port map (
            O => \N__71505\,
            I => \N__71467\
        );

    \I__17673\ : InMux
    port map (
            O => \N__71504\,
            I => \N__71459\
        );

    \I__17672\ : InMux
    port map (
            O => \N__71503\,
            I => \N__71459\
        );

    \I__17671\ : LocalMux
    port map (
            O => \N__71500\,
            I => \N__71456\
        );

    \I__17670\ : LocalMux
    port map (
            O => \N__71497\,
            I => \N__71453\
        );

    \I__17669\ : InMux
    port map (
            O => \N__71496\,
            I => \N__71450\
        );

    \I__17668\ : InMux
    port map (
            O => \N__71493\,
            I => \N__71445\
        );

    \I__17667\ : InMux
    port map (
            O => \N__71492\,
            I => \N__71445\
        );

    \I__17666\ : LocalMux
    port map (
            O => \N__71489\,
            I => \N__71442\
        );

    \I__17665\ : InMux
    port map (
            O => \N__71488\,
            I => \N__71437\
        );

    \I__17664\ : InMux
    port map (
            O => \N__71487\,
            I => \N__71437\
        );

    \I__17663\ : InMux
    port map (
            O => \N__71486\,
            I => \N__71433\
        );

    \I__17662\ : InMux
    port map (
            O => \N__71485\,
            I => \N__71430\
        );

    \I__17661\ : Span4Mux_v
    port map (
            O => \N__71480\,
            I => \N__71427\
        );

    \I__17660\ : Span4Mux_h
    port map (
            O => \N__71473\,
            I => \N__71420\
        );

    \I__17659\ : LocalMux
    port map (
            O => \N__71470\,
            I => \N__71420\
        );

    \I__17658\ : LocalMux
    port map (
            O => \N__71467\,
            I => \N__71420\
        );

    \I__17657\ : InMux
    port map (
            O => \N__71466\,
            I => \N__71412\
        );

    \I__17656\ : InMux
    port map (
            O => \N__71465\,
            I => \N__71412\
        );

    \I__17655\ : InMux
    port map (
            O => \N__71464\,
            I => \N__71412\
        );

    \I__17654\ : LocalMux
    port map (
            O => \N__71459\,
            I => \N__71409\
        );

    \I__17653\ : Span4Mux_v
    port map (
            O => \N__71456\,
            I => \N__71404\
        );

    \I__17652\ : Span4Mux_v
    port map (
            O => \N__71453\,
            I => \N__71404\
        );

    \I__17651\ : LocalMux
    port map (
            O => \N__71450\,
            I => \N__71399\
        );

    \I__17650\ : LocalMux
    port map (
            O => \N__71445\,
            I => \N__71399\
        );

    \I__17649\ : Span4Mux_v
    port map (
            O => \N__71442\,
            I => \N__71394\
        );

    \I__17648\ : LocalMux
    port map (
            O => \N__71437\,
            I => \N__71394\
        );

    \I__17647\ : InMux
    port map (
            O => \N__71436\,
            I => \N__71390\
        );

    \I__17646\ : LocalMux
    port map (
            O => \N__71433\,
            I => \N__71385\
        );

    \I__17645\ : LocalMux
    port map (
            O => \N__71430\,
            I => \N__71385\
        );

    \I__17644\ : Sp12to4
    port map (
            O => \N__71427\,
            I => \N__71380\
        );

    \I__17643\ : Sp12to4
    port map (
            O => \N__71420\,
            I => \N__71380\
        );

    \I__17642\ : InMux
    port map (
            O => \N__71419\,
            I => \N__71377\
        );

    \I__17641\ : LocalMux
    port map (
            O => \N__71412\,
            I => \N__71369\
        );

    \I__17640\ : Span12Mux_v
    port map (
            O => \N__71409\,
            I => \N__71369\
        );

    \I__17639\ : Span4Mux_h
    port map (
            O => \N__71404\,
            I => \N__71362\
        );

    \I__17638\ : Span4Mux_h
    port map (
            O => \N__71399\,
            I => \N__71362\
        );

    \I__17637\ : Span4Mux_v
    port map (
            O => \N__71394\,
            I => \N__71362\
        );

    \I__17636\ : InMux
    port map (
            O => \N__71393\,
            I => \N__71359\
        );

    \I__17635\ : LocalMux
    port map (
            O => \N__71390\,
            I => \N__71356\
        );

    \I__17634\ : Span4Mux_h
    port map (
            O => \N__71385\,
            I => \N__71353\
        );

    \I__17633\ : Span12Mux_h
    port map (
            O => \N__71380\,
            I => \N__71350\
        );

    \I__17632\ : LocalMux
    port map (
            O => \N__71377\,
            I => \N__71344\
        );

    \I__17631\ : InMux
    port map (
            O => \N__71376\,
            I => \N__71341\
        );

    \I__17630\ : InMux
    port map (
            O => \N__71375\,
            I => \N__71336\
        );

    \I__17629\ : InMux
    port map (
            O => \N__71374\,
            I => \N__71336\
        );

    \I__17628\ : Span12Mux_h
    port map (
            O => \N__71369\,
            I => \N__71333\
        );

    \I__17627\ : Sp12to4
    port map (
            O => \N__71362\,
            I => \N__71330\
        );

    \I__17626\ : LocalMux
    port map (
            O => \N__71359\,
            I => \N__71323\
        );

    \I__17625\ : Span4Mux_h
    port map (
            O => \N__71356\,
            I => \N__71323\
        );

    \I__17624\ : Span4Mux_v
    port map (
            O => \N__71353\,
            I => \N__71323\
        );

    \I__17623\ : Span12Mux_v
    port map (
            O => \N__71350\,
            I => \N__71320\
        );

    \I__17622\ : InMux
    port map (
            O => \N__71349\,
            I => \N__71315\
        );

    \I__17621\ : InMux
    port map (
            O => \N__71348\,
            I => \N__71315\
        );

    \I__17620\ : InMux
    port map (
            O => \N__71347\,
            I => \N__71312\
        );

    \I__17619\ : Span4Mux_h
    port map (
            O => \N__71344\,
            I => \N__71307\
        );

    \I__17618\ : LocalMux
    port map (
            O => \N__71341\,
            I => \N__71307\
        );

    \I__17617\ : LocalMux
    port map (
            O => \N__71336\,
            I => \N__71302\
        );

    \I__17616\ : Span12Mux_v
    port map (
            O => \N__71333\,
            I => \N__71302\
        );

    \I__17615\ : Span12Mux_h
    port map (
            O => \N__71330\,
            I => \N__71295\
        );

    \I__17614\ : Sp12to4
    port map (
            O => \N__71323\,
            I => \N__71295\
        );

    \I__17613\ : Span12Mux_h
    port map (
            O => \N__71320\,
            I => \N__71295\
        );

    \I__17612\ : LocalMux
    port map (
            O => \N__71315\,
            I => rx_data_1
        );

    \I__17611\ : LocalMux
    port map (
            O => \N__71312\,
            I => rx_data_1
        );

    \I__17610\ : Odrv4
    port map (
            O => \N__71307\,
            I => rx_data_1
        );

    \I__17609\ : Odrv12
    port map (
            O => \N__71302\,
            I => rx_data_1
        );

    \I__17608\ : Odrv12
    port map (
            O => \N__71295\,
            I => rx_data_1
        );

    \I__17607\ : CascadeMux
    port map (
            O => \N__71284\,
            I => \N__71280\
        );

    \I__17606\ : InMux
    port map (
            O => \N__71283\,
            I => \N__71277\
        );

    \I__17605\ : InMux
    port map (
            O => \N__71280\,
            I => \N__71274\
        );

    \I__17604\ : LocalMux
    port map (
            O => \N__71277\,
            I => \N__71270\
        );

    \I__17603\ : LocalMux
    port map (
            O => \N__71274\,
            I => \N__71267\
        );

    \I__17602\ : CascadeMux
    port map (
            O => \N__71273\,
            I => \N__71262\
        );

    \I__17601\ : Span4Mux_h
    port map (
            O => \N__71270\,
            I => \N__71259\
        );

    \I__17600\ : Span4Mux_h
    port map (
            O => \N__71267\,
            I => \N__71256\
        );

    \I__17599\ : InMux
    port map (
            O => \N__71266\,
            I => \N__71251\
        );

    \I__17598\ : InMux
    port map (
            O => \N__71265\,
            I => \N__71251\
        );

    \I__17597\ : InMux
    port map (
            O => \N__71262\,
            I => \N__71248\
        );

    \I__17596\ : Span4Mux_h
    port map (
            O => \N__71259\,
            I => \N__71245\
        );

    \I__17595\ : Span4Mux_h
    port map (
            O => \N__71256\,
            I => \N__71240\
        );

    \I__17594\ : LocalMux
    port map (
            O => \N__71251\,
            I => \N__71240\
        );

    \I__17593\ : LocalMux
    port map (
            O => \N__71248\,
            I => \c0.data_in_frame_21_1\
        );

    \I__17592\ : Odrv4
    port map (
            O => \N__71245\,
            I => \c0.data_in_frame_21_1\
        );

    \I__17591\ : Odrv4
    port map (
            O => \N__71240\,
            I => \c0.data_in_frame_21_1\
        );

    \I__17590\ : ClkMux
    port map (
            O => \N__71233\,
            I => \N__70504\
        );

    \I__17589\ : ClkMux
    port map (
            O => \N__71232\,
            I => \N__70504\
        );

    \I__17588\ : ClkMux
    port map (
            O => \N__71231\,
            I => \N__70504\
        );

    \I__17587\ : ClkMux
    port map (
            O => \N__71230\,
            I => \N__70504\
        );

    \I__17586\ : ClkMux
    port map (
            O => \N__71229\,
            I => \N__70504\
        );

    \I__17585\ : ClkMux
    port map (
            O => \N__71228\,
            I => \N__70504\
        );

    \I__17584\ : ClkMux
    port map (
            O => \N__71227\,
            I => \N__70504\
        );

    \I__17583\ : ClkMux
    port map (
            O => \N__71226\,
            I => \N__70504\
        );

    \I__17582\ : ClkMux
    port map (
            O => \N__71225\,
            I => \N__70504\
        );

    \I__17581\ : ClkMux
    port map (
            O => \N__71224\,
            I => \N__70504\
        );

    \I__17580\ : ClkMux
    port map (
            O => \N__71223\,
            I => \N__70504\
        );

    \I__17579\ : ClkMux
    port map (
            O => \N__71222\,
            I => \N__70504\
        );

    \I__17578\ : ClkMux
    port map (
            O => \N__71221\,
            I => \N__70504\
        );

    \I__17577\ : ClkMux
    port map (
            O => \N__71220\,
            I => \N__70504\
        );

    \I__17576\ : ClkMux
    port map (
            O => \N__71219\,
            I => \N__70504\
        );

    \I__17575\ : ClkMux
    port map (
            O => \N__71218\,
            I => \N__70504\
        );

    \I__17574\ : ClkMux
    port map (
            O => \N__71217\,
            I => \N__70504\
        );

    \I__17573\ : ClkMux
    port map (
            O => \N__71216\,
            I => \N__70504\
        );

    \I__17572\ : ClkMux
    port map (
            O => \N__71215\,
            I => \N__70504\
        );

    \I__17571\ : ClkMux
    port map (
            O => \N__71214\,
            I => \N__70504\
        );

    \I__17570\ : ClkMux
    port map (
            O => \N__71213\,
            I => \N__70504\
        );

    \I__17569\ : ClkMux
    port map (
            O => \N__71212\,
            I => \N__70504\
        );

    \I__17568\ : ClkMux
    port map (
            O => \N__71211\,
            I => \N__70504\
        );

    \I__17567\ : ClkMux
    port map (
            O => \N__71210\,
            I => \N__70504\
        );

    \I__17566\ : ClkMux
    port map (
            O => \N__71209\,
            I => \N__70504\
        );

    \I__17565\ : ClkMux
    port map (
            O => \N__71208\,
            I => \N__70504\
        );

    \I__17564\ : ClkMux
    port map (
            O => \N__71207\,
            I => \N__70504\
        );

    \I__17563\ : ClkMux
    port map (
            O => \N__71206\,
            I => \N__70504\
        );

    \I__17562\ : ClkMux
    port map (
            O => \N__71205\,
            I => \N__70504\
        );

    \I__17561\ : ClkMux
    port map (
            O => \N__71204\,
            I => \N__70504\
        );

    \I__17560\ : ClkMux
    port map (
            O => \N__71203\,
            I => \N__70504\
        );

    \I__17559\ : ClkMux
    port map (
            O => \N__71202\,
            I => \N__70504\
        );

    \I__17558\ : ClkMux
    port map (
            O => \N__71201\,
            I => \N__70504\
        );

    \I__17557\ : ClkMux
    port map (
            O => \N__71200\,
            I => \N__70504\
        );

    \I__17556\ : ClkMux
    port map (
            O => \N__71199\,
            I => \N__70504\
        );

    \I__17555\ : ClkMux
    port map (
            O => \N__71198\,
            I => \N__70504\
        );

    \I__17554\ : ClkMux
    port map (
            O => \N__71197\,
            I => \N__70504\
        );

    \I__17553\ : ClkMux
    port map (
            O => \N__71196\,
            I => \N__70504\
        );

    \I__17552\ : ClkMux
    port map (
            O => \N__71195\,
            I => \N__70504\
        );

    \I__17551\ : ClkMux
    port map (
            O => \N__71194\,
            I => \N__70504\
        );

    \I__17550\ : ClkMux
    port map (
            O => \N__71193\,
            I => \N__70504\
        );

    \I__17549\ : ClkMux
    port map (
            O => \N__71192\,
            I => \N__70504\
        );

    \I__17548\ : ClkMux
    port map (
            O => \N__71191\,
            I => \N__70504\
        );

    \I__17547\ : ClkMux
    port map (
            O => \N__71190\,
            I => \N__70504\
        );

    \I__17546\ : ClkMux
    port map (
            O => \N__71189\,
            I => \N__70504\
        );

    \I__17545\ : ClkMux
    port map (
            O => \N__71188\,
            I => \N__70504\
        );

    \I__17544\ : ClkMux
    port map (
            O => \N__71187\,
            I => \N__70504\
        );

    \I__17543\ : ClkMux
    port map (
            O => \N__71186\,
            I => \N__70504\
        );

    \I__17542\ : ClkMux
    port map (
            O => \N__71185\,
            I => \N__70504\
        );

    \I__17541\ : ClkMux
    port map (
            O => \N__71184\,
            I => \N__70504\
        );

    \I__17540\ : ClkMux
    port map (
            O => \N__71183\,
            I => \N__70504\
        );

    \I__17539\ : ClkMux
    port map (
            O => \N__71182\,
            I => \N__70504\
        );

    \I__17538\ : ClkMux
    port map (
            O => \N__71181\,
            I => \N__70504\
        );

    \I__17537\ : ClkMux
    port map (
            O => \N__71180\,
            I => \N__70504\
        );

    \I__17536\ : ClkMux
    port map (
            O => \N__71179\,
            I => \N__70504\
        );

    \I__17535\ : ClkMux
    port map (
            O => \N__71178\,
            I => \N__70504\
        );

    \I__17534\ : ClkMux
    port map (
            O => \N__71177\,
            I => \N__70504\
        );

    \I__17533\ : ClkMux
    port map (
            O => \N__71176\,
            I => \N__70504\
        );

    \I__17532\ : ClkMux
    port map (
            O => \N__71175\,
            I => \N__70504\
        );

    \I__17531\ : ClkMux
    port map (
            O => \N__71174\,
            I => \N__70504\
        );

    \I__17530\ : ClkMux
    port map (
            O => \N__71173\,
            I => \N__70504\
        );

    \I__17529\ : ClkMux
    port map (
            O => \N__71172\,
            I => \N__70504\
        );

    \I__17528\ : ClkMux
    port map (
            O => \N__71171\,
            I => \N__70504\
        );

    \I__17527\ : ClkMux
    port map (
            O => \N__71170\,
            I => \N__70504\
        );

    \I__17526\ : ClkMux
    port map (
            O => \N__71169\,
            I => \N__70504\
        );

    \I__17525\ : ClkMux
    port map (
            O => \N__71168\,
            I => \N__70504\
        );

    \I__17524\ : ClkMux
    port map (
            O => \N__71167\,
            I => \N__70504\
        );

    \I__17523\ : ClkMux
    port map (
            O => \N__71166\,
            I => \N__70504\
        );

    \I__17522\ : ClkMux
    port map (
            O => \N__71165\,
            I => \N__70504\
        );

    \I__17521\ : ClkMux
    port map (
            O => \N__71164\,
            I => \N__70504\
        );

    \I__17520\ : ClkMux
    port map (
            O => \N__71163\,
            I => \N__70504\
        );

    \I__17519\ : ClkMux
    port map (
            O => \N__71162\,
            I => \N__70504\
        );

    \I__17518\ : ClkMux
    port map (
            O => \N__71161\,
            I => \N__70504\
        );

    \I__17517\ : ClkMux
    port map (
            O => \N__71160\,
            I => \N__70504\
        );

    \I__17516\ : ClkMux
    port map (
            O => \N__71159\,
            I => \N__70504\
        );

    \I__17515\ : ClkMux
    port map (
            O => \N__71158\,
            I => \N__70504\
        );

    \I__17514\ : ClkMux
    port map (
            O => \N__71157\,
            I => \N__70504\
        );

    \I__17513\ : ClkMux
    port map (
            O => \N__71156\,
            I => \N__70504\
        );

    \I__17512\ : ClkMux
    port map (
            O => \N__71155\,
            I => \N__70504\
        );

    \I__17511\ : ClkMux
    port map (
            O => \N__71154\,
            I => \N__70504\
        );

    \I__17510\ : ClkMux
    port map (
            O => \N__71153\,
            I => \N__70504\
        );

    \I__17509\ : ClkMux
    port map (
            O => \N__71152\,
            I => \N__70504\
        );

    \I__17508\ : ClkMux
    port map (
            O => \N__71151\,
            I => \N__70504\
        );

    \I__17507\ : ClkMux
    port map (
            O => \N__71150\,
            I => \N__70504\
        );

    \I__17506\ : ClkMux
    port map (
            O => \N__71149\,
            I => \N__70504\
        );

    \I__17505\ : ClkMux
    port map (
            O => \N__71148\,
            I => \N__70504\
        );

    \I__17504\ : ClkMux
    port map (
            O => \N__71147\,
            I => \N__70504\
        );

    \I__17503\ : ClkMux
    port map (
            O => \N__71146\,
            I => \N__70504\
        );

    \I__17502\ : ClkMux
    port map (
            O => \N__71145\,
            I => \N__70504\
        );

    \I__17501\ : ClkMux
    port map (
            O => \N__71144\,
            I => \N__70504\
        );

    \I__17500\ : ClkMux
    port map (
            O => \N__71143\,
            I => \N__70504\
        );

    \I__17499\ : ClkMux
    port map (
            O => \N__71142\,
            I => \N__70504\
        );

    \I__17498\ : ClkMux
    port map (
            O => \N__71141\,
            I => \N__70504\
        );

    \I__17497\ : ClkMux
    port map (
            O => \N__71140\,
            I => \N__70504\
        );

    \I__17496\ : ClkMux
    port map (
            O => \N__71139\,
            I => \N__70504\
        );

    \I__17495\ : ClkMux
    port map (
            O => \N__71138\,
            I => \N__70504\
        );

    \I__17494\ : ClkMux
    port map (
            O => \N__71137\,
            I => \N__70504\
        );

    \I__17493\ : ClkMux
    port map (
            O => \N__71136\,
            I => \N__70504\
        );

    \I__17492\ : ClkMux
    port map (
            O => \N__71135\,
            I => \N__70504\
        );

    \I__17491\ : ClkMux
    port map (
            O => \N__71134\,
            I => \N__70504\
        );

    \I__17490\ : ClkMux
    port map (
            O => \N__71133\,
            I => \N__70504\
        );

    \I__17489\ : ClkMux
    port map (
            O => \N__71132\,
            I => \N__70504\
        );

    \I__17488\ : ClkMux
    port map (
            O => \N__71131\,
            I => \N__70504\
        );

    \I__17487\ : ClkMux
    port map (
            O => \N__71130\,
            I => \N__70504\
        );

    \I__17486\ : ClkMux
    port map (
            O => \N__71129\,
            I => \N__70504\
        );

    \I__17485\ : ClkMux
    port map (
            O => \N__71128\,
            I => \N__70504\
        );

    \I__17484\ : ClkMux
    port map (
            O => \N__71127\,
            I => \N__70504\
        );

    \I__17483\ : ClkMux
    port map (
            O => \N__71126\,
            I => \N__70504\
        );

    \I__17482\ : ClkMux
    port map (
            O => \N__71125\,
            I => \N__70504\
        );

    \I__17481\ : ClkMux
    port map (
            O => \N__71124\,
            I => \N__70504\
        );

    \I__17480\ : ClkMux
    port map (
            O => \N__71123\,
            I => \N__70504\
        );

    \I__17479\ : ClkMux
    port map (
            O => \N__71122\,
            I => \N__70504\
        );

    \I__17478\ : ClkMux
    port map (
            O => \N__71121\,
            I => \N__70504\
        );

    \I__17477\ : ClkMux
    port map (
            O => \N__71120\,
            I => \N__70504\
        );

    \I__17476\ : ClkMux
    port map (
            O => \N__71119\,
            I => \N__70504\
        );

    \I__17475\ : ClkMux
    port map (
            O => \N__71118\,
            I => \N__70504\
        );

    \I__17474\ : ClkMux
    port map (
            O => \N__71117\,
            I => \N__70504\
        );

    \I__17473\ : ClkMux
    port map (
            O => \N__71116\,
            I => \N__70504\
        );

    \I__17472\ : ClkMux
    port map (
            O => \N__71115\,
            I => \N__70504\
        );

    \I__17471\ : ClkMux
    port map (
            O => \N__71114\,
            I => \N__70504\
        );

    \I__17470\ : ClkMux
    port map (
            O => \N__71113\,
            I => \N__70504\
        );

    \I__17469\ : ClkMux
    port map (
            O => \N__71112\,
            I => \N__70504\
        );

    \I__17468\ : ClkMux
    port map (
            O => \N__71111\,
            I => \N__70504\
        );

    \I__17467\ : ClkMux
    port map (
            O => \N__71110\,
            I => \N__70504\
        );

    \I__17466\ : ClkMux
    port map (
            O => \N__71109\,
            I => \N__70504\
        );

    \I__17465\ : ClkMux
    port map (
            O => \N__71108\,
            I => \N__70504\
        );

    \I__17464\ : ClkMux
    port map (
            O => \N__71107\,
            I => \N__70504\
        );

    \I__17463\ : ClkMux
    port map (
            O => \N__71106\,
            I => \N__70504\
        );

    \I__17462\ : ClkMux
    port map (
            O => \N__71105\,
            I => \N__70504\
        );

    \I__17461\ : ClkMux
    port map (
            O => \N__71104\,
            I => \N__70504\
        );

    \I__17460\ : ClkMux
    port map (
            O => \N__71103\,
            I => \N__70504\
        );

    \I__17459\ : ClkMux
    port map (
            O => \N__71102\,
            I => \N__70504\
        );

    \I__17458\ : ClkMux
    port map (
            O => \N__71101\,
            I => \N__70504\
        );

    \I__17457\ : ClkMux
    port map (
            O => \N__71100\,
            I => \N__70504\
        );

    \I__17456\ : ClkMux
    port map (
            O => \N__71099\,
            I => \N__70504\
        );

    \I__17455\ : ClkMux
    port map (
            O => \N__71098\,
            I => \N__70504\
        );

    \I__17454\ : ClkMux
    port map (
            O => \N__71097\,
            I => \N__70504\
        );

    \I__17453\ : ClkMux
    port map (
            O => \N__71096\,
            I => \N__70504\
        );

    \I__17452\ : ClkMux
    port map (
            O => \N__71095\,
            I => \N__70504\
        );

    \I__17451\ : ClkMux
    port map (
            O => \N__71094\,
            I => \N__70504\
        );

    \I__17450\ : ClkMux
    port map (
            O => \N__71093\,
            I => \N__70504\
        );

    \I__17449\ : ClkMux
    port map (
            O => \N__71092\,
            I => \N__70504\
        );

    \I__17448\ : ClkMux
    port map (
            O => \N__71091\,
            I => \N__70504\
        );

    \I__17447\ : ClkMux
    port map (
            O => \N__71090\,
            I => \N__70504\
        );

    \I__17446\ : ClkMux
    port map (
            O => \N__71089\,
            I => \N__70504\
        );

    \I__17445\ : ClkMux
    port map (
            O => \N__71088\,
            I => \N__70504\
        );

    \I__17444\ : ClkMux
    port map (
            O => \N__71087\,
            I => \N__70504\
        );

    \I__17443\ : ClkMux
    port map (
            O => \N__71086\,
            I => \N__70504\
        );

    \I__17442\ : ClkMux
    port map (
            O => \N__71085\,
            I => \N__70504\
        );

    \I__17441\ : ClkMux
    port map (
            O => \N__71084\,
            I => \N__70504\
        );

    \I__17440\ : ClkMux
    port map (
            O => \N__71083\,
            I => \N__70504\
        );

    \I__17439\ : ClkMux
    port map (
            O => \N__71082\,
            I => \N__70504\
        );

    \I__17438\ : ClkMux
    port map (
            O => \N__71081\,
            I => \N__70504\
        );

    \I__17437\ : ClkMux
    port map (
            O => \N__71080\,
            I => \N__70504\
        );

    \I__17436\ : ClkMux
    port map (
            O => \N__71079\,
            I => \N__70504\
        );

    \I__17435\ : ClkMux
    port map (
            O => \N__71078\,
            I => \N__70504\
        );

    \I__17434\ : ClkMux
    port map (
            O => \N__71077\,
            I => \N__70504\
        );

    \I__17433\ : ClkMux
    port map (
            O => \N__71076\,
            I => \N__70504\
        );

    \I__17432\ : ClkMux
    port map (
            O => \N__71075\,
            I => \N__70504\
        );

    \I__17431\ : ClkMux
    port map (
            O => \N__71074\,
            I => \N__70504\
        );

    \I__17430\ : ClkMux
    port map (
            O => \N__71073\,
            I => \N__70504\
        );

    \I__17429\ : ClkMux
    port map (
            O => \N__71072\,
            I => \N__70504\
        );

    \I__17428\ : ClkMux
    port map (
            O => \N__71071\,
            I => \N__70504\
        );

    \I__17427\ : ClkMux
    port map (
            O => \N__71070\,
            I => \N__70504\
        );

    \I__17426\ : ClkMux
    port map (
            O => \N__71069\,
            I => \N__70504\
        );

    \I__17425\ : ClkMux
    port map (
            O => \N__71068\,
            I => \N__70504\
        );

    \I__17424\ : ClkMux
    port map (
            O => \N__71067\,
            I => \N__70504\
        );

    \I__17423\ : ClkMux
    port map (
            O => \N__71066\,
            I => \N__70504\
        );

    \I__17422\ : ClkMux
    port map (
            O => \N__71065\,
            I => \N__70504\
        );

    \I__17421\ : ClkMux
    port map (
            O => \N__71064\,
            I => \N__70504\
        );

    \I__17420\ : ClkMux
    port map (
            O => \N__71063\,
            I => \N__70504\
        );

    \I__17419\ : ClkMux
    port map (
            O => \N__71062\,
            I => \N__70504\
        );

    \I__17418\ : ClkMux
    port map (
            O => \N__71061\,
            I => \N__70504\
        );

    \I__17417\ : ClkMux
    port map (
            O => \N__71060\,
            I => \N__70504\
        );

    \I__17416\ : ClkMux
    port map (
            O => \N__71059\,
            I => \N__70504\
        );

    \I__17415\ : ClkMux
    port map (
            O => \N__71058\,
            I => \N__70504\
        );

    \I__17414\ : ClkMux
    port map (
            O => \N__71057\,
            I => \N__70504\
        );

    \I__17413\ : ClkMux
    port map (
            O => \N__71056\,
            I => \N__70504\
        );

    \I__17412\ : ClkMux
    port map (
            O => \N__71055\,
            I => \N__70504\
        );

    \I__17411\ : ClkMux
    port map (
            O => \N__71054\,
            I => \N__70504\
        );

    \I__17410\ : ClkMux
    port map (
            O => \N__71053\,
            I => \N__70504\
        );

    \I__17409\ : ClkMux
    port map (
            O => \N__71052\,
            I => \N__70504\
        );

    \I__17408\ : ClkMux
    port map (
            O => \N__71051\,
            I => \N__70504\
        );

    \I__17407\ : ClkMux
    port map (
            O => \N__71050\,
            I => \N__70504\
        );

    \I__17406\ : ClkMux
    port map (
            O => \N__71049\,
            I => \N__70504\
        );

    \I__17405\ : ClkMux
    port map (
            O => \N__71048\,
            I => \N__70504\
        );

    \I__17404\ : ClkMux
    port map (
            O => \N__71047\,
            I => \N__70504\
        );

    \I__17403\ : ClkMux
    port map (
            O => \N__71046\,
            I => \N__70504\
        );

    \I__17402\ : ClkMux
    port map (
            O => \N__71045\,
            I => \N__70504\
        );

    \I__17401\ : ClkMux
    port map (
            O => \N__71044\,
            I => \N__70504\
        );

    \I__17400\ : ClkMux
    port map (
            O => \N__71043\,
            I => \N__70504\
        );

    \I__17399\ : ClkMux
    port map (
            O => \N__71042\,
            I => \N__70504\
        );

    \I__17398\ : ClkMux
    port map (
            O => \N__71041\,
            I => \N__70504\
        );

    \I__17397\ : ClkMux
    port map (
            O => \N__71040\,
            I => \N__70504\
        );

    \I__17396\ : ClkMux
    port map (
            O => \N__71039\,
            I => \N__70504\
        );

    \I__17395\ : ClkMux
    port map (
            O => \N__71038\,
            I => \N__70504\
        );

    \I__17394\ : ClkMux
    port map (
            O => \N__71037\,
            I => \N__70504\
        );

    \I__17393\ : ClkMux
    port map (
            O => \N__71036\,
            I => \N__70504\
        );

    \I__17392\ : ClkMux
    port map (
            O => \N__71035\,
            I => \N__70504\
        );

    \I__17391\ : ClkMux
    port map (
            O => \N__71034\,
            I => \N__70504\
        );

    \I__17390\ : ClkMux
    port map (
            O => \N__71033\,
            I => \N__70504\
        );

    \I__17389\ : ClkMux
    port map (
            O => \N__71032\,
            I => \N__70504\
        );

    \I__17388\ : ClkMux
    port map (
            O => \N__71031\,
            I => \N__70504\
        );

    \I__17387\ : ClkMux
    port map (
            O => \N__71030\,
            I => \N__70504\
        );

    \I__17386\ : ClkMux
    port map (
            O => \N__71029\,
            I => \N__70504\
        );

    \I__17385\ : ClkMux
    port map (
            O => \N__71028\,
            I => \N__70504\
        );

    \I__17384\ : ClkMux
    port map (
            O => \N__71027\,
            I => \N__70504\
        );

    \I__17383\ : ClkMux
    port map (
            O => \N__71026\,
            I => \N__70504\
        );

    \I__17382\ : ClkMux
    port map (
            O => \N__71025\,
            I => \N__70504\
        );

    \I__17381\ : ClkMux
    port map (
            O => \N__71024\,
            I => \N__70504\
        );

    \I__17380\ : ClkMux
    port map (
            O => \N__71023\,
            I => \N__70504\
        );

    \I__17379\ : ClkMux
    port map (
            O => \N__71022\,
            I => \N__70504\
        );

    \I__17378\ : ClkMux
    port map (
            O => \N__71021\,
            I => \N__70504\
        );

    \I__17377\ : ClkMux
    port map (
            O => \N__71020\,
            I => \N__70504\
        );

    \I__17376\ : ClkMux
    port map (
            O => \N__71019\,
            I => \N__70504\
        );

    \I__17375\ : ClkMux
    port map (
            O => \N__71018\,
            I => \N__70504\
        );

    \I__17374\ : ClkMux
    port map (
            O => \N__71017\,
            I => \N__70504\
        );

    \I__17373\ : ClkMux
    port map (
            O => \N__71016\,
            I => \N__70504\
        );

    \I__17372\ : ClkMux
    port map (
            O => \N__71015\,
            I => \N__70504\
        );

    \I__17371\ : ClkMux
    port map (
            O => \N__71014\,
            I => \N__70504\
        );

    \I__17370\ : ClkMux
    port map (
            O => \N__71013\,
            I => \N__70504\
        );

    \I__17369\ : ClkMux
    port map (
            O => \N__71012\,
            I => \N__70504\
        );

    \I__17368\ : ClkMux
    port map (
            O => \N__71011\,
            I => \N__70504\
        );

    \I__17367\ : ClkMux
    port map (
            O => \N__71010\,
            I => \N__70504\
        );

    \I__17366\ : ClkMux
    port map (
            O => \N__71009\,
            I => \N__70504\
        );

    \I__17365\ : ClkMux
    port map (
            O => \N__71008\,
            I => \N__70504\
        );

    \I__17364\ : ClkMux
    port map (
            O => \N__71007\,
            I => \N__70504\
        );

    \I__17363\ : ClkMux
    port map (
            O => \N__71006\,
            I => \N__70504\
        );

    \I__17362\ : ClkMux
    port map (
            O => \N__71005\,
            I => \N__70504\
        );

    \I__17361\ : ClkMux
    port map (
            O => \N__71004\,
            I => \N__70504\
        );

    \I__17360\ : ClkMux
    port map (
            O => \N__71003\,
            I => \N__70504\
        );

    \I__17359\ : ClkMux
    port map (
            O => \N__71002\,
            I => \N__70504\
        );

    \I__17358\ : ClkMux
    port map (
            O => \N__71001\,
            I => \N__70504\
        );

    \I__17357\ : ClkMux
    port map (
            O => \N__71000\,
            I => \N__70504\
        );

    \I__17356\ : ClkMux
    port map (
            O => \N__70999\,
            I => \N__70504\
        );

    \I__17355\ : ClkMux
    port map (
            O => \N__70998\,
            I => \N__70504\
        );

    \I__17354\ : ClkMux
    port map (
            O => \N__70997\,
            I => \N__70504\
        );

    \I__17353\ : ClkMux
    port map (
            O => \N__70996\,
            I => \N__70504\
        );

    \I__17352\ : ClkMux
    port map (
            O => \N__70995\,
            I => \N__70504\
        );

    \I__17351\ : ClkMux
    port map (
            O => \N__70994\,
            I => \N__70504\
        );

    \I__17350\ : ClkMux
    port map (
            O => \N__70993\,
            I => \N__70504\
        );

    \I__17349\ : ClkMux
    port map (
            O => \N__70992\,
            I => \N__70504\
        );

    \I__17348\ : ClkMux
    port map (
            O => \N__70991\,
            I => \N__70504\
        );

    \I__17347\ : GlobalMux
    port map (
            O => \N__70504\,
            I => \N__70501\
        );

    \I__17346\ : gio2CtrlBuf
    port map (
            O => \N__70501\,
            I => \CLK_c\
        );

    \I__17345\ : CascadeMux
    port map (
            O => \N__70498\,
            I => \N__70495\
        );

    \I__17344\ : InMux
    port map (
            O => \N__70495\,
            I => \N__70491\
        );

    \I__17343\ : InMux
    port map (
            O => \N__70494\,
            I => \N__70488\
        );

    \I__17342\ : LocalMux
    port map (
            O => \N__70491\,
            I => \N__70485\
        );

    \I__17341\ : LocalMux
    port map (
            O => \N__70488\,
            I => \N__70482\
        );

    \I__17340\ : Span4Mux_v
    port map (
            O => \N__70485\,
            I => \N__70478\
        );

    \I__17339\ : Span4Mux_h
    port map (
            O => \N__70482\,
            I => \N__70475\
        );

    \I__17338\ : InMux
    port map (
            O => \N__70481\,
            I => \N__70472\
        );

    \I__17337\ : Odrv4
    port map (
            O => \N__70478\,
            I => \c0.n19162\
        );

    \I__17336\ : Odrv4
    port map (
            O => \N__70475\,
            I => \c0.n19162\
        );

    \I__17335\ : LocalMux
    port map (
            O => \N__70472\,
            I => \c0.n19162\
        );

    \I__17334\ : CascadeMux
    port map (
            O => \N__70465\,
            I => \N__70461\
        );

    \I__17333\ : InMux
    port map (
            O => \N__70464\,
            I => \N__70457\
        );

    \I__17332\ : InMux
    port map (
            O => \N__70461\,
            I => \N__70451\
        );

    \I__17331\ : InMux
    port map (
            O => \N__70460\,
            I => \N__70451\
        );

    \I__17330\ : LocalMux
    port map (
            O => \N__70457\,
            I => \N__70448\
        );

    \I__17329\ : InMux
    port map (
            O => \N__70456\,
            I => \N__70445\
        );

    \I__17328\ : LocalMux
    port map (
            O => \N__70451\,
            I => \N__70442\
        );

    \I__17327\ : Span4Mux_v
    port map (
            O => \N__70448\,
            I => \N__70439\
        );

    \I__17326\ : LocalMux
    port map (
            O => \N__70445\,
            I => \N__70435\
        );

    \I__17325\ : Span4Mux_v
    port map (
            O => \N__70442\,
            I => \N__70432\
        );

    \I__17324\ : Span4Mux_h
    port map (
            O => \N__70439\,
            I => \N__70429\
        );

    \I__17323\ : InMux
    port map (
            O => \N__70438\,
            I => \N__70425\
        );

    \I__17322\ : Span4Mux_v
    port map (
            O => \N__70435\,
            I => \N__70420\
        );

    \I__17321\ : Span4Mux_h
    port map (
            O => \N__70432\,
            I => \N__70420\
        );

    \I__17320\ : Span4Mux_h
    port map (
            O => \N__70429\,
            I => \N__70417\
        );

    \I__17319\ : InMux
    port map (
            O => \N__70428\,
            I => \N__70414\
        );

    \I__17318\ : LocalMux
    port map (
            O => \N__70425\,
            I => data_in_frame_22_1
        );

    \I__17317\ : Odrv4
    port map (
            O => \N__70420\,
            I => data_in_frame_22_1
        );

    \I__17316\ : Odrv4
    port map (
            O => \N__70417\,
            I => data_in_frame_22_1
        );

    \I__17315\ : LocalMux
    port map (
            O => \N__70414\,
            I => data_in_frame_22_1
        );

    \I__17314\ : InMux
    port map (
            O => \N__70405\,
            I => \N__70402\
        );

    \I__17313\ : LocalMux
    port map (
            O => \N__70402\,
            I => \N__70399\
        );

    \I__17312\ : Span4Mux_v
    port map (
            O => \N__70399\,
            I => \N__70396\
        );

    \I__17311\ : Span4Mux_h
    port map (
            O => \N__70396\,
            I => \N__70393\
        );

    \I__17310\ : Odrv4
    port map (
            O => \N__70393\,
            I => \c0.n20332\
        );

    \I__17309\ : InMux
    port map (
            O => \N__70390\,
            I => \N__70386\
        );

    \I__17308\ : InMux
    port map (
            O => \N__70389\,
            I => \N__70383\
        );

    \I__17307\ : LocalMux
    port map (
            O => \N__70386\,
            I => \N__70379\
        );

    \I__17306\ : LocalMux
    port map (
            O => \N__70383\,
            I => \N__70376\
        );

    \I__17305\ : InMux
    port map (
            O => \N__70382\,
            I => \N__70371\
        );

    \I__17304\ : Span4Mux_v
    port map (
            O => \N__70379\,
            I => \N__70368\
        );

    \I__17303\ : Span4Mux_h
    port map (
            O => \N__70376\,
            I => \N__70365\
        );

    \I__17302\ : InMux
    port map (
            O => \N__70375\,
            I => \N__70362\
        );

    \I__17301\ : InMux
    port map (
            O => \N__70374\,
            I => \N__70359\
        );

    \I__17300\ : LocalMux
    port map (
            O => \N__70371\,
            I => \N__70354\
        );

    \I__17299\ : Span4Mux_v
    port map (
            O => \N__70368\,
            I => \N__70354\
        );

    \I__17298\ : Span4Mux_h
    port map (
            O => \N__70365\,
            I => \N__70351\
        );

    \I__17297\ : LocalMux
    port map (
            O => \N__70362\,
            I => \N__70348\
        );

    \I__17296\ : LocalMux
    port map (
            O => \N__70359\,
            I => data_in_frame_24_1
        );

    \I__17295\ : Odrv4
    port map (
            O => \N__70354\,
            I => data_in_frame_24_1
        );

    \I__17294\ : Odrv4
    port map (
            O => \N__70351\,
            I => data_in_frame_24_1
        );

    \I__17293\ : Odrv4
    port map (
            O => \N__70348\,
            I => data_in_frame_24_1
        );

    \I__17292\ : InMux
    port map (
            O => \N__70339\,
            I => \N__70334\
        );

    \I__17291\ : CascadeMux
    port map (
            O => \N__70338\,
            I => \N__70331\
        );

    \I__17290\ : InMux
    port map (
            O => \N__70337\,
            I => \N__70328\
        );

    \I__17289\ : LocalMux
    port map (
            O => \N__70334\,
            I => \N__70325\
        );

    \I__17288\ : InMux
    port map (
            O => \N__70331\,
            I => \N__70321\
        );

    \I__17287\ : LocalMux
    port map (
            O => \N__70328\,
            I => \N__70318\
        );

    \I__17286\ : Span4Mux_h
    port map (
            O => \N__70325\,
            I => \N__70315\
        );

    \I__17285\ : InMux
    port map (
            O => \N__70324\,
            I => \N__70311\
        );

    \I__17284\ : LocalMux
    port map (
            O => \N__70321\,
            I => \N__70308\
        );

    \I__17283\ : Span4Mux_v
    port map (
            O => \N__70318\,
            I => \N__70303\
        );

    \I__17282\ : Span4Mux_v
    port map (
            O => \N__70315\,
            I => \N__70303\
        );

    \I__17281\ : InMux
    port map (
            O => \N__70314\,
            I => \N__70300\
        );

    \I__17280\ : LocalMux
    port map (
            O => \N__70311\,
            I => data_in_frame_24_3
        );

    \I__17279\ : Odrv12
    port map (
            O => \N__70308\,
            I => data_in_frame_24_3
        );

    \I__17278\ : Odrv4
    port map (
            O => \N__70303\,
            I => data_in_frame_24_3
        );

    \I__17277\ : LocalMux
    port map (
            O => \N__70300\,
            I => data_in_frame_24_3
        );

    \I__17276\ : CascadeMux
    port map (
            O => \N__70291\,
            I => \c0.n20332_cascade_\
        );

    \I__17275\ : InMux
    port map (
            O => \N__70288\,
            I => \N__70285\
        );

    \I__17274\ : LocalMux
    port map (
            O => \N__70285\,
            I => \N__70282\
        );

    \I__17273\ : Odrv4
    port map (
            O => \N__70282\,
            I => \c0.n18413\
        );

    \I__17272\ : InMux
    port map (
            O => \N__70279\,
            I => \N__70276\
        );

    \I__17271\ : LocalMux
    port map (
            O => \N__70276\,
            I => \N__70273\
        );

    \I__17270\ : Span4Mux_v
    port map (
            O => \N__70273\,
            I => \N__70270\
        );

    \I__17269\ : Span4Mux_h
    port map (
            O => \N__70270\,
            I => \N__70267\
        );

    \I__17268\ : Odrv4
    port map (
            O => \N__70267\,
            I => \c0.n36\
        );

    \I__17267\ : InMux
    port map (
            O => \N__70264\,
            I => \N__70261\
        );

    \I__17266\ : LocalMux
    port map (
            O => \N__70261\,
            I => \N__70258\
        );

    \I__17265\ : Span4Mux_h
    port map (
            O => \N__70258\,
            I => \N__70254\
        );

    \I__17264\ : InMux
    port map (
            O => \N__70257\,
            I => \N__70251\
        );

    \I__17263\ : Span4Mux_v
    port map (
            O => \N__70254\,
            I => \N__70248\
        );

    \I__17262\ : LocalMux
    port map (
            O => \N__70251\,
            I => \c0.n20642\
        );

    \I__17261\ : Odrv4
    port map (
            O => \N__70248\,
            I => \c0.n20642\
        );

    \I__17260\ : InMux
    port map (
            O => \N__70243\,
            I => \N__70239\
        );

    \I__17259\ : InMux
    port map (
            O => \N__70242\,
            I => \N__70236\
        );

    \I__17258\ : LocalMux
    port map (
            O => \N__70239\,
            I => \N__70233\
        );

    \I__17257\ : LocalMux
    port map (
            O => \N__70236\,
            I => \N__70230\
        );

    \I__17256\ : Odrv4
    port map (
            O => \N__70233\,
            I => \c0.n18525\
        );

    \I__17255\ : Odrv4
    port map (
            O => \N__70230\,
            I => \c0.n18525\
        );

    \I__17254\ : CascadeMux
    port map (
            O => \N__70225\,
            I => \N__70221\
        );

    \I__17253\ : CascadeMux
    port map (
            O => \N__70224\,
            I => \N__70218\
        );

    \I__17252\ : InMux
    port map (
            O => \N__70221\,
            I => \N__70213\
        );

    \I__17251\ : InMux
    port map (
            O => \N__70218\,
            I => \N__70213\
        );

    \I__17250\ : LocalMux
    port map (
            O => \N__70213\,
            I => \N__70210\
        );

    \I__17249\ : Span4Mux_h
    port map (
            O => \N__70210\,
            I => \N__70205\
        );

    \I__17248\ : InMux
    port map (
            O => \N__70209\,
            I => \N__70202\
        );

    \I__17247\ : InMux
    port map (
            O => \N__70208\,
            I => \N__70199\
        );

    \I__17246\ : Span4Mux_h
    port map (
            O => \N__70205\,
            I => \N__70196\
        );

    \I__17245\ : LocalMux
    port map (
            O => \N__70202\,
            I => data_in_frame_24_2
        );

    \I__17244\ : LocalMux
    port map (
            O => \N__70199\,
            I => data_in_frame_24_2
        );

    \I__17243\ : Odrv4
    port map (
            O => \N__70196\,
            I => data_in_frame_24_2
        );

    \I__17242\ : InMux
    port map (
            O => \N__70189\,
            I => \N__70183\
        );

    \I__17241\ : InMux
    port map (
            O => \N__70188\,
            I => \N__70183\
        );

    \I__17240\ : LocalMux
    port map (
            O => \N__70183\,
            I => \c0.n18498\
        );

    \I__17239\ : InMux
    port map (
            O => \N__70180\,
            I => \N__70177\
        );

    \I__17238\ : LocalMux
    port map (
            O => \N__70177\,
            I => \N__70174\
        );

    \I__17237\ : Span4Mux_h
    port map (
            O => \N__70174\,
            I => \N__70171\
        );

    \I__17236\ : Span4Mux_h
    port map (
            O => \N__70171\,
            I => \N__70168\
        );

    \I__17235\ : Odrv4
    port map (
            O => \N__70168\,
            I => \c0.n10_adj_3410\
        );

    \I__17234\ : CascadeMux
    port map (
            O => \N__70165\,
            I => \N__70162\
        );

    \I__17233\ : InMux
    port map (
            O => \N__70162\,
            I => \N__70158\
        );

    \I__17232\ : InMux
    port map (
            O => \N__70161\,
            I => \N__70155\
        );

    \I__17231\ : LocalMux
    port map (
            O => \N__70158\,
            I => \N__70151\
        );

    \I__17230\ : LocalMux
    port map (
            O => \N__70155\,
            I => \N__70148\
        );

    \I__17229\ : CascadeMux
    port map (
            O => \N__70154\,
            I => \N__70144\
        );

    \I__17228\ : Span4Mux_v
    port map (
            O => \N__70151\,
            I => \N__70139\
        );

    \I__17227\ : Span4Mux_v
    port map (
            O => \N__70148\,
            I => \N__70139\
        );

    \I__17226\ : InMux
    port map (
            O => \N__70147\,
            I => \N__70134\
        );

    \I__17225\ : InMux
    port map (
            O => \N__70144\,
            I => \N__70134\
        );

    \I__17224\ : Span4Mux_h
    port map (
            O => \N__70139\,
            I => \N__70131\
        );

    \I__17223\ : LocalMux
    port map (
            O => \N__70134\,
            I => \c0.data_in_frame_20_7\
        );

    \I__17222\ : Odrv4
    port map (
            O => \N__70131\,
            I => \c0.data_in_frame_20_7\
        );

    \I__17221\ : InMux
    port map (
            O => \N__70126\,
            I => \N__70120\
        );

    \I__17220\ : CascadeMux
    port map (
            O => \N__70125\,
            I => \N__70117\
        );

    \I__17219\ : InMux
    port map (
            O => \N__70124\,
            I => \N__70114\
        );

    \I__17218\ : InMux
    port map (
            O => \N__70123\,
            I => \N__70111\
        );

    \I__17217\ : LocalMux
    port map (
            O => \N__70120\,
            I => \N__70108\
        );

    \I__17216\ : InMux
    port map (
            O => \N__70117\,
            I => \N__70105\
        );

    \I__17215\ : LocalMux
    port map (
            O => \N__70114\,
            I => \N__70102\
        );

    \I__17214\ : LocalMux
    port map (
            O => \N__70111\,
            I => \N__70099\
        );

    \I__17213\ : Span12Mux_h
    port map (
            O => \N__70108\,
            I => \N__70096\
        );

    \I__17212\ : LocalMux
    port map (
            O => \N__70105\,
            I => \N__70091\
        );

    \I__17211\ : Span12Mux_v
    port map (
            O => \N__70102\,
            I => \N__70091\
        );

    \I__17210\ : Odrv4
    port map (
            O => \N__70099\,
            I => \c0.data_in_frame_20_6\
        );

    \I__17209\ : Odrv12
    port map (
            O => \N__70096\,
            I => \c0.data_in_frame_20_6\
        );

    \I__17208\ : Odrv12
    port map (
            O => \N__70091\,
            I => \c0.data_in_frame_20_6\
        );

    \I__17207\ : InMux
    port map (
            O => \N__70084\,
            I => \N__70080\
        );

    \I__17206\ : InMux
    port map (
            O => \N__70083\,
            I => \N__70077\
        );

    \I__17205\ : LocalMux
    port map (
            O => \N__70080\,
            I => \N__70074\
        );

    \I__17204\ : LocalMux
    port map (
            O => \N__70077\,
            I => \c0.n20576\
        );

    \I__17203\ : Odrv12
    port map (
            O => \N__70074\,
            I => \c0.n20576\
        );

    \I__17202\ : InMux
    port map (
            O => \N__70069\,
            I => \N__70066\
        );

    \I__17201\ : LocalMux
    port map (
            O => \N__70066\,
            I => \c0.n12_adj_3439\
        );

    \I__17200\ : InMux
    port map (
            O => \N__70063\,
            I => \N__70060\
        );

    \I__17199\ : LocalMux
    port map (
            O => \N__70060\,
            I => \N__70057\
        );

    \I__17198\ : Span4Mux_v
    port map (
            O => \N__70057\,
            I => \N__70053\
        );

    \I__17197\ : InMux
    port map (
            O => \N__70056\,
            I => \N__70050\
        );

    \I__17196\ : Span4Mux_h
    port map (
            O => \N__70053\,
            I => \N__70045\
        );

    \I__17195\ : LocalMux
    port map (
            O => \N__70050\,
            I => \N__70045\
        );

    \I__17194\ : Span4Mux_v
    port map (
            O => \N__70045\,
            I => \N__70041\
        );

    \I__17193\ : InMux
    port map (
            O => \N__70044\,
            I => \N__70038\
        );

    \I__17192\ : Sp12to4
    port map (
            O => \N__70041\,
            I => \N__70032\
        );

    \I__17191\ : LocalMux
    port map (
            O => \N__70038\,
            I => \N__70032\
        );

    \I__17190\ : InMux
    port map (
            O => \N__70037\,
            I => \N__70029\
        );

    \I__17189\ : Span12Mux_h
    port map (
            O => \N__70032\,
            I => \N__70026\
        );

    \I__17188\ : LocalMux
    port map (
            O => \N__70029\,
            I => data_in_frame_22_0
        );

    \I__17187\ : Odrv12
    port map (
            O => \N__70026\,
            I => data_in_frame_22_0
        );

    \I__17186\ : InMux
    port map (
            O => \N__70021\,
            I => \N__70018\
        );

    \I__17185\ : LocalMux
    port map (
            O => \N__70018\,
            I => \N__70013\
        );

    \I__17184\ : InMux
    port map (
            O => \N__70017\,
            I => \N__70010\
        );

    \I__17183\ : InMux
    port map (
            O => \N__70016\,
            I => \N__70007\
        );

    \I__17182\ : Span4Mux_h
    port map (
            O => \N__70013\,
            I => \N__70004\
        );

    \I__17181\ : LocalMux
    port map (
            O => \N__70010\,
            I => \N__70001\
        );

    \I__17180\ : LocalMux
    port map (
            O => \N__70007\,
            I => \N__69998\
        );

    \I__17179\ : Odrv4
    port map (
            O => \N__70004\,
            I => \c0.n18415\
        );

    \I__17178\ : Odrv4
    port map (
            O => \N__70001\,
            I => \c0.n18415\
        );

    \I__17177\ : Odrv4
    port map (
            O => \N__69998\,
            I => \c0.n18415\
        );

    \I__17176\ : CascadeMux
    port map (
            O => \N__69991\,
            I => \c0.n4_adj_3067_cascade_\
        );

    \I__17175\ : InMux
    port map (
            O => \N__69988\,
            I => \N__69983\
        );

    \I__17174\ : InMux
    port map (
            O => \N__69987\,
            I => \N__69980\
        );

    \I__17173\ : InMux
    port map (
            O => \N__69986\,
            I => \N__69977\
        );

    \I__17172\ : LocalMux
    port map (
            O => \N__69983\,
            I => \N__69974\
        );

    \I__17171\ : LocalMux
    port map (
            O => \N__69980\,
            I => \N__69971\
        );

    \I__17170\ : LocalMux
    port map (
            O => \N__69977\,
            I => \N__69968\
        );

    \I__17169\ : Span4Mux_v
    port map (
            O => \N__69974\,
            I => \N__69961\
        );

    \I__17168\ : Span4Mux_h
    port map (
            O => \N__69971\,
            I => \N__69958\
        );

    \I__17167\ : Span4Mux_h
    port map (
            O => \N__69968\,
            I => \N__69955\
        );

    \I__17166\ : InMux
    port map (
            O => \N__69967\,
            I => \N__69946\
        );

    \I__17165\ : InMux
    port map (
            O => \N__69966\,
            I => \N__69946\
        );

    \I__17164\ : InMux
    port map (
            O => \N__69965\,
            I => \N__69946\
        );

    \I__17163\ : InMux
    port map (
            O => \N__69964\,
            I => \N__69946\
        );

    \I__17162\ : Odrv4
    port map (
            O => \N__69961\,
            I => \c0.n6009\
        );

    \I__17161\ : Odrv4
    port map (
            O => \N__69958\,
            I => \c0.n6009\
        );

    \I__17160\ : Odrv4
    port map (
            O => \N__69955\,
            I => \c0.n6009\
        );

    \I__17159\ : LocalMux
    port map (
            O => \N__69946\,
            I => \c0.n6009\
        );

    \I__17158\ : InMux
    port map (
            O => \N__69937\,
            I => \N__69934\
        );

    \I__17157\ : LocalMux
    port map (
            O => \N__69934\,
            I => \N__69930\
        );

    \I__17156\ : InMux
    port map (
            O => \N__69933\,
            I => \N__69927\
        );

    \I__17155\ : Odrv12
    port map (
            O => \N__69930\,
            I => \c0.n19369\
        );

    \I__17154\ : LocalMux
    port map (
            O => \N__69927\,
            I => \c0.n19369\
        );

    \I__17153\ : CascadeMux
    port map (
            O => \N__69922\,
            I => \c0.n22_adj_3322_cascade_\
        );

    \I__17152\ : InMux
    port map (
            O => \N__69919\,
            I => \N__69913\
        );

    \I__17151\ : InMux
    port map (
            O => \N__69918\,
            I => \N__69913\
        );

    \I__17150\ : LocalMux
    port map (
            O => \N__69913\,
            I => \N__69910\
        );

    \I__17149\ : Odrv4
    port map (
            O => \N__69910\,
            I => \c0.n36_adj_3090\
        );

    \I__17148\ : CascadeMux
    port map (
            O => \N__69907\,
            I => \N__69904\
        );

    \I__17147\ : InMux
    port map (
            O => \N__69904\,
            I => \N__69900\
        );

    \I__17146\ : InMux
    port map (
            O => \N__69903\,
            I => \N__69897\
        );

    \I__17145\ : LocalMux
    port map (
            O => \N__69900\,
            I => \N__69893\
        );

    \I__17144\ : LocalMux
    port map (
            O => \N__69897\,
            I => \N__69890\
        );

    \I__17143\ : CascadeMux
    port map (
            O => \N__69896\,
            I => \N__69886\
        );

    \I__17142\ : Span4Mux_h
    port map (
            O => \N__69893\,
            I => \N__69883\
        );

    \I__17141\ : Span4Mux_v
    port map (
            O => \N__69890\,
            I => \N__69880\
        );

    \I__17140\ : CascadeMux
    port map (
            O => \N__69889\,
            I => \N__69876\
        );

    \I__17139\ : InMux
    port map (
            O => \N__69886\,
            I => \N__69873\
        );

    \I__17138\ : Span4Mux_h
    port map (
            O => \N__69883\,
            I => \N__69870\
        );

    \I__17137\ : Sp12to4
    port map (
            O => \N__69880\,
            I => \N__69867\
        );

    \I__17136\ : InMux
    port map (
            O => \N__69879\,
            I => \N__69862\
        );

    \I__17135\ : InMux
    port map (
            O => \N__69876\,
            I => \N__69862\
        );

    \I__17134\ : LocalMux
    port map (
            O => \N__69873\,
            I => \c0.data_in_frame_21_2\
        );

    \I__17133\ : Odrv4
    port map (
            O => \N__69870\,
            I => \c0.data_in_frame_21_2\
        );

    \I__17132\ : Odrv12
    port map (
            O => \N__69867\,
            I => \c0.data_in_frame_21_2\
        );

    \I__17131\ : LocalMux
    port map (
            O => \N__69862\,
            I => \c0.data_in_frame_21_2\
        );

    \I__17130\ : InMux
    port map (
            O => \N__69853\,
            I => \N__69850\
        );

    \I__17129\ : LocalMux
    port map (
            O => \N__69850\,
            I => \N__69845\
        );

    \I__17128\ : InMux
    port map (
            O => \N__69849\,
            I => \N__69840\
        );

    \I__17127\ : InMux
    port map (
            O => \N__69848\,
            I => \N__69840\
        );

    \I__17126\ : Odrv4
    port map (
            O => \N__69845\,
            I => \c0.n29_adj_3383\
        );

    \I__17125\ : LocalMux
    port map (
            O => \N__69840\,
            I => \c0.n29_adj_3383\
        );

    \I__17124\ : InMux
    port map (
            O => \N__69835\,
            I => \N__69831\
        );

    \I__17123\ : InMux
    port map (
            O => \N__69834\,
            I => \N__69828\
        );

    \I__17122\ : LocalMux
    port map (
            O => \N__69831\,
            I => \N__69822\
        );

    \I__17121\ : LocalMux
    port map (
            O => \N__69828\,
            I => \N__69819\
        );

    \I__17120\ : InMux
    port map (
            O => \N__69827\,
            I => \N__69812\
        );

    \I__17119\ : InMux
    port map (
            O => \N__69826\,
            I => \N__69812\
        );

    \I__17118\ : InMux
    port map (
            O => \N__69825\,
            I => \N__69809\
        );

    \I__17117\ : Span4Mux_h
    port map (
            O => \N__69822\,
            I => \N__69804\
        );

    \I__17116\ : Span4Mux_h
    port map (
            O => \N__69819\,
            I => \N__69804\
        );

    \I__17115\ : InMux
    port map (
            O => \N__69818\,
            I => \N__69801\
        );

    \I__17114\ : InMux
    port map (
            O => \N__69817\,
            I => \N__69798\
        );

    \I__17113\ : LocalMux
    port map (
            O => \N__69812\,
            I => \c0.n20917\
        );

    \I__17112\ : LocalMux
    port map (
            O => \N__69809\,
            I => \c0.n20917\
        );

    \I__17111\ : Odrv4
    port map (
            O => \N__69804\,
            I => \c0.n20917\
        );

    \I__17110\ : LocalMux
    port map (
            O => \N__69801\,
            I => \c0.n20917\
        );

    \I__17109\ : LocalMux
    port map (
            O => \N__69798\,
            I => \c0.n20917\
        );

    \I__17108\ : InMux
    port map (
            O => \N__69787\,
            I => \N__69784\
        );

    \I__17107\ : LocalMux
    port map (
            O => \N__69784\,
            I => \N__69781\
        );

    \I__17106\ : Span4Mux_h
    port map (
            O => \N__69781\,
            I => \N__69778\
        );

    \I__17105\ : Span4Mux_v
    port map (
            O => \N__69778\,
            I => \N__69774\
        );

    \I__17104\ : CascadeMux
    port map (
            O => \N__69777\,
            I => \N__69769\
        );

    \I__17103\ : Sp12to4
    port map (
            O => \N__69774\,
            I => \N__69766\
        );

    \I__17102\ : InMux
    port map (
            O => \N__69773\,
            I => \N__69761\
        );

    \I__17101\ : InMux
    port map (
            O => \N__69772\,
            I => \N__69761\
        );

    \I__17100\ : InMux
    port map (
            O => \N__69769\,
            I => \N__69758\
        );

    \I__17099\ : Span12Mux_s8_h
    port map (
            O => \N__69766\,
            I => \N__69753\
        );

    \I__17098\ : LocalMux
    port map (
            O => \N__69761\,
            I => \N__69753\
        );

    \I__17097\ : LocalMux
    port map (
            O => \N__69758\,
            I => \c0.data_in_frame_20_0\
        );

    \I__17096\ : Odrv12
    port map (
            O => \N__69753\,
            I => \c0.data_in_frame_20_0\
        );

    \I__17095\ : InMux
    port map (
            O => \N__69748\,
            I => \N__69739\
        );

    \I__17094\ : InMux
    port map (
            O => \N__69747\,
            I => \N__69739\
        );

    \I__17093\ : InMux
    port map (
            O => \N__69746\,
            I => \N__69734\
        );

    \I__17092\ : InMux
    port map (
            O => \N__69745\,
            I => \N__69734\
        );

    \I__17091\ : InMux
    port map (
            O => \N__69744\,
            I => \N__69731\
        );

    \I__17090\ : LocalMux
    port map (
            O => \N__69739\,
            I => \N__69726\
        );

    \I__17089\ : LocalMux
    port map (
            O => \N__69734\,
            I => \N__69726\
        );

    \I__17088\ : LocalMux
    port map (
            O => \N__69731\,
            I => \N__69723\
        );

    \I__17087\ : Span4Mux_v
    port map (
            O => \N__69726\,
            I => \N__69718\
        );

    \I__17086\ : Span4Mux_v
    port map (
            O => \N__69723\,
            I => \N__69718\
        );

    \I__17085\ : Odrv4
    port map (
            O => \N__69718\,
            I => \c0.n4_adj_3435\
        );

    \I__17084\ : CascadeMux
    port map (
            O => \N__69715\,
            I => \N__69711\
        );

    \I__17083\ : InMux
    port map (
            O => \N__69714\,
            I => \N__69708\
        );

    \I__17082\ : InMux
    port map (
            O => \N__69711\,
            I => \N__69704\
        );

    \I__17081\ : LocalMux
    port map (
            O => \N__69708\,
            I => \N__69701\
        );

    \I__17080\ : InMux
    port map (
            O => \N__69707\,
            I => \N__69698\
        );

    \I__17079\ : LocalMux
    port map (
            O => \N__69704\,
            I => \N__69695\
        );

    \I__17078\ : Odrv4
    port map (
            O => \N__69701\,
            I => \c0.n6_adj_3091\
        );

    \I__17077\ : LocalMux
    port map (
            O => \N__69698\,
            I => \c0.n6_adj_3091\
        );

    \I__17076\ : Odrv12
    port map (
            O => \N__69695\,
            I => \c0.n6_adj_3091\
        );

    \I__17075\ : InMux
    port map (
            O => \N__69688\,
            I => \N__69685\
        );

    \I__17074\ : LocalMux
    port map (
            O => \N__69685\,
            I => \N__69679\
        );

    \I__17073\ : InMux
    port map (
            O => \N__69684\,
            I => \N__69676\
        );

    \I__17072\ : InMux
    port map (
            O => \N__69683\,
            I => \N__69673\
        );

    \I__17071\ : InMux
    port map (
            O => \N__69682\,
            I => \N__69670\
        );

    \I__17070\ : Odrv12
    port map (
            O => \N__69679\,
            I => \c0.n18375\
        );

    \I__17069\ : LocalMux
    port map (
            O => \N__69676\,
            I => \c0.n18375\
        );

    \I__17068\ : LocalMux
    port map (
            O => \N__69673\,
            I => \c0.n18375\
        );

    \I__17067\ : LocalMux
    port map (
            O => \N__69670\,
            I => \c0.n18375\
        );

    \I__17066\ : CascadeMux
    port map (
            O => \N__69661\,
            I => \c0.n6_adj_3091_cascade_\
        );

    \I__17065\ : InMux
    port map (
            O => \N__69658\,
            I => \N__69653\
        );

    \I__17064\ : CascadeMux
    port map (
            O => \N__69657\,
            I => \N__69649\
        );

    \I__17063\ : InMux
    port map (
            O => \N__69656\,
            I => \N__69645\
        );

    \I__17062\ : LocalMux
    port map (
            O => \N__69653\,
            I => \N__69642\
        );

    \I__17061\ : InMux
    port map (
            O => \N__69652\,
            I => \N__69637\
        );

    \I__17060\ : InMux
    port map (
            O => \N__69649\,
            I => \N__69637\
        );

    \I__17059\ : InMux
    port map (
            O => \N__69648\,
            I => \N__69633\
        );

    \I__17058\ : LocalMux
    port map (
            O => \N__69645\,
            I => \N__69630\
        );

    \I__17057\ : Span4Mux_v
    port map (
            O => \N__69642\,
            I => \N__69625\
        );

    \I__17056\ : LocalMux
    port map (
            O => \N__69637\,
            I => \N__69625\
        );

    \I__17055\ : InMux
    port map (
            O => \N__69636\,
            I => \N__69622\
        );

    \I__17054\ : LocalMux
    port map (
            O => \N__69633\,
            I => \N__69619\
        );

    \I__17053\ : Span4Mux_h
    port map (
            O => \N__69630\,
            I => \N__69614\
        );

    \I__17052\ : Span4Mux_h
    port map (
            O => \N__69625\,
            I => \N__69614\
        );

    \I__17051\ : LocalMux
    port map (
            O => \N__69622\,
            I => \c0.n17900\
        );

    \I__17050\ : Odrv12
    port map (
            O => \N__69619\,
            I => \c0.n17900\
        );

    \I__17049\ : Odrv4
    port map (
            O => \N__69614\,
            I => \c0.n17900\
        );

    \I__17048\ : CascadeMux
    port map (
            O => \N__69607\,
            I => \N__69603\
        );

    \I__17047\ : CascadeMux
    port map (
            O => \N__69606\,
            I => \N__69599\
        );

    \I__17046\ : InMux
    port map (
            O => \N__69603\,
            I => \N__69596\
        );

    \I__17045\ : CascadeMux
    port map (
            O => \N__69602\,
            I => \N__69592\
        );

    \I__17044\ : InMux
    port map (
            O => \N__69599\,
            I => \N__69589\
        );

    \I__17043\ : LocalMux
    port map (
            O => \N__69596\,
            I => \N__69586\
        );

    \I__17042\ : InMux
    port map (
            O => \N__69595\,
            I => \N__69583\
        );

    \I__17041\ : InMux
    port map (
            O => \N__69592\,
            I => \N__69580\
        );

    \I__17040\ : LocalMux
    port map (
            O => \N__69589\,
            I => \N__69577\
        );

    \I__17039\ : Span4Mux_h
    port map (
            O => \N__69586\,
            I => \N__69572\
        );

    \I__17038\ : LocalMux
    port map (
            O => \N__69583\,
            I => \N__69572\
        );

    \I__17037\ : LocalMux
    port map (
            O => \N__69580\,
            I => \c0.data_in_frame_21_3\
        );

    \I__17036\ : Odrv4
    port map (
            O => \N__69577\,
            I => \c0.data_in_frame_21_3\
        );

    \I__17035\ : Odrv4
    port map (
            O => \N__69572\,
            I => \c0.data_in_frame_21_3\
        );

    \I__17034\ : InMux
    port map (
            O => \N__69565\,
            I => \N__69561\
        );

    \I__17033\ : CascadeMux
    port map (
            O => \N__69564\,
            I => \N__69558\
        );

    \I__17032\ : LocalMux
    port map (
            O => \N__69561\,
            I => \N__69552\
        );

    \I__17031\ : InMux
    port map (
            O => \N__69558\,
            I => \N__69547\
        );

    \I__17030\ : InMux
    port map (
            O => \N__69557\,
            I => \N__69547\
        );

    \I__17029\ : CascadeMux
    port map (
            O => \N__69556\,
            I => \N__69544\
        );

    \I__17028\ : CascadeMux
    port map (
            O => \N__69555\,
            I => \N__69540\
        );

    \I__17027\ : Span4Mux_v
    port map (
            O => \N__69552\,
            I => \N__69537\
        );

    \I__17026\ : LocalMux
    port map (
            O => \N__69547\,
            I => \N__69534\
        );

    \I__17025\ : InMux
    port map (
            O => \N__69544\,
            I => \N__69529\
        );

    \I__17024\ : InMux
    port map (
            O => \N__69543\,
            I => \N__69529\
        );

    \I__17023\ : InMux
    port map (
            O => \N__69540\,
            I => \N__69526\
        );

    \I__17022\ : Odrv4
    port map (
            O => \N__69537\,
            I => \c0.data_in_frame_21_5\
        );

    \I__17021\ : Odrv4
    port map (
            O => \N__69534\,
            I => \c0.data_in_frame_21_5\
        );

    \I__17020\ : LocalMux
    port map (
            O => \N__69529\,
            I => \c0.data_in_frame_21_5\
        );

    \I__17019\ : LocalMux
    port map (
            O => \N__69526\,
            I => \c0.data_in_frame_21_5\
        );

    \I__17018\ : InMux
    port map (
            O => \N__69517\,
            I => \N__69514\
        );

    \I__17017\ : LocalMux
    port map (
            O => \N__69514\,
            I => \N__69511\
        );

    \I__17016\ : Span4Mux_h
    port map (
            O => \N__69511\,
            I => \N__69506\
        );

    \I__17015\ : InMux
    port map (
            O => \N__69510\,
            I => \N__69501\
        );

    \I__17014\ : InMux
    port map (
            O => \N__69509\,
            I => \N__69501\
        );

    \I__17013\ : Odrv4
    port map (
            O => \N__69506\,
            I => \c0.n19321\
        );

    \I__17012\ : LocalMux
    port map (
            O => \N__69501\,
            I => \c0.n19321\
        );

    \I__17011\ : InMux
    port map (
            O => \N__69496\,
            I => \N__69493\
        );

    \I__17010\ : LocalMux
    port map (
            O => \N__69493\,
            I => \N__69489\
        );

    \I__17009\ : InMux
    port map (
            O => \N__69492\,
            I => \N__69486\
        );

    \I__17008\ : Span4Mux_h
    port map (
            O => \N__69489\,
            I => \N__69483\
        );

    \I__17007\ : LocalMux
    port map (
            O => \N__69486\,
            I => \N__69480\
        );

    \I__17006\ : Odrv4
    port map (
            O => \N__69483\,
            I => \c0.n12037\
        );

    \I__17005\ : Odrv12
    port map (
            O => \N__69480\,
            I => \c0.n12037\
        );

    \I__17004\ : CascadeMux
    port map (
            O => \N__69475\,
            I => \N__69472\
        );

    \I__17003\ : InMux
    port map (
            O => \N__69472\,
            I => \N__69469\
        );

    \I__17002\ : LocalMux
    port map (
            O => \N__69469\,
            I => \N__69466\
        );

    \I__17001\ : Span4Mux_h
    port map (
            O => \N__69466\,
            I => \N__69462\
        );

    \I__17000\ : CascadeMux
    port map (
            O => \N__69465\,
            I => \N__69459\
        );

    \I__16999\ : Span4Mux_v
    port map (
            O => \N__69462\,
            I => \N__69455\
        );

    \I__16998\ : InMux
    port map (
            O => \N__69459\,
            I => \N__69450\
        );

    \I__16997\ : InMux
    port map (
            O => \N__69458\,
            I => \N__69450\
        );

    \I__16996\ : Odrv4
    port map (
            O => \N__69455\,
            I => data_in_frame_19_7
        );

    \I__16995\ : LocalMux
    port map (
            O => \N__69450\,
            I => data_in_frame_19_7
        );

    \I__16994\ : InMux
    port map (
            O => \N__69445\,
            I => \N__69439\
        );

    \I__16993\ : CascadeMux
    port map (
            O => \N__69444\,
            I => \N__69432\
        );

    \I__16992\ : InMux
    port map (
            O => \N__69443\,
            I => \N__69429\
        );

    \I__16991\ : InMux
    port map (
            O => \N__69442\,
            I => \N__69426\
        );

    \I__16990\ : LocalMux
    port map (
            O => \N__69439\,
            I => \N__69418\
        );

    \I__16989\ : InMux
    port map (
            O => \N__69438\,
            I => \N__69415\
        );

    \I__16988\ : CascadeMux
    port map (
            O => \N__69437\,
            I => \N__69411\
        );

    \I__16987\ : InMux
    port map (
            O => \N__69436\,
            I => \N__69405\
        );

    \I__16986\ : InMux
    port map (
            O => \N__69435\,
            I => \N__69402\
        );

    \I__16985\ : InMux
    port map (
            O => \N__69432\,
            I => \N__69399\
        );

    \I__16984\ : LocalMux
    port map (
            O => \N__69429\,
            I => \N__69396\
        );

    \I__16983\ : LocalMux
    port map (
            O => \N__69426\,
            I => \N__69393\
        );

    \I__16982\ : InMux
    port map (
            O => \N__69425\,
            I => \N__69390\
        );

    \I__16981\ : InMux
    port map (
            O => \N__69424\,
            I => \N__69385\
        );

    \I__16980\ : InMux
    port map (
            O => \N__69423\,
            I => \N__69385\
        );

    \I__16979\ : InMux
    port map (
            O => \N__69422\,
            I => \N__69382\
        );

    \I__16978\ : InMux
    port map (
            O => \N__69421\,
            I => \N__69377\
        );

    \I__16977\ : Span4Mux_h
    port map (
            O => \N__69418\,
            I => \N__69371\
        );

    \I__16976\ : LocalMux
    port map (
            O => \N__69415\,
            I => \N__69371\
        );

    \I__16975\ : InMux
    port map (
            O => \N__69414\,
            I => \N__69364\
        );

    \I__16974\ : InMux
    port map (
            O => \N__69411\,
            I => \N__69364\
        );

    \I__16973\ : InMux
    port map (
            O => \N__69410\,
            I => \N__69364\
        );

    \I__16972\ : InMux
    port map (
            O => \N__69409\,
            I => \N__69360\
        );

    \I__16971\ : InMux
    port map (
            O => \N__69408\,
            I => \N__69357\
        );

    \I__16970\ : LocalMux
    port map (
            O => \N__69405\,
            I => \N__69352\
        );

    \I__16969\ : LocalMux
    port map (
            O => \N__69402\,
            I => \N__69352\
        );

    \I__16968\ : LocalMux
    port map (
            O => \N__69399\,
            I => \N__69349\
        );

    \I__16967\ : Span4Mux_v
    port map (
            O => \N__69396\,
            I => \N__69342\
        );

    \I__16966\ : Span4Mux_v
    port map (
            O => \N__69393\,
            I => \N__69342\
        );

    \I__16965\ : LocalMux
    port map (
            O => \N__69390\,
            I => \N__69342\
        );

    \I__16964\ : LocalMux
    port map (
            O => \N__69385\,
            I => \N__69339\
        );

    \I__16963\ : LocalMux
    port map (
            O => \N__69382\,
            I => \N__69336\
        );

    \I__16962\ : InMux
    port map (
            O => \N__69381\,
            I => \N__69331\
        );

    \I__16961\ : InMux
    port map (
            O => \N__69380\,
            I => \N__69331\
        );

    \I__16960\ : LocalMux
    port map (
            O => \N__69377\,
            I => \N__69328\
        );

    \I__16959\ : InMux
    port map (
            O => \N__69376\,
            I => \N__69325\
        );

    \I__16958\ : Span4Mux_v
    port map (
            O => \N__69371\,
            I => \N__69320\
        );

    \I__16957\ : LocalMux
    port map (
            O => \N__69364\,
            I => \N__69320\
        );

    \I__16956\ : CascadeMux
    port map (
            O => \N__69363\,
            I => \N__69317\
        );

    \I__16955\ : LocalMux
    port map (
            O => \N__69360\,
            I => \N__69311\
        );

    \I__16954\ : LocalMux
    port map (
            O => \N__69357\,
            I => \N__69308\
        );

    \I__16953\ : Span4Mux_v
    port map (
            O => \N__69352\,
            I => \N__69301\
        );

    \I__16952\ : Span4Mux_h
    port map (
            O => \N__69349\,
            I => \N__69301\
        );

    \I__16951\ : Span4Mux_h
    port map (
            O => \N__69342\,
            I => \N__69301\
        );

    \I__16950\ : Span4Mux_v
    port map (
            O => \N__69339\,
            I => \N__69298\
        );

    \I__16949\ : Span4Mux_h
    port map (
            O => \N__69336\,
            I => \N__69293\
        );

    \I__16948\ : LocalMux
    port map (
            O => \N__69331\,
            I => \N__69293\
        );

    \I__16947\ : Span4Mux_h
    port map (
            O => \N__69328\,
            I => \N__69288\
        );

    \I__16946\ : LocalMux
    port map (
            O => \N__69325\,
            I => \N__69288\
        );

    \I__16945\ : Span4Mux_h
    port map (
            O => \N__69320\,
            I => \N__69284\
        );

    \I__16944\ : InMux
    port map (
            O => \N__69317\,
            I => \N__69279\
        );

    \I__16943\ : InMux
    port map (
            O => \N__69316\,
            I => \N__69279\
        );

    \I__16942\ : InMux
    port map (
            O => \N__69315\,
            I => \N__69274\
        );

    \I__16941\ : InMux
    port map (
            O => \N__69314\,
            I => \N__69271\
        );

    \I__16940\ : Span4Mux_h
    port map (
            O => \N__69311\,
            I => \N__69264\
        );

    \I__16939\ : Span4Mux_v
    port map (
            O => \N__69308\,
            I => \N__69264\
        );

    \I__16938\ : Span4Mux_v
    port map (
            O => \N__69301\,
            I => \N__69264\
        );

    \I__16937\ : Span4Mux_v
    port map (
            O => \N__69298\,
            I => \N__69261\
        );

    \I__16936\ : Span4Mux_h
    port map (
            O => \N__69293\,
            I => \N__69256\
        );

    \I__16935\ : Span4Mux_v
    port map (
            O => \N__69288\,
            I => \N__69256\
        );

    \I__16934\ : InMux
    port map (
            O => \N__69287\,
            I => \N__69253\
        );

    \I__16933\ : Span4Mux_v
    port map (
            O => \N__69284\,
            I => \N__69248\
        );

    \I__16932\ : LocalMux
    port map (
            O => \N__69279\,
            I => \N__69248\
        );

    \I__16931\ : InMux
    port map (
            O => \N__69278\,
            I => \N__69242\
        );

    \I__16930\ : InMux
    port map (
            O => \N__69277\,
            I => \N__69242\
        );

    \I__16929\ : LocalMux
    port map (
            O => \N__69274\,
            I => \N__69239\
        );

    \I__16928\ : LocalMux
    port map (
            O => \N__69271\,
            I => \N__69236\
        );

    \I__16927\ : Span4Mux_v
    port map (
            O => \N__69264\,
            I => \N__69233\
        );

    \I__16926\ : Span4Mux_v
    port map (
            O => \N__69261\,
            I => \N__69228\
        );

    \I__16925\ : Span4Mux_h
    port map (
            O => \N__69256\,
            I => \N__69228\
        );

    \I__16924\ : LocalMux
    port map (
            O => \N__69253\,
            I => \N__69225\
        );

    \I__16923\ : Span4Mux_h
    port map (
            O => \N__69248\,
            I => \N__69222\
        );

    \I__16922\ : InMux
    port map (
            O => \N__69247\,
            I => \N__69219\
        );

    \I__16921\ : LocalMux
    port map (
            O => \N__69242\,
            I => \N__69212\
        );

    \I__16920\ : Span4Mux_h
    port map (
            O => \N__69239\,
            I => \N__69207\
        );

    \I__16919\ : Span4Mux_h
    port map (
            O => \N__69236\,
            I => \N__69207\
        );

    \I__16918\ : Span4Mux_h
    port map (
            O => \N__69233\,
            I => \N__69204\
        );

    \I__16917\ : Span4Mux_v
    port map (
            O => \N__69228\,
            I => \N__69201\
        );

    \I__16916\ : Span4Mux_h
    port map (
            O => \N__69225\,
            I => \N__69194\
        );

    \I__16915\ : Span4Mux_h
    port map (
            O => \N__69222\,
            I => \N__69194\
        );

    \I__16914\ : LocalMux
    port map (
            O => \N__69219\,
            I => \N__69194\
        );

    \I__16913\ : InMux
    port map (
            O => \N__69218\,
            I => \N__69189\
        );

    \I__16912\ : InMux
    port map (
            O => \N__69217\,
            I => \N__69189\
        );

    \I__16911\ : InMux
    port map (
            O => \N__69216\,
            I => \N__69184\
        );

    \I__16910\ : InMux
    port map (
            O => \N__69215\,
            I => \N__69184\
        );

    \I__16909\ : Odrv12
    port map (
            O => \N__69212\,
            I => rx_data_3
        );

    \I__16908\ : Odrv4
    port map (
            O => \N__69207\,
            I => rx_data_3
        );

    \I__16907\ : Odrv4
    port map (
            O => \N__69204\,
            I => rx_data_3
        );

    \I__16906\ : Odrv4
    port map (
            O => \N__69201\,
            I => rx_data_3
        );

    \I__16905\ : Odrv4
    port map (
            O => \N__69194\,
            I => rx_data_3
        );

    \I__16904\ : LocalMux
    port map (
            O => \N__69189\,
            I => rx_data_3
        );

    \I__16903\ : LocalMux
    port map (
            O => \N__69184\,
            I => rx_data_3
        );

    \I__16902\ : InMux
    port map (
            O => \N__69169\,
            I => \N__69164\
        );

    \I__16901\ : InMux
    port map (
            O => \N__69168\,
            I => \N__69161\
        );

    \I__16900\ : InMux
    port map (
            O => \N__69167\,
            I => \N__69158\
        );

    \I__16899\ : LocalMux
    port map (
            O => \N__69164\,
            I => \N__69155\
        );

    \I__16898\ : LocalMux
    port map (
            O => \N__69161\,
            I => \N__69152\
        );

    \I__16897\ : LocalMux
    port map (
            O => \N__69158\,
            I => \N__69147\
        );

    \I__16896\ : Span4Mux_h
    port map (
            O => \N__69155\,
            I => \N__69143\
        );

    \I__16895\ : Span4Mux_v
    port map (
            O => \N__69152\,
            I => \N__69140\
        );

    \I__16894\ : InMux
    port map (
            O => \N__69151\,
            I => \N__69133\
        );

    \I__16893\ : InMux
    port map (
            O => \N__69150\,
            I => \N__69133\
        );

    \I__16892\ : Span4Mux_h
    port map (
            O => \N__69147\,
            I => \N__69130\
        );

    \I__16891\ : InMux
    port map (
            O => \N__69146\,
            I => \N__69127\
        );

    \I__16890\ : Span4Mux_v
    port map (
            O => \N__69143\,
            I => \N__69124\
        );

    \I__16889\ : Sp12to4
    port map (
            O => \N__69140\,
            I => \N__69121\
        );

    \I__16888\ : InMux
    port map (
            O => \N__69139\,
            I => \N__69116\
        );

    \I__16887\ : InMux
    port map (
            O => \N__69138\,
            I => \N__69116\
        );

    \I__16886\ : LocalMux
    port map (
            O => \N__69133\,
            I => \N__69111\
        );

    \I__16885\ : Span4Mux_v
    port map (
            O => \N__69130\,
            I => \N__69111\
        );

    \I__16884\ : LocalMux
    port map (
            O => \N__69127\,
            I => \N__69108\
        );

    \I__16883\ : Span4Mux_v
    port map (
            O => \N__69124\,
            I => \N__69105\
        );

    \I__16882\ : Span12Mux_s10_v
    port map (
            O => \N__69121\,
            I => \N__69102\
        );

    \I__16881\ : LocalMux
    port map (
            O => \N__69116\,
            I => \N__69097\
        );

    \I__16880\ : Span4Mux_h
    port map (
            O => \N__69111\,
            I => \N__69097\
        );

    \I__16879\ : Span4Mux_h
    port map (
            O => \N__69108\,
            I => \N__69092\
        );

    \I__16878\ : Span4Mux_h
    port map (
            O => \N__69105\,
            I => \N__69092\
        );

    \I__16877\ : Span12Mux_v
    port map (
            O => \N__69102\,
            I => \N__69089\
        );

    \I__16876\ : Odrv4
    port map (
            O => \N__69097\,
            I => n19128
        );

    \I__16875\ : Odrv4
    port map (
            O => \N__69092\,
            I => n19128
        );

    \I__16874\ : Odrv12
    port map (
            O => \N__69089\,
            I => n19128
        );

    \I__16873\ : InMux
    port map (
            O => \N__69082\,
            I => \N__69071\
        );

    \I__16872\ : InMux
    port map (
            O => \N__69081\,
            I => \N__69071\
        );

    \I__16871\ : InMux
    port map (
            O => \N__69080\,
            I => \N__69071\
        );

    \I__16870\ : InMux
    port map (
            O => \N__69079\,
            I => \N__69066\
        );

    \I__16869\ : InMux
    port map (
            O => \N__69078\,
            I => \N__69066\
        );

    \I__16868\ : LocalMux
    port map (
            O => \N__69071\,
            I => \N__69063\
        );

    \I__16867\ : LocalMux
    port map (
            O => \N__69066\,
            I => \N__69060\
        );

    \I__16866\ : Span4Mux_v
    port map (
            O => \N__69063\,
            I => \N__69057\
        );

    \I__16865\ : Span4Mux_v
    port map (
            O => \N__69060\,
            I => \N__69050\
        );

    \I__16864\ : Span4Mux_v
    port map (
            O => \N__69057\,
            I => \N__69050\
        );

    \I__16863\ : InMux
    port map (
            O => \N__69056\,
            I => \N__69045\
        );

    \I__16862\ : InMux
    port map (
            O => \N__69055\,
            I => \N__69045\
        );

    \I__16861\ : Odrv4
    port map (
            O => \N__69050\,
            I => data_in_frame_19_3
        );

    \I__16860\ : LocalMux
    port map (
            O => \N__69045\,
            I => data_in_frame_19_3
        );

    \I__16859\ : InMux
    port map (
            O => \N__69040\,
            I => \N__69037\
        );

    \I__16858\ : LocalMux
    port map (
            O => \N__69037\,
            I => \N__69032\
        );

    \I__16857\ : InMux
    port map (
            O => \N__69036\,
            I => \N__69026\
        );

    \I__16856\ : InMux
    port map (
            O => \N__69035\,
            I => \N__69026\
        );

    \I__16855\ : Span4Mux_v
    port map (
            O => \N__69032\,
            I => \N__69019\
        );

    \I__16854\ : InMux
    port map (
            O => \N__69031\,
            I => \N__69016\
        );

    \I__16853\ : LocalMux
    port map (
            O => \N__69026\,
            I => \N__69008\
        );

    \I__16852\ : CascadeMux
    port map (
            O => \N__69025\,
            I => \N__69003\
        );

    \I__16851\ : InMux
    port map (
            O => \N__69024\,
            I => \N__68998\
        );

    \I__16850\ : CascadeMux
    port map (
            O => \N__69023\,
            I => \N__68995\
        );

    \I__16849\ : InMux
    port map (
            O => \N__69022\,
            I => \N__68991\
        );

    \I__16848\ : Span4Mux_h
    port map (
            O => \N__69019\,
            I => \N__68986\
        );

    \I__16847\ : LocalMux
    port map (
            O => \N__69016\,
            I => \N__68986\
        );

    \I__16846\ : InMux
    port map (
            O => \N__69015\,
            I => \N__68981\
        );

    \I__16845\ : InMux
    port map (
            O => \N__69014\,
            I => \N__68981\
        );

    \I__16844\ : InMux
    port map (
            O => \N__69013\,
            I => \N__68977\
        );

    \I__16843\ : InMux
    port map (
            O => \N__69012\,
            I => \N__68974\
        );

    \I__16842\ : InMux
    port map (
            O => \N__69011\,
            I => \N__68970\
        );

    \I__16841\ : Span4Mux_v
    port map (
            O => \N__69008\,
            I => \N__68967\
        );

    \I__16840\ : InMux
    port map (
            O => \N__69007\,
            I => \N__68964\
        );

    \I__16839\ : InMux
    port map (
            O => \N__69006\,
            I => \N__68961\
        );

    \I__16838\ : InMux
    port map (
            O => \N__69003\,
            I => \N__68956\
        );

    \I__16837\ : InMux
    port map (
            O => \N__69002\,
            I => \N__68956\
        );

    \I__16836\ : InMux
    port map (
            O => \N__69001\,
            I => \N__68953\
        );

    \I__16835\ : LocalMux
    port map (
            O => \N__68998\,
            I => \N__68950\
        );

    \I__16834\ : InMux
    port map (
            O => \N__68995\,
            I => \N__68945\
        );

    \I__16833\ : InMux
    port map (
            O => \N__68994\,
            I => \N__68945\
        );

    \I__16832\ : LocalMux
    port map (
            O => \N__68991\,
            I => \N__68938\
        );

    \I__16831\ : Span4Mux_v
    port map (
            O => \N__68986\,
            I => \N__68938\
        );

    \I__16830\ : LocalMux
    port map (
            O => \N__68981\,
            I => \N__68938\
        );

    \I__16829\ : InMux
    port map (
            O => \N__68980\,
            I => \N__68935\
        );

    \I__16828\ : LocalMux
    port map (
            O => \N__68977\,
            I => \N__68932\
        );

    \I__16827\ : LocalMux
    port map (
            O => \N__68974\,
            I => \N__68929\
        );

    \I__16826\ : CascadeMux
    port map (
            O => \N__68973\,
            I => \N__68924\
        );

    \I__16825\ : LocalMux
    port map (
            O => \N__68970\,
            I => \N__68920\
        );

    \I__16824\ : Span4Mux_h
    port map (
            O => \N__68967\,
            I => \N__68917\
        );

    \I__16823\ : LocalMux
    port map (
            O => \N__68964\,
            I => \N__68912\
        );

    \I__16822\ : LocalMux
    port map (
            O => \N__68961\,
            I => \N__68912\
        );

    \I__16821\ : LocalMux
    port map (
            O => \N__68956\,
            I => \N__68909\
        );

    \I__16820\ : LocalMux
    port map (
            O => \N__68953\,
            I => \N__68904\
        );

    \I__16819\ : Span4Mux_v
    port map (
            O => \N__68950\,
            I => \N__68904\
        );

    \I__16818\ : LocalMux
    port map (
            O => \N__68945\,
            I => \N__68898\
        );

    \I__16817\ : Span4Mux_v
    port map (
            O => \N__68938\,
            I => \N__68898\
        );

    \I__16816\ : LocalMux
    port map (
            O => \N__68935\,
            I => \N__68895\
        );

    \I__16815\ : Span4Mux_v
    port map (
            O => \N__68932\,
            I => \N__68890\
        );

    \I__16814\ : Span4Mux_h
    port map (
            O => \N__68929\,
            I => \N__68890\
        );

    \I__16813\ : InMux
    port map (
            O => \N__68928\,
            I => \N__68887\
        );

    \I__16812\ : InMux
    port map (
            O => \N__68927\,
            I => \N__68882\
        );

    \I__16811\ : InMux
    port map (
            O => \N__68924\,
            I => \N__68882\
        );

    \I__16810\ : InMux
    port map (
            O => \N__68923\,
            I => \N__68879\
        );

    \I__16809\ : Span4Mux_h
    port map (
            O => \N__68920\,
            I => \N__68872\
        );

    \I__16808\ : Span4Mux_v
    port map (
            O => \N__68917\,
            I => \N__68872\
        );

    \I__16807\ : Span4Mux_v
    port map (
            O => \N__68912\,
            I => \N__68872\
        );

    \I__16806\ : Span4Mux_h
    port map (
            O => \N__68909\,
            I => \N__68867\
        );

    \I__16805\ : Span4Mux_v
    port map (
            O => \N__68904\,
            I => \N__68867\
        );

    \I__16804\ : InMux
    port map (
            O => \N__68903\,
            I => \N__68863\
        );

    \I__16803\ : Span4Mux_h
    port map (
            O => \N__68898\,
            I => \N__68860\
        );

    \I__16802\ : Span4Mux_v
    port map (
            O => \N__68895\,
            I => \N__68855\
        );

    \I__16801\ : Span4Mux_v
    port map (
            O => \N__68890\,
            I => \N__68855\
        );

    \I__16800\ : LocalMux
    port map (
            O => \N__68887\,
            I => \N__68850\
        );

    \I__16799\ : LocalMux
    port map (
            O => \N__68882\,
            I => \N__68845\
        );

    \I__16798\ : LocalMux
    port map (
            O => \N__68879\,
            I => \N__68845\
        );

    \I__16797\ : Span4Mux_v
    port map (
            O => \N__68872\,
            I => \N__68840\
        );

    \I__16796\ : Span4Mux_v
    port map (
            O => \N__68867\,
            I => \N__68837\
        );

    \I__16795\ : InMux
    port map (
            O => \N__68866\,
            I => \N__68834\
        );

    \I__16794\ : LocalMux
    port map (
            O => \N__68863\,
            I => \N__68827\
        );

    \I__16793\ : Span4Mux_v
    port map (
            O => \N__68860\,
            I => \N__68827\
        );

    \I__16792\ : Span4Mux_v
    port map (
            O => \N__68855\,
            I => \N__68827\
        );

    \I__16791\ : CascadeMux
    port map (
            O => \N__68854\,
            I => \N__68821\
        );

    \I__16790\ : InMux
    port map (
            O => \N__68853\,
            I => \N__68818\
        );

    \I__16789\ : Span4Mux_v
    port map (
            O => \N__68850\,
            I => \N__68813\
        );

    \I__16788\ : Span4Mux_v
    port map (
            O => \N__68845\,
            I => \N__68813\
        );

    \I__16787\ : InMux
    port map (
            O => \N__68844\,
            I => \N__68808\
        );

    \I__16786\ : InMux
    port map (
            O => \N__68843\,
            I => \N__68808\
        );

    \I__16785\ : Span4Mux_h
    port map (
            O => \N__68840\,
            I => \N__68803\
        );

    \I__16784\ : Span4Mux_h
    port map (
            O => \N__68837\,
            I => \N__68803\
        );

    \I__16783\ : LocalMux
    port map (
            O => \N__68834\,
            I => \N__68800\
        );

    \I__16782\ : Span4Mux_h
    port map (
            O => \N__68827\,
            I => \N__68797\
        );

    \I__16781\ : InMux
    port map (
            O => \N__68826\,
            I => \N__68794\
        );

    \I__16780\ : InMux
    port map (
            O => \N__68825\,
            I => \N__68789\
        );

    \I__16779\ : InMux
    port map (
            O => \N__68824\,
            I => \N__68789\
        );

    \I__16778\ : InMux
    port map (
            O => \N__68821\,
            I => \N__68786\
        );

    \I__16777\ : LocalMux
    port map (
            O => \N__68818\,
            I => \N__68781\
        );

    \I__16776\ : Span4Mux_h
    port map (
            O => \N__68813\,
            I => \N__68781\
        );

    \I__16775\ : LocalMux
    port map (
            O => \N__68808\,
            I => \N__68776\
        );

    \I__16774\ : Span4Mux_h
    port map (
            O => \N__68803\,
            I => \N__68776\
        );

    \I__16773\ : Span4Mux_v
    port map (
            O => \N__68800\,
            I => \N__68771\
        );

    \I__16772\ : Span4Mux_h
    port map (
            O => \N__68797\,
            I => \N__68771\
        );

    \I__16771\ : LocalMux
    port map (
            O => \N__68794\,
            I => rx_data_6
        );

    \I__16770\ : LocalMux
    port map (
            O => \N__68789\,
            I => rx_data_6
        );

    \I__16769\ : LocalMux
    port map (
            O => \N__68786\,
            I => rx_data_6
        );

    \I__16768\ : Odrv4
    port map (
            O => \N__68781\,
            I => rx_data_6
        );

    \I__16767\ : Odrv4
    port map (
            O => \N__68776\,
            I => rx_data_6
        );

    \I__16766\ : Odrv4
    port map (
            O => \N__68771\,
            I => rx_data_6
        );

    \I__16765\ : CascadeMux
    port map (
            O => \N__68758\,
            I => \N__68755\
        );

    \I__16764\ : InMux
    port map (
            O => \N__68755\,
            I => \N__68752\
        );

    \I__16763\ : LocalMux
    port map (
            O => \N__68752\,
            I => \N__68747\
        );

    \I__16762\ : CascadeMux
    port map (
            O => \N__68751\,
            I => \N__68741\
        );

    \I__16761\ : InMux
    port map (
            O => \N__68750\,
            I => \N__68737\
        );

    \I__16760\ : Span4Mux_v
    port map (
            O => \N__68747\,
            I => \N__68734\
        );

    \I__16759\ : InMux
    port map (
            O => \N__68746\,
            I => \N__68731\
        );

    \I__16758\ : InMux
    port map (
            O => \N__68745\,
            I => \N__68728\
        );

    \I__16757\ : InMux
    port map (
            O => \N__68744\,
            I => \N__68719\
        );

    \I__16756\ : InMux
    port map (
            O => \N__68741\,
            I => \N__68716\
        );

    \I__16755\ : InMux
    port map (
            O => \N__68740\,
            I => \N__68713\
        );

    \I__16754\ : LocalMux
    port map (
            O => \N__68737\,
            I => \N__68708\
        );

    \I__16753\ : Span4Mux_h
    port map (
            O => \N__68734\,
            I => \N__68701\
        );

    \I__16752\ : LocalMux
    port map (
            O => \N__68731\,
            I => \N__68701\
        );

    \I__16751\ : LocalMux
    port map (
            O => \N__68728\,
            I => \N__68701\
        );

    \I__16750\ : InMux
    port map (
            O => \N__68727\,
            I => \N__68698\
        );

    \I__16749\ : InMux
    port map (
            O => \N__68726\,
            I => \N__68695\
        );

    \I__16748\ : InMux
    port map (
            O => \N__68725\,
            I => \N__68692\
        );

    \I__16747\ : CascadeMux
    port map (
            O => \N__68724\,
            I => \N__68688\
        );

    \I__16746\ : InMux
    port map (
            O => \N__68723\,
            I => \N__68683\
        );

    \I__16745\ : InMux
    port map (
            O => \N__68722\,
            I => \N__68683\
        );

    \I__16744\ : LocalMux
    port map (
            O => \N__68719\,
            I => \N__68675\
        );

    \I__16743\ : LocalMux
    port map (
            O => \N__68716\,
            I => \N__68675\
        );

    \I__16742\ : LocalMux
    port map (
            O => \N__68713\,
            I => \N__68675\
        );

    \I__16741\ : InMux
    port map (
            O => \N__68712\,
            I => \N__68671\
        );

    \I__16740\ : InMux
    port map (
            O => \N__68711\,
            I => \N__68668\
        );

    \I__16739\ : Span4Mux_v
    port map (
            O => \N__68708\,
            I => \N__68657\
        );

    \I__16738\ : Span4Mux_v
    port map (
            O => \N__68701\,
            I => \N__68657\
        );

    \I__16737\ : LocalMux
    port map (
            O => \N__68698\,
            I => \N__68657\
        );

    \I__16736\ : LocalMux
    port map (
            O => \N__68695\,
            I => \N__68657\
        );

    \I__16735\ : LocalMux
    port map (
            O => \N__68692\,
            I => \N__68657\
        );

    \I__16734\ : InMux
    port map (
            O => \N__68691\,
            I => \N__68652\
        );

    \I__16733\ : InMux
    port map (
            O => \N__68688\,
            I => \N__68649\
        );

    \I__16732\ : LocalMux
    port map (
            O => \N__68683\,
            I => \N__68641\
        );

    \I__16731\ : InMux
    port map (
            O => \N__68682\,
            I => \N__68638\
        );

    \I__16730\ : Span4Mux_v
    port map (
            O => \N__68675\,
            I => \N__68635\
        );

    \I__16729\ : InMux
    port map (
            O => \N__68674\,
            I => \N__68632\
        );

    \I__16728\ : LocalMux
    port map (
            O => \N__68671\,
            I => \N__68629\
        );

    \I__16727\ : LocalMux
    port map (
            O => \N__68668\,
            I => \N__68626\
        );

    \I__16726\ : Span4Mux_v
    port map (
            O => \N__68657\,
            I => \N__68623\
        );

    \I__16725\ : InMux
    port map (
            O => \N__68656\,
            I => \N__68619\
        );

    \I__16724\ : InMux
    port map (
            O => \N__68655\,
            I => \N__68616\
        );

    \I__16723\ : LocalMux
    port map (
            O => \N__68652\,
            I => \N__68613\
        );

    \I__16722\ : LocalMux
    port map (
            O => \N__68649\,
            I => \N__68609\
        );

    \I__16721\ : InMux
    port map (
            O => \N__68648\,
            I => \N__68604\
        );

    \I__16720\ : InMux
    port map (
            O => \N__68647\,
            I => \N__68604\
        );

    \I__16719\ : InMux
    port map (
            O => \N__68646\,
            I => \N__68601\
        );

    \I__16718\ : InMux
    port map (
            O => \N__68645\,
            I => \N__68598\
        );

    \I__16717\ : InMux
    port map (
            O => \N__68644\,
            I => \N__68595\
        );

    \I__16716\ : Span4Mux_h
    port map (
            O => \N__68641\,
            I => \N__68590\
        );

    \I__16715\ : LocalMux
    port map (
            O => \N__68638\,
            I => \N__68587\
        );

    \I__16714\ : Span4Mux_h
    port map (
            O => \N__68635\,
            I => \N__68584\
        );

    \I__16713\ : LocalMux
    port map (
            O => \N__68632\,
            I => \N__68581\
        );

    \I__16712\ : Span4Mux_h
    port map (
            O => \N__68629\,
            I => \N__68576\
        );

    \I__16711\ : Span4Mux_h
    port map (
            O => \N__68626\,
            I => \N__68576\
        );

    \I__16710\ : Span4Mux_h
    port map (
            O => \N__68623\,
            I => \N__68573\
        );

    \I__16709\ : InMux
    port map (
            O => \N__68622\,
            I => \N__68570\
        );

    \I__16708\ : LocalMux
    port map (
            O => \N__68619\,
            I => \N__68565\
        );

    \I__16707\ : LocalMux
    port map (
            O => \N__68616\,
            I => \N__68565\
        );

    \I__16706\ : Span4Mux_h
    port map (
            O => \N__68613\,
            I => \N__68562\
        );

    \I__16705\ : InMux
    port map (
            O => \N__68612\,
            I => \N__68559\
        );

    \I__16704\ : Span4Mux_h
    port map (
            O => \N__68609\,
            I => \N__68554\
        );

    \I__16703\ : LocalMux
    port map (
            O => \N__68604\,
            I => \N__68554\
        );

    \I__16702\ : LocalMux
    port map (
            O => \N__68601\,
            I => \N__68546\
        );

    \I__16701\ : LocalMux
    port map (
            O => \N__68598\,
            I => \N__68546\
        );

    \I__16700\ : LocalMux
    port map (
            O => \N__68595\,
            I => \N__68546\
        );

    \I__16699\ : InMux
    port map (
            O => \N__68594\,
            I => \N__68543\
        );

    \I__16698\ : InMux
    port map (
            O => \N__68593\,
            I => \N__68540\
        );

    \I__16697\ : Span4Mux_v
    port map (
            O => \N__68590\,
            I => \N__68535\
        );

    \I__16696\ : Span4Mux_h
    port map (
            O => \N__68587\,
            I => \N__68535\
        );

    \I__16695\ : Sp12to4
    port map (
            O => \N__68584\,
            I => \N__68532\
        );

    \I__16694\ : Span4Mux_h
    port map (
            O => \N__68581\,
            I => \N__68529\
        );

    \I__16693\ : Span4Mux_v
    port map (
            O => \N__68576\,
            I => \N__68526\
        );

    \I__16692\ : Span4Mux_v
    port map (
            O => \N__68573\,
            I => \N__68523\
        );

    \I__16691\ : LocalMux
    port map (
            O => \N__68570\,
            I => \N__68518\
        );

    \I__16690\ : Sp12to4
    port map (
            O => \N__68565\,
            I => \N__68515\
        );

    \I__16689\ : Span4Mux_h
    port map (
            O => \N__68562\,
            I => \N__68512\
        );

    \I__16688\ : LocalMux
    port map (
            O => \N__68559\,
            I => \N__68509\
        );

    \I__16687\ : Span4Mux_v
    port map (
            O => \N__68554\,
            I => \N__68506\
        );

    \I__16686\ : InMux
    port map (
            O => \N__68553\,
            I => \N__68503\
        );

    \I__16685\ : Span4Mux_v
    port map (
            O => \N__68546\,
            I => \N__68500\
        );

    \I__16684\ : LocalMux
    port map (
            O => \N__68543\,
            I => \N__68495\
        );

    \I__16683\ : LocalMux
    port map (
            O => \N__68540\,
            I => \N__68495\
        );

    \I__16682\ : Sp12to4
    port map (
            O => \N__68535\,
            I => \N__68492\
        );

    \I__16681\ : Span12Mux_h
    port map (
            O => \N__68532\,
            I => \N__68489\
        );

    \I__16680\ : Span4Mux_v
    port map (
            O => \N__68529\,
            I => \N__68484\
        );

    \I__16679\ : Span4Mux_v
    port map (
            O => \N__68526\,
            I => \N__68484\
        );

    \I__16678\ : Sp12to4
    port map (
            O => \N__68523\,
            I => \N__68481\
        );

    \I__16677\ : InMux
    port map (
            O => \N__68522\,
            I => \N__68476\
        );

    \I__16676\ : InMux
    port map (
            O => \N__68521\,
            I => \N__68476\
        );

    \I__16675\ : Span4Mux_v
    port map (
            O => \N__68518\,
            I => \N__68473\
        );

    \I__16674\ : Span12Mux_v
    port map (
            O => \N__68515\,
            I => \N__68470\
        );

    \I__16673\ : Span4Mux_v
    port map (
            O => \N__68512\,
            I => \N__68463\
        );

    \I__16672\ : Span4Mux_v
    port map (
            O => \N__68509\,
            I => \N__68463\
        );

    \I__16671\ : Span4Mux_v
    port map (
            O => \N__68506\,
            I => \N__68463\
        );

    \I__16670\ : LocalMux
    port map (
            O => \N__68503\,
            I => \N__68456\
        );

    \I__16669\ : Span4Mux_v
    port map (
            O => \N__68500\,
            I => \N__68456\
        );

    \I__16668\ : Span4Mux_h
    port map (
            O => \N__68495\,
            I => \N__68456\
        );

    \I__16667\ : Span12Mux_v
    port map (
            O => \N__68492\,
            I => \N__68447\
        );

    \I__16666\ : Span12Mux_v
    port map (
            O => \N__68489\,
            I => \N__68447\
        );

    \I__16665\ : Sp12to4
    port map (
            O => \N__68484\,
            I => \N__68447\
        );

    \I__16664\ : Span12Mux_s6_h
    port map (
            O => \N__68481\,
            I => \N__68447\
        );

    \I__16663\ : LocalMux
    port map (
            O => \N__68476\,
            I => rx_data_2
        );

    \I__16662\ : Odrv4
    port map (
            O => \N__68473\,
            I => rx_data_2
        );

    \I__16661\ : Odrv12
    port map (
            O => \N__68470\,
            I => rx_data_2
        );

    \I__16660\ : Odrv4
    port map (
            O => \N__68463\,
            I => rx_data_2
        );

    \I__16659\ : Odrv4
    port map (
            O => \N__68456\,
            I => rx_data_2
        );

    \I__16658\ : Odrv12
    port map (
            O => \N__68447\,
            I => rx_data_2
        );

    \I__16657\ : InMux
    port map (
            O => \N__68434\,
            I => \N__68431\
        );

    \I__16656\ : LocalMux
    port map (
            O => \N__68431\,
            I => \N__68425\
        );

    \I__16655\ : InMux
    port map (
            O => \N__68430\,
            I => \N__68422\
        );

    \I__16654\ : InMux
    port map (
            O => \N__68429\,
            I => \N__68419\
        );

    \I__16653\ : InMux
    port map (
            O => \N__68428\,
            I => \N__68416\
        );

    \I__16652\ : Span4Mux_v
    port map (
            O => \N__68425\,
            I => \N__68413\
        );

    \I__16651\ : LocalMux
    port map (
            O => \N__68422\,
            I => \N__68410\
        );

    \I__16650\ : LocalMux
    port map (
            O => \N__68419\,
            I => \N__68405\
        );

    \I__16649\ : LocalMux
    port map (
            O => \N__68416\,
            I => \N__68405\
        );

    \I__16648\ : Span4Mux_h
    port map (
            O => \N__68413\,
            I => \N__68398\
        );

    \I__16647\ : Span4Mux_v
    port map (
            O => \N__68410\,
            I => \N__68398\
        );

    \I__16646\ : Span4Mux_h
    port map (
            O => \N__68405\,
            I => \N__68398\
        );

    \I__16645\ : Span4Mux_v
    port map (
            O => \N__68398\,
            I => \N__68395\
        );

    \I__16644\ : Odrv4
    port map (
            O => \N__68395\,
            I => \c0.n19474\
        );

    \I__16643\ : CascadeMux
    port map (
            O => \N__68392\,
            I => \N__68388\
        );

    \I__16642\ : CascadeMux
    port map (
            O => \N__68391\,
            I => \N__68385\
        );

    \I__16641\ : InMux
    port map (
            O => \N__68388\,
            I => \N__68378\
        );

    \I__16640\ : InMux
    port map (
            O => \N__68385\,
            I => \N__68378\
        );

    \I__16639\ : InMux
    port map (
            O => \N__68384\,
            I => \N__68375\
        );

    \I__16638\ : InMux
    port map (
            O => \N__68383\,
            I => \N__68371\
        );

    \I__16637\ : LocalMux
    port map (
            O => \N__68378\,
            I => \N__68368\
        );

    \I__16636\ : LocalMux
    port map (
            O => \N__68375\,
            I => \N__68365\
        );

    \I__16635\ : InMux
    port map (
            O => \N__68374\,
            I => \N__68361\
        );

    \I__16634\ : LocalMux
    port map (
            O => \N__68371\,
            I => \N__68356\
        );

    \I__16633\ : Span4Mux_v
    port map (
            O => \N__68368\,
            I => \N__68356\
        );

    \I__16632\ : Span4Mux_v
    port map (
            O => \N__68365\,
            I => \N__68352\
        );

    \I__16631\ : CascadeMux
    port map (
            O => \N__68364\,
            I => \N__68349\
        );

    \I__16630\ : LocalMux
    port map (
            O => \N__68361\,
            I => \N__68345\
        );

    \I__16629\ : Span4Mux_v
    port map (
            O => \N__68356\,
            I => \N__68342\
        );

    \I__16628\ : InMux
    port map (
            O => \N__68355\,
            I => \N__68339\
        );

    \I__16627\ : Span4Mux_h
    port map (
            O => \N__68352\,
            I => \N__68336\
        );

    \I__16626\ : InMux
    port map (
            O => \N__68349\,
            I => \N__68333\
        );

    \I__16625\ : InMux
    port map (
            O => \N__68348\,
            I => \N__68330\
        );

    \I__16624\ : Span12Mux_h
    port map (
            O => \N__68345\,
            I => \N__68327\
        );

    \I__16623\ : Span4Mux_h
    port map (
            O => \N__68342\,
            I => \N__68324\
        );

    \I__16622\ : LocalMux
    port map (
            O => \N__68339\,
            I => \N__68317\
        );

    \I__16621\ : Span4Mux_h
    port map (
            O => \N__68336\,
            I => \N__68317\
        );

    \I__16620\ : LocalMux
    port map (
            O => \N__68333\,
            I => \N__68317\
        );

    \I__16619\ : LocalMux
    port map (
            O => \N__68330\,
            I => \c0.data_in_frame_17_2\
        );

    \I__16618\ : Odrv12
    port map (
            O => \N__68327\,
            I => \c0.data_in_frame_17_2\
        );

    \I__16617\ : Odrv4
    port map (
            O => \N__68324\,
            I => \c0.data_in_frame_17_2\
        );

    \I__16616\ : Odrv4
    port map (
            O => \N__68317\,
            I => \c0.data_in_frame_17_2\
        );

    \I__16615\ : InMux
    port map (
            O => \N__68308\,
            I => \N__68304\
        );

    \I__16614\ : InMux
    port map (
            O => \N__68307\,
            I => \N__68301\
        );

    \I__16613\ : LocalMux
    port map (
            O => \N__68304\,
            I => \N__68296\
        );

    \I__16612\ : LocalMux
    port map (
            O => \N__68301\,
            I => \N__68293\
        );

    \I__16611\ : InMux
    port map (
            O => \N__68300\,
            I => \N__68290\
        );

    \I__16610\ : InMux
    port map (
            O => \N__68299\,
            I => \N__68286\
        );

    \I__16609\ : Span4Mux_h
    port map (
            O => \N__68296\,
            I => \N__68283\
        );

    \I__16608\ : Span4Mux_h
    port map (
            O => \N__68293\,
            I => \N__68278\
        );

    \I__16607\ : LocalMux
    port map (
            O => \N__68290\,
            I => \N__68278\
        );

    \I__16606\ : InMux
    port map (
            O => \N__68289\,
            I => \N__68275\
        );

    \I__16605\ : LocalMux
    port map (
            O => \N__68286\,
            I => \N__68271\
        );

    \I__16604\ : Span4Mux_h
    port map (
            O => \N__68283\,
            I => \N__68266\
        );

    \I__16603\ : Span4Mux_h
    port map (
            O => \N__68278\,
            I => \N__68266\
        );

    \I__16602\ : LocalMux
    port map (
            O => \N__68275\,
            I => \N__68263\
        );

    \I__16601\ : InMux
    port map (
            O => \N__68274\,
            I => \N__68260\
        );

    \I__16600\ : Span4Mux_v
    port map (
            O => \N__68271\,
            I => \N__68257\
        );

    \I__16599\ : Span4Mux_v
    port map (
            O => \N__68266\,
            I => \N__68252\
        );

    \I__16598\ : Span4Mux_h
    port map (
            O => \N__68263\,
            I => \N__68252\
        );

    \I__16597\ : LocalMux
    port map (
            O => \N__68260\,
            I => \c0.data_in_frame_17_3\
        );

    \I__16596\ : Odrv4
    port map (
            O => \N__68257\,
            I => \c0.data_in_frame_17_3\
        );

    \I__16595\ : Odrv4
    port map (
            O => \N__68252\,
            I => \c0.data_in_frame_17_3\
        );

    \I__16594\ : InMux
    port map (
            O => \N__68245\,
            I => \N__68242\
        );

    \I__16593\ : LocalMux
    port map (
            O => \N__68242\,
            I => \N__68239\
        );

    \I__16592\ : Odrv4
    port map (
            O => \N__68239\,
            I => \c0.n14_adj_3436\
        );

    \I__16591\ : InMux
    port map (
            O => \N__68236\,
            I => \N__68229\
        );

    \I__16590\ : InMux
    port map (
            O => \N__68235\,
            I => \N__68229\
        );

    \I__16589\ : InMux
    port map (
            O => \N__68234\,
            I => \N__68224\
        );

    \I__16588\ : LocalMux
    port map (
            O => \N__68229\,
            I => \N__68221\
        );

    \I__16587\ : CascadeMux
    port map (
            O => \N__68228\,
            I => \N__68218\
        );

    \I__16586\ : InMux
    port map (
            O => \N__68227\,
            I => \N__68214\
        );

    \I__16585\ : LocalMux
    port map (
            O => \N__68224\,
            I => \N__68208\
        );

    \I__16584\ : Span4Mux_h
    port map (
            O => \N__68221\,
            I => \N__68208\
        );

    \I__16583\ : InMux
    port map (
            O => \N__68218\,
            I => \N__68203\
        );

    \I__16582\ : InMux
    port map (
            O => \N__68217\,
            I => \N__68203\
        );

    \I__16581\ : LocalMux
    port map (
            O => \N__68214\,
            I => \N__68200\
        );

    \I__16580\ : InMux
    port map (
            O => \N__68213\,
            I => \N__68197\
        );

    \I__16579\ : Span4Mux_v
    port map (
            O => \N__68208\,
            I => \N__68192\
        );

    \I__16578\ : LocalMux
    port map (
            O => \N__68203\,
            I => \N__68185\
        );

    \I__16577\ : Span4Mux_h
    port map (
            O => \N__68200\,
            I => \N__68185\
        );

    \I__16576\ : LocalMux
    port map (
            O => \N__68197\,
            I => \N__68185\
        );

    \I__16575\ : InMux
    port map (
            O => \N__68196\,
            I => \N__68180\
        );

    \I__16574\ : InMux
    port map (
            O => \N__68195\,
            I => \N__68180\
        );

    \I__16573\ : Odrv4
    port map (
            O => \N__68192\,
            I => \c0.data_in_frame_20_4\
        );

    \I__16572\ : Odrv4
    port map (
            O => \N__68185\,
            I => \c0.data_in_frame_20_4\
        );

    \I__16571\ : LocalMux
    port map (
            O => \N__68180\,
            I => \c0.data_in_frame_20_4\
        );

    \I__16570\ : CascadeMux
    port map (
            O => \N__68173\,
            I => \N__68170\
        );

    \I__16569\ : InMux
    port map (
            O => \N__68170\,
            I => \N__68166\
        );

    \I__16568\ : InMux
    port map (
            O => \N__68169\,
            I => \N__68162\
        );

    \I__16567\ : LocalMux
    port map (
            O => \N__68166\,
            I => \N__68159\
        );

    \I__16566\ : InMux
    port map (
            O => \N__68165\,
            I => \N__68154\
        );

    \I__16565\ : LocalMux
    port map (
            O => \N__68162\,
            I => \N__68151\
        );

    \I__16564\ : Span4Mux_v
    port map (
            O => \N__68159\,
            I => \N__68148\
        );

    \I__16563\ : InMux
    port map (
            O => \N__68158\,
            I => \N__68143\
        );

    \I__16562\ : InMux
    port map (
            O => \N__68157\,
            I => \N__68143\
        );

    \I__16561\ : LocalMux
    port map (
            O => \N__68154\,
            I => \N__68140\
        );

    \I__16560\ : Span4Mux_v
    port map (
            O => \N__68151\,
            I => \N__68133\
        );

    \I__16559\ : Span4Mux_h
    port map (
            O => \N__68148\,
            I => \N__68133\
        );

    \I__16558\ : LocalMux
    port map (
            O => \N__68143\,
            I => \N__68133\
        );

    \I__16557\ : Span12Mux_v
    port map (
            O => \N__68140\,
            I => \N__68130\
        );

    \I__16556\ : Odrv4
    port map (
            O => \N__68133\,
            I => \c0.n19274\
        );

    \I__16555\ : Odrv12
    port map (
            O => \N__68130\,
            I => \c0.n19274\
        );

    \I__16554\ : CascadeMux
    port map (
            O => \N__68125\,
            I => \N__68121\
        );

    \I__16553\ : InMux
    port map (
            O => \N__68124\,
            I => \N__68114\
        );

    \I__16552\ : InMux
    port map (
            O => \N__68121\,
            I => \N__68114\
        );

    \I__16551\ : InMux
    port map (
            O => \N__68120\,
            I => \N__68109\
        );

    \I__16550\ : InMux
    port map (
            O => \N__68119\,
            I => \N__68106\
        );

    \I__16549\ : LocalMux
    port map (
            O => \N__68114\,
            I => \N__68101\
        );

    \I__16548\ : InMux
    port map (
            O => \N__68113\,
            I => \N__68096\
        );

    \I__16547\ : InMux
    port map (
            O => \N__68112\,
            I => \N__68096\
        );

    \I__16546\ : LocalMux
    port map (
            O => \N__68109\,
            I => \N__68093\
        );

    \I__16545\ : LocalMux
    port map (
            O => \N__68106\,
            I => \N__68090\
        );

    \I__16544\ : InMux
    port map (
            O => \N__68105\,
            I => \N__68085\
        );

    \I__16543\ : InMux
    port map (
            O => \N__68104\,
            I => \N__68085\
        );

    \I__16542\ : Span4Mux_h
    port map (
            O => \N__68101\,
            I => \N__68081\
        );

    \I__16541\ : LocalMux
    port map (
            O => \N__68096\,
            I => \N__68076\
        );

    \I__16540\ : Span4Mux_v
    port map (
            O => \N__68093\,
            I => \N__68076\
        );

    \I__16539\ : Span4Mux_h
    port map (
            O => \N__68090\,
            I => \N__68071\
        );

    \I__16538\ : LocalMux
    port map (
            O => \N__68085\,
            I => \N__68071\
        );

    \I__16537\ : InMux
    port map (
            O => \N__68084\,
            I => \N__68067\
        );

    \I__16536\ : Span4Mux_v
    port map (
            O => \N__68081\,
            I => \N__68064\
        );

    \I__16535\ : Span4Mux_h
    port map (
            O => \N__68076\,
            I => \N__68059\
        );

    \I__16534\ : Span4Mux_v
    port map (
            O => \N__68071\,
            I => \N__68059\
        );

    \I__16533\ : InMux
    port map (
            O => \N__68070\,
            I => \N__68056\
        );

    \I__16532\ : LocalMux
    port map (
            O => \N__68067\,
            I => \c0.data_in_frame_20_3\
        );

    \I__16531\ : Odrv4
    port map (
            O => \N__68064\,
            I => \c0.data_in_frame_20_3\
        );

    \I__16530\ : Odrv4
    port map (
            O => \N__68059\,
            I => \c0.data_in_frame_20_3\
        );

    \I__16529\ : LocalMux
    port map (
            O => \N__68056\,
            I => \c0.data_in_frame_20_3\
        );

    \I__16528\ : CascadeMux
    port map (
            O => \N__68047\,
            I => \N__68044\
        );

    \I__16527\ : InMux
    port map (
            O => \N__68044\,
            I => \N__68040\
        );

    \I__16526\ : InMux
    port map (
            O => \N__68043\,
            I => \N__68037\
        );

    \I__16525\ : LocalMux
    port map (
            O => \N__68040\,
            I => \N__68034\
        );

    \I__16524\ : LocalMux
    port map (
            O => \N__68037\,
            I => \N__68031\
        );

    \I__16523\ : Span4Mux_h
    port map (
            O => \N__68034\,
            I => \N__68026\
        );

    \I__16522\ : Span4Mux_v
    port map (
            O => \N__68031\,
            I => \N__68026\
        );

    \I__16521\ : Odrv4
    port map (
            O => \N__68026\,
            I => \c0.n54_adj_3388\
        );

    \I__16520\ : InMux
    port map (
            O => \N__68023\,
            I => \N__68019\
        );

    \I__16519\ : InMux
    port map (
            O => \N__68022\,
            I => \N__68014\
        );

    \I__16518\ : LocalMux
    port map (
            O => \N__68019\,
            I => \N__68011\
        );

    \I__16517\ : InMux
    port map (
            O => \N__68018\,
            I => \N__68008\
        );

    \I__16516\ : InMux
    port map (
            O => \N__68017\,
            I => \N__68005\
        );

    \I__16515\ : LocalMux
    port map (
            O => \N__68014\,
            I => \N__68002\
        );

    \I__16514\ : Odrv12
    port map (
            O => \N__68011\,
            I => \c0.n32_adj_3310\
        );

    \I__16513\ : LocalMux
    port map (
            O => \N__68008\,
            I => \c0.n32_adj_3310\
        );

    \I__16512\ : LocalMux
    port map (
            O => \N__68005\,
            I => \c0.n32_adj_3310\
        );

    \I__16511\ : Odrv4
    port map (
            O => \N__68002\,
            I => \c0.n32_adj_3310\
        );

    \I__16510\ : InMux
    port map (
            O => \N__67993\,
            I => \N__67990\
        );

    \I__16509\ : LocalMux
    port map (
            O => \N__67990\,
            I => \c0.n43_adj_3131\
        );

    \I__16508\ : InMux
    port map (
            O => \N__67987\,
            I => \N__67984\
        );

    \I__16507\ : LocalMux
    port map (
            O => \N__67984\,
            I => \N__67976\
        );

    \I__16506\ : InMux
    port map (
            O => \N__67983\,
            I => \N__67973\
        );

    \I__16505\ : InMux
    port map (
            O => \N__67982\,
            I => \N__67968\
        );

    \I__16504\ : InMux
    port map (
            O => \N__67981\,
            I => \N__67965\
        );

    \I__16503\ : InMux
    port map (
            O => \N__67980\,
            I => \N__67961\
        );

    \I__16502\ : InMux
    port map (
            O => \N__67979\,
            I => \N__67958\
        );

    \I__16501\ : Span4Mux_h
    port map (
            O => \N__67976\,
            I => \N__67953\
        );

    \I__16500\ : LocalMux
    port map (
            O => \N__67973\,
            I => \N__67953\
        );

    \I__16499\ : InMux
    port map (
            O => \N__67972\,
            I => \N__67941\
        );

    \I__16498\ : InMux
    port map (
            O => \N__67971\,
            I => \N__67936\
        );

    \I__16497\ : LocalMux
    port map (
            O => \N__67968\,
            I => \N__67933\
        );

    \I__16496\ : LocalMux
    port map (
            O => \N__67965\,
            I => \N__67929\
        );

    \I__16495\ : InMux
    port map (
            O => \N__67964\,
            I => \N__67926\
        );

    \I__16494\ : LocalMux
    port map (
            O => \N__67961\,
            I => \N__67923\
        );

    \I__16493\ : LocalMux
    port map (
            O => \N__67958\,
            I => \N__67916\
        );

    \I__16492\ : Span4Mux_v
    port map (
            O => \N__67953\,
            I => \N__67913\
        );

    \I__16491\ : InMux
    port map (
            O => \N__67952\,
            I => \N__67908\
        );

    \I__16490\ : InMux
    port map (
            O => \N__67951\,
            I => \N__67905\
        );

    \I__16489\ : InMux
    port map (
            O => \N__67950\,
            I => \N__67900\
        );

    \I__16488\ : InMux
    port map (
            O => \N__67949\,
            I => \N__67900\
        );

    \I__16487\ : InMux
    port map (
            O => \N__67948\,
            I => \N__67897\
        );

    \I__16486\ : InMux
    port map (
            O => \N__67947\,
            I => \N__67890\
        );

    \I__16485\ : InMux
    port map (
            O => \N__67946\,
            I => \N__67890\
        );

    \I__16484\ : InMux
    port map (
            O => \N__67945\,
            I => \N__67890\
        );

    \I__16483\ : CascadeMux
    port map (
            O => \N__67944\,
            I => \N__67886\
        );

    \I__16482\ : LocalMux
    port map (
            O => \N__67941\,
            I => \N__67883\
        );

    \I__16481\ : InMux
    port map (
            O => \N__67940\,
            I => \N__67880\
        );

    \I__16480\ : InMux
    port map (
            O => \N__67939\,
            I => \N__67877\
        );

    \I__16479\ : LocalMux
    port map (
            O => \N__67936\,
            I => \N__67872\
        );

    \I__16478\ : Span4Mux_h
    port map (
            O => \N__67933\,
            I => \N__67872\
        );

    \I__16477\ : InMux
    port map (
            O => \N__67932\,
            I => \N__67869\
        );

    \I__16476\ : Span4Mux_h
    port map (
            O => \N__67929\,
            I => \N__67866\
        );

    \I__16475\ : LocalMux
    port map (
            O => \N__67926\,
            I => \N__67861\
        );

    \I__16474\ : Span4Mux_h
    port map (
            O => \N__67923\,
            I => \N__67861\
        );

    \I__16473\ : InMux
    port map (
            O => \N__67922\,
            I => \N__67858\
        );

    \I__16472\ : InMux
    port map (
            O => \N__67921\,
            I => \N__67855\
        );

    \I__16471\ : InMux
    port map (
            O => \N__67920\,
            I => \N__67849\
        );

    \I__16470\ : InMux
    port map (
            O => \N__67919\,
            I => \N__67849\
        );

    \I__16469\ : Span4Mux_h
    port map (
            O => \N__67916\,
            I => \N__67846\
        );

    \I__16468\ : Span4Mux_v
    port map (
            O => \N__67913\,
            I => \N__67843\
        );

    \I__16467\ : InMux
    port map (
            O => \N__67912\,
            I => \N__67840\
        );

    \I__16466\ : InMux
    port map (
            O => \N__67911\,
            I => \N__67837\
        );

    \I__16465\ : LocalMux
    port map (
            O => \N__67908\,
            I => \N__67826\
        );

    \I__16464\ : LocalMux
    port map (
            O => \N__67905\,
            I => \N__67826\
        );

    \I__16463\ : LocalMux
    port map (
            O => \N__67900\,
            I => \N__67826\
        );

    \I__16462\ : LocalMux
    port map (
            O => \N__67897\,
            I => \N__67826\
        );

    \I__16461\ : LocalMux
    port map (
            O => \N__67890\,
            I => \N__67826\
        );

    \I__16460\ : InMux
    port map (
            O => \N__67889\,
            I => \N__67821\
        );

    \I__16459\ : InMux
    port map (
            O => \N__67886\,
            I => \N__67821\
        );

    \I__16458\ : Span4Mux_v
    port map (
            O => \N__67883\,
            I => \N__67818\
        );

    \I__16457\ : LocalMux
    port map (
            O => \N__67880\,
            I => \N__67813\
        );

    \I__16456\ : LocalMux
    port map (
            O => \N__67877\,
            I => \N__67813\
        );

    \I__16455\ : Span4Mux_h
    port map (
            O => \N__67872\,
            I => \N__67808\
        );

    \I__16454\ : LocalMux
    port map (
            O => \N__67869\,
            I => \N__67808\
        );

    \I__16453\ : Span4Mux_h
    port map (
            O => \N__67866\,
            I => \N__67803\
        );

    \I__16452\ : Span4Mux_v
    port map (
            O => \N__67861\,
            I => \N__67803\
        );

    \I__16451\ : LocalMux
    port map (
            O => \N__67858\,
            I => \N__67799\
        );

    \I__16450\ : LocalMux
    port map (
            O => \N__67855\,
            I => \N__67796\
        );

    \I__16449\ : InMux
    port map (
            O => \N__67854\,
            I => \N__67793\
        );

    \I__16448\ : LocalMux
    port map (
            O => \N__67849\,
            I => \N__67790\
        );

    \I__16447\ : Span4Mux_h
    port map (
            O => \N__67846\,
            I => \N__67785\
        );

    \I__16446\ : Span4Mux_v
    port map (
            O => \N__67843\,
            I => \N__67785\
        );

    \I__16445\ : LocalMux
    port map (
            O => \N__67840\,
            I => \N__67778\
        );

    \I__16444\ : LocalMux
    port map (
            O => \N__67837\,
            I => \N__67778\
        );

    \I__16443\ : Span4Mux_v
    port map (
            O => \N__67826\,
            I => \N__67778\
        );

    \I__16442\ : LocalMux
    port map (
            O => \N__67821\,
            I => \N__67773\
        );

    \I__16441\ : Sp12to4
    port map (
            O => \N__67818\,
            I => \N__67770\
        );

    \I__16440\ : Span12Mux_h
    port map (
            O => \N__67813\,
            I => \N__67763\
        );

    \I__16439\ : Sp12to4
    port map (
            O => \N__67808\,
            I => \N__67763\
        );

    \I__16438\ : Sp12to4
    port map (
            O => \N__67803\,
            I => \N__67763\
        );

    \I__16437\ : InMux
    port map (
            O => \N__67802\,
            I => \N__67760\
        );

    \I__16436\ : Span4Mux_v
    port map (
            O => \N__67799\,
            I => \N__67757\
        );

    \I__16435\ : Span4Mux_h
    port map (
            O => \N__67796\,
            I => \N__67750\
        );

    \I__16434\ : LocalMux
    port map (
            O => \N__67793\,
            I => \N__67750\
        );

    \I__16433\ : Span4Mux_h
    port map (
            O => \N__67790\,
            I => \N__67750\
        );

    \I__16432\ : Span4Mux_h
    port map (
            O => \N__67785\,
            I => \N__67747\
        );

    \I__16431\ : Span4Mux_v
    port map (
            O => \N__67778\,
            I => \N__67744\
        );

    \I__16430\ : InMux
    port map (
            O => \N__67777\,
            I => \N__67741\
        );

    \I__16429\ : InMux
    port map (
            O => \N__67776\,
            I => \N__67738\
        );

    \I__16428\ : Span12Mux_h
    port map (
            O => \N__67773\,
            I => \N__67733\
        );

    \I__16427\ : Span12Mux_v
    port map (
            O => \N__67770\,
            I => \N__67733\
        );

    \I__16426\ : Span12Mux_v
    port map (
            O => \N__67763\,
            I => \N__67730\
        );

    \I__16425\ : LocalMux
    port map (
            O => \N__67760\,
            I => \N__67723\
        );

    \I__16424\ : Span4Mux_h
    port map (
            O => \N__67757\,
            I => \N__67723\
        );

    \I__16423\ : Span4Mux_v
    port map (
            O => \N__67750\,
            I => \N__67723\
        );

    \I__16422\ : Span4Mux_v
    port map (
            O => \N__67747\,
            I => \N__67718\
        );

    \I__16421\ : Span4Mux_h
    port map (
            O => \N__67744\,
            I => \N__67718\
        );

    \I__16420\ : LocalMux
    port map (
            O => \N__67741\,
            I => rx_data_5
        );

    \I__16419\ : LocalMux
    port map (
            O => \N__67738\,
            I => rx_data_5
        );

    \I__16418\ : Odrv12
    port map (
            O => \N__67733\,
            I => rx_data_5
        );

    \I__16417\ : Odrv12
    port map (
            O => \N__67730\,
            I => rx_data_5
        );

    \I__16416\ : Odrv4
    port map (
            O => \N__67723\,
            I => rx_data_5
        );

    \I__16415\ : Odrv4
    port map (
            O => \N__67718\,
            I => rx_data_5
        );

    \I__16414\ : CascadeMux
    port map (
            O => \N__67705\,
            I => \N__67701\
        );

    \I__16413\ : CascadeMux
    port map (
            O => \N__67704\,
            I => \N__67698\
        );

    \I__16412\ : InMux
    port map (
            O => \N__67701\,
            I => \N__67693\
        );

    \I__16411\ : InMux
    port map (
            O => \N__67698\,
            I => \N__67690\
        );

    \I__16410\ : InMux
    port map (
            O => \N__67697\,
            I => \N__67685\
        );

    \I__16409\ : InMux
    port map (
            O => \N__67696\,
            I => \N__67685\
        );

    \I__16408\ : LocalMux
    port map (
            O => \N__67693\,
            I => \N__67682\
        );

    \I__16407\ : LocalMux
    port map (
            O => \N__67690\,
            I => \c0.data_in_frame_20_2\
        );

    \I__16406\ : LocalMux
    port map (
            O => \N__67685\,
            I => \c0.data_in_frame_20_2\
        );

    \I__16405\ : Odrv4
    port map (
            O => \N__67682\,
            I => \c0.data_in_frame_20_2\
        );

    \I__16404\ : InMux
    port map (
            O => \N__67675\,
            I => \N__67670\
        );

    \I__16403\ : InMux
    port map (
            O => \N__67674\,
            I => \N__67667\
        );

    \I__16402\ : InMux
    port map (
            O => \N__67673\,
            I => \N__67663\
        );

    \I__16401\ : LocalMux
    port map (
            O => \N__67670\,
            I => \N__67658\
        );

    \I__16400\ : LocalMux
    port map (
            O => \N__67667\,
            I => \N__67658\
        );

    \I__16399\ : InMux
    port map (
            O => \N__67666\,
            I => \N__67654\
        );

    \I__16398\ : LocalMux
    port map (
            O => \N__67663\,
            I => \N__67649\
        );

    \I__16397\ : Span4Mux_v
    port map (
            O => \N__67658\,
            I => \N__67649\
        );

    \I__16396\ : InMux
    port map (
            O => \N__67657\,
            I => \N__67646\
        );

    \I__16395\ : LocalMux
    port map (
            O => \N__67654\,
            I => \c0.n20840\
        );

    \I__16394\ : Odrv4
    port map (
            O => \N__67649\,
            I => \c0.n20840\
        );

    \I__16393\ : LocalMux
    port map (
            O => \N__67646\,
            I => \c0.n20840\
        );

    \I__16392\ : InMux
    port map (
            O => \N__67639\,
            I => \N__67636\
        );

    \I__16391\ : LocalMux
    port map (
            O => \N__67636\,
            I => \N__67633\
        );

    \I__16390\ : Span4Mux_v
    port map (
            O => \N__67633\,
            I => \N__67630\
        );

    \I__16389\ : Span4Mux_h
    port map (
            O => \N__67630\,
            I => \N__67626\
        );

    \I__16388\ : InMux
    port map (
            O => \N__67629\,
            I => \N__67623\
        );

    \I__16387\ : Odrv4
    port map (
            O => \N__67626\,
            I => \c0.n22_adj_3322\
        );

    \I__16386\ : LocalMux
    port map (
            O => \N__67623\,
            I => \c0.n22_adj_3322\
        );

    \I__16385\ : InMux
    port map (
            O => \N__67618\,
            I => \N__67615\
        );

    \I__16384\ : LocalMux
    port map (
            O => \N__67615\,
            I => \N__67610\
        );

    \I__16383\ : InMux
    port map (
            O => \N__67614\,
            I => \N__67607\
        );

    \I__16382\ : InMux
    port map (
            O => \N__67613\,
            I => \N__67604\
        );

    \I__16381\ : Span4Mux_h
    port map (
            O => \N__67610\,
            I => \N__67601\
        );

    \I__16380\ : LocalMux
    port map (
            O => \N__67607\,
            I => \N__67598\
        );

    \I__16379\ : LocalMux
    port map (
            O => \N__67604\,
            I => \N__67595\
        );

    \I__16378\ : Span4Mux_v
    port map (
            O => \N__67601\,
            I => \N__67590\
        );

    \I__16377\ : Span4Mux_v
    port map (
            O => \N__67598\,
            I => \N__67590\
        );

    \I__16376\ : Span4Mux_h
    port map (
            O => \N__67595\,
            I => \N__67587\
        );

    \I__16375\ : Odrv4
    port map (
            O => \N__67590\,
            I => \c0.n11971\
        );

    \I__16374\ : Odrv4
    port map (
            O => \N__67587\,
            I => \c0.n11971\
        );

    \I__16373\ : InMux
    port map (
            O => \N__67582\,
            I => \N__67579\
        );

    \I__16372\ : LocalMux
    port map (
            O => \N__67579\,
            I => \c0.n19484\
        );

    \I__16371\ : CascadeMux
    port map (
            O => \N__67576\,
            I => \c0.n7_adj_3072_cascade_\
        );

    \I__16370\ : CascadeMux
    port map (
            O => \N__67573\,
            I => \c0.n18413_cascade_\
        );

    \I__16369\ : InMux
    port map (
            O => \N__67570\,
            I => \N__67567\
        );

    \I__16368\ : LocalMux
    port map (
            O => \N__67567\,
            I => \N__67563\
        );

    \I__16367\ : InMux
    port map (
            O => \N__67566\,
            I => \N__67559\
        );

    \I__16366\ : Span4Mux_v
    port map (
            O => \N__67563\,
            I => \N__67556\
        );

    \I__16365\ : CascadeMux
    port map (
            O => \N__67562\,
            I => \N__67553\
        );

    \I__16364\ : LocalMux
    port map (
            O => \N__67559\,
            I => \N__67550\
        );

    \I__16363\ : Span4Mux_h
    port map (
            O => \N__67556\,
            I => \N__67547\
        );

    \I__16362\ : InMux
    port map (
            O => \N__67553\,
            I => \N__67544\
        );

    \I__16361\ : Span4Mux_h
    port map (
            O => \N__67550\,
            I => \N__67541\
        );

    \I__16360\ : Span4Mux_h
    port map (
            O => \N__67547\,
            I => \N__67538\
        );

    \I__16359\ : LocalMux
    port map (
            O => \N__67544\,
            I => \c0.data_in_frame_26_3\
        );

    \I__16358\ : Odrv4
    port map (
            O => \N__67541\,
            I => \c0.data_in_frame_26_3\
        );

    \I__16357\ : Odrv4
    port map (
            O => \N__67538\,
            I => \c0.data_in_frame_26_3\
        );

    \I__16356\ : InMux
    port map (
            O => \N__67531\,
            I => \N__67523\
        );

    \I__16355\ : InMux
    port map (
            O => \N__67530\,
            I => \N__67519\
        );

    \I__16354\ : InMux
    port map (
            O => \N__67529\,
            I => \N__67516\
        );

    \I__16353\ : InMux
    port map (
            O => \N__67528\,
            I => \N__67511\
        );

    \I__16352\ : InMux
    port map (
            O => \N__67527\,
            I => \N__67511\
        );

    \I__16351\ : InMux
    port map (
            O => \N__67526\,
            I => \N__67508\
        );

    \I__16350\ : LocalMux
    port map (
            O => \N__67523\,
            I => \N__67505\
        );

    \I__16349\ : InMux
    port map (
            O => \N__67522\,
            I => \N__67501\
        );

    \I__16348\ : LocalMux
    port map (
            O => \N__67519\,
            I => \N__67498\
        );

    \I__16347\ : LocalMux
    port map (
            O => \N__67516\,
            I => \N__67495\
        );

    \I__16346\ : LocalMux
    port map (
            O => \N__67511\,
            I => \N__67492\
        );

    \I__16345\ : LocalMux
    port map (
            O => \N__67508\,
            I => \N__67489\
        );

    \I__16344\ : Span4Mux_h
    port map (
            O => \N__67505\,
            I => \N__67486\
        );

    \I__16343\ : InMux
    port map (
            O => \N__67504\,
            I => \N__67483\
        );

    \I__16342\ : LocalMux
    port map (
            O => \N__67501\,
            I => \N__67478\
        );

    \I__16341\ : Span4Mux_v
    port map (
            O => \N__67498\,
            I => \N__67478\
        );

    \I__16340\ : Span4Mux_v
    port map (
            O => \N__67495\,
            I => \N__67475\
        );

    \I__16339\ : Span4Mux_h
    port map (
            O => \N__67492\,
            I => \N__67472\
        );

    \I__16338\ : Span4Mux_h
    port map (
            O => \N__67489\,
            I => \N__67467\
        );

    \I__16337\ : Span4Mux_h
    port map (
            O => \N__67486\,
            I => \N__67467\
        );

    \I__16336\ : LocalMux
    port map (
            O => \N__67483\,
            I => \N__67462\
        );

    \I__16335\ : Span4Mux_v
    port map (
            O => \N__67478\,
            I => \N__67462\
        );

    \I__16334\ : Span4Mux_h
    port map (
            O => \N__67475\,
            I => \N__67459\
        );

    \I__16333\ : Span4Mux_h
    port map (
            O => \N__67472\,
            I => \N__67456\
        );

    \I__16332\ : Span4Mux_v
    port map (
            O => \N__67467\,
            I => \N__67453\
        );

    \I__16331\ : Span4Mux_h
    port map (
            O => \N__67462\,
            I => \N__67450\
        );

    \I__16330\ : Sp12to4
    port map (
            O => \N__67459\,
            I => \N__67447\
        );

    \I__16329\ : Odrv4
    port map (
            O => \N__67456\,
            I => n19127
        );

    \I__16328\ : Odrv4
    port map (
            O => \N__67453\,
            I => n19127
        );

    \I__16327\ : Odrv4
    port map (
            O => \N__67450\,
            I => n19127
        );

    \I__16326\ : Odrv12
    port map (
            O => \N__67447\,
            I => n19127
        );

    \I__16325\ : InMux
    port map (
            O => \N__67438\,
            I => \N__67435\
        );

    \I__16324\ : LocalMux
    port map (
            O => \N__67435\,
            I => \N__67431\
        );

    \I__16323\ : CascadeMux
    port map (
            O => \N__67434\,
            I => \N__67428\
        );

    \I__16322\ : Span4Mux_v
    port map (
            O => \N__67431\,
            I => \N__67424\
        );

    \I__16321\ : InMux
    port map (
            O => \N__67428\,
            I => \N__67421\
        );

    \I__16320\ : InMux
    port map (
            O => \N__67427\,
            I => \N__67418\
        );

    \I__16319\ : Sp12to4
    port map (
            O => \N__67424\,
            I => \N__67413\
        );

    \I__16318\ : LocalMux
    port map (
            O => \N__67421\,
            I => \N__67413\
        );

    \I__16317\ : LocalMux
    port map (
            O => \N__67418\,
            I => data_in_frame_22_5
        );

    \I__16316\ : Odrv12
    port map (
            O => \N__67413\,
            I => data_in_frame_22_5
        );

    \I__16315\ : InMux
    port map (
            O => \N__67408\,
            I => \N__67405\
        );

    \I__16314\ : LocalMux
    port map (
            O => \N__67405\,
            I => \N__67401\
        );

    \I__16313\ : InMux
    port map (
            O => \N__67404\,
            I => \N__67398\
        );

    \I__16312\ : Span4Mux_v
    port map (
            O => \N__67401\,
            I => \N__67393\
        );

    \I__16311\ : LocalMux
    port map (
            O => \N__67398\,
            I => \N__67393\
        );

    \I__16310\ : Span4Mux_h
    port map (
            O => \N__67393\,
            I => \N__67390\
        );

    \I__16309\ : Odrv4
    port map (
            O => \N__67390\,
            I => \c0.n9_adj_3069\
        );

    \I__16308\ : InMux
    port map (
            O => \N__67387\,
            I => \N__67383\
        );

    \I__16307\ : InMux
    port map (
            O => \N__67386\,
            I => \N__67380\
        );

    \I__16306\ : LocalMux
    port map (
            O => \N__67383\,
            I => \N__67373\
        );

    \I__16305\ : LocalMux
    port map (
            O => \N__67380\,
            I => \N__67373\
        );

    \I__16304\ : InMux
    port map (
            O => \N__67379\,
            I => \N__67368\
        );

    \I__16303\ : InMux
    port map (
            O => \N__67378\,
            I => \N__67368\
        );

    \I__16302\ : Span4Mux_v
    port map (
            O => \N__67373\,
            I => \N__67365\
        );

    \I__16301\ : LocalMux
    port map (
            O => \N__67368\,
            I => \c0.n20451\
        );

    \I__16300\ : Odrv4
    port map (
            O => \N__67365\,
            I => \c0.n20451\
        );

    \I__16299\ : InMux
    port map (
            O => \N__67360\,
            I => \N__67357\
        );

    \I__16298\ : LocalMux
    port map (
            O => \N__67357\,
            I => \c0.n8_adj_3070\
        );

    \I__16297\ : InMux
    port map (
            O => \N__67354\,
            I => \N__67351\
        );

    \I__16296\ : LocalMux
    port map (
            O => \N__67351\,
            I => \c0.n19315\
        );

    \I__16295\ : InMux
    port map (
            O => \N__67348\,
            I => \N__67345\
        );

    \I__16294\ : LocalMux
    port map (
            O => \N__67345\,
            I => \N__67342\
        );

    \I__16293\ : Span4Mux_v
    port map (
            O => \N__67342\,
            I => \N__67339\
        );

    \I__16292\ : Span4Mux_h
    port map (
            O => \N__67339\,
            I => \N__67336\
        );

    \I__16291\ : Span4Mux_v
    port map (
            O => \N__67336\,
            I => \N__67333\
        );

    \I__16290\ : Odrv4
    port map (
            O => \N__67333\,
            I => \c0.n26_adj_3550\
        );

    \I__16289\ : InMux
    port map (
            O => \N__67330\,
            I => \N__67327\
        );

    \I__16288\ : LocalMux
    port map (
            O => \N__67327\,
            I => \N__67324\
        );

    \I__16287\ : Span4Mux_h
    port map (
            O => \N__67324\,
            I => \N__67321\
        );

    \I__16286\ : Span4Mux_v
    port map (
            O => \N__67321\,
            I => \N__67318\
        );

    \I__16285\ : Odrv4
    port map (
            O => \N__67318\,
            I => \c0.n27_adj_3551\
        );

    \I__16284\ : CascadeMux
    port map (
            O => \N__67315\,
            I => \N__67312\
        );

    \I__16283\ : InMux
    port map (
            O => \N__67312\,
            I => \N__67309\
        );

    \I__16282\ : LocalMux
    port map (
            O => \N__67309\,
            I => \N__67306\
        );

    \I__16281\ : Odrv12
    port map (
            O => \N__67306\,
            I => \c0.n25_adj_3553\
        );

    \I__16280\ : InMux
    port map (
            O => \N__67303\,
            I => \N__67299\
        );

    \I__16279\ : InMux
    port map (
            O => \N__67302\,
            I => \N__67296\
        );

    \I__16278\ : LocalMux
    port map (
            O => \N__67299\,
            I => \N__67293\
        );

    \I__16277\ : LocalMux
    port map (
            O => \N__67296\,
            I => \N__67290\
        );

    \I__16276\ : Span4Mux_h
    port map (
            O => \N__67293\,
            I => \N__67285\
        );

    \I__16275\ : Span4Mux_h
    port map (
            O => \N__67290\,
            I => \N__67282\
        );

    \I__16274\ : InMux
    port map (
            O => \N__67289\,
            I => \N__67277\
        );

    \I__16273\ : InMux
    port map (
            O => \N__67288\,
            I => \N__67277\
        );

    \I__16272\ : Odrv4
    port map (
            O => \N__67285\,
            I => \c0.n49_adj_3358\
        );

    \I__16271\ : Odrv4
    port map (
            O => \N__67282\,
            I => \c0.n49_adj_3358\
        );

    \I__16270\ : LocalMux
    port map (
            O => \N__67277\,
            I => \c0.n49_adj_3358\
        );

    \I__16269\ : CascadeMux
    port map (
            O => \N__67270\,
            I => \N__67267\
        );

    \I__16268\ : InMux
    port map (
            O => \N__67267\,
            I => \N__67260\
        );

    \I__16267\ : InMux
    port map (
            O => \N__67266\,
            I => \N__67255\
        );

    \I__16266\ : InMux
    port map (
            O => \N__67265\,
            I => \N__67255\
        );

    \I__16265\ : InMux
    port map (
            O => \N__67264\,
            I => \N__67250\
        );

    \I__16264\ : InMux
    port map (
            O => \N__67263\,
            I => \N__67250\
        );

    \I__16263\ : LocalMux
    port map (
            O => \N__67260\,
            I => \c0.n17832\
        );

    \I__16262\ : LocalMux
    port map (
            O => \N__67255\,
            I => \c0.n17832\
        );

    \I__16261\ : LocalMux
    port map (
            O => \N__67250\,
            I => \c0.n17832\
        );

    \I__16260\ : InMux
    port map (
            O => \N__67243\,
            I => \N__67234\
        );

    \I__16259\ : InMux
    port map (
            O => \N__67242\,
            I => \N__67234\
        );

    \I__16258\ : InMux
    port map (
            O => \N__67241\,
            I => \N__67234\
        );

    \I__16257\ : LocalMux
    port map (
            O => \N__67234\,
            I => \c0.n40_adj_3271\
        );

    \I__16256\ : CascadeMux
    port map (
            O => \N__67231\,
            I => \N__67228\
        );

    \I__16255\ : InMux
    port map (
            O => \N__67228\,
            I => \N__67213\
        );

    \I__16254\ : InMux
    port map (
            O => \N__67227\,
            I => \N__67213\
        );

    \I__16253\ : InMux
    port map (
            O => \N__67226\,
            I => \N__67204\
        );

    \I__16252\ : InMux
    port map (
            O => \N__67225\,
            I => \N__67204\
        );

    \I__16251\ : InMux
    port map (
            O => \N__67224\,
            I => \N__67204\
        );

    \I__16250\ : InMux
    port map (
            O => \N__67223\,
            I => \N__67204\
        );

    \I__16249\ : CascadeMux
    port map (
            O => \N__67222\,
            I => \N__67201\
        );

    \I__16248\ : InMux
    port map (
            O => \N__67221\,
            I => \N__67191\
        );

    \I__16247\ : InMux
    port map (
            O => \N__67220\,
            I => \N__67191\
        );

    \I__16246\ : CascadeMux
    port map (
            O => \N__67219\,
            I => \N__67188\
        );

    \I__16245\ : InMux
    port map (
            O => \N__67218\,
            I => \N__67184\
        );

    \I__16244\ : LocalMux
    port map (
            O => \N__67213\,
            I => \N__67179\
        );

    \I__16243\ : LocalMux
    port map (
            O => \N__67204\,
            I => \N__67179\
        );

    \I__16242\ : InMux
    port map (
            O => \N__67201\,
            I => \N__67173\
        );

    \I__16241\ : InMux
    port map (
            O => \N__67200\,
            I => \N__67173\
        );

    \I__16240\ : InMux
    port map (
            O => \N__67199\,
            I => \N__67170\
        );

    \I__16239\ : InMux
    port map (
            O => \N__67198\,
            I => \N__67167\
        );

    \I__16238\ : InMux
    port map (
            O => \N__67197\,
            I => \N__67163\
        );

    \I__16237\ : InMux
    port map (
            O => \N__67196\,
            I => \N__67160\
        );

    \I__16236\ : LocalMux
    port map (
            O => \N__67191\,
            I => \N__67157\
        );

    \I__16235\ : InMux
    port map (
            O => \N__67188\,
            I => \N__67154\
        );

    \I__16234\ : InMux
    port map (
            O => \N__67187\,
            I => \N__67151\
        );

    \I__16233\ : LocalMux
    port map (
            O => \N__67184\,
            I => \N__67148\
        );

    \I__16232\ : Span4Mux_v
    port map (
            O => \N__67179\,
            I => \N__67145\
        );

    \I__16231\ : InMux
    port map (
            O => \N__67178\,
            I => \N__67141\
        );

    \I__16230\ : LocalMux
    port map (
            O => \N__67173\,
            I => \N__67138\
        );

    \I__16229\ : LocalMux
    port map (
            O => \N__67170\,
            I => \N__67135\
        );

    \I__16228\ : LocalMux
    port map (
            O => \N__67167\,
            I => \N__67132\
        );

    \I__16227\ : InMux
    port map (
            O => \N__67166\,
            I => \N__67127\
        );

    \I__16226\ : LocalMux
    port map (
            O => \N__67163\,
            I => \N__67122\
        );

    \I__16225\ : LocalMux
    port map (
            O => \N__67160\,
            I => \N__67122\
        );

    \I__16224\ : Span4Mux_h
    port map (
            O => \N__67157\,
            I => \N__67119\
        );

    \I__16223\ : LocalMux
    port map (
            O => \N__67154\,
            I => \N__67113\
        );

    \I__16222\ : LocalMux
    port map (
            O => \N__67151\,
            I => \N__67113\
        );

    \I__16221\ : Span4Mux_v
    port map (
            O => \N__67148\,
            I => \N__67108\
        );

    \I__16220\ : Span4Mux_h
    port map (
            O => \N__67145\,
            I => \N__67108\
        );

    \I__16219\ : InMux
    port map (
            O => \N__67144\,
            I => \N__67105\
        );

    \I__16218\ : LocalMux
    port map (
            O => \N__67141\,
            I => \N__67102\
        );

    \I__16217\ : Span4Mux_v
    port map (
            O => \N__67138\,
            I => \N__67095\
        );

    \I__16216\ : Span4Mux_v
    port map (
            O => \N__67135\,
            I => \N__67095\
        );

    \I__16215\ : Span4Mux_h
    port map (
            O => \N__67132\,
            I => \N__67095\
        );

    \I__16214\ : InMux
    port map (
            O => \N__67131\,
            I => \N__67092\
        );

    \I__16213\ : InMux
    port map (
            O => \N__67130\,
            I => \N__67089\
        );

    \I__16212\ : LocalMux
    port map (
            O => \N__67127\,
            I => \N__67086\
        );

    \I__16211\ : Span4Mux_v
    port map (
            O => \N__67122\,
            I => \N__67081\
        );

    \I__16210\ : Span4Mux_v
    port map (
            O => \N__67119\,
            I => \N__67081\
        );

    \I__16209\ : InMux
    port map (
            O => \N__67118\,
            I => \N__67078\
        );

    \I__16208\ : Span4Mux_h
    port map (
            O => \N__67113\,
            I => \N__67075\
        );

    \I__16207\ : Span4Mux_h
    port map (
            O => \N__67108\,
            I => \N__67072\
        );

    \I__16206\ : LocalMux
    port map (
            O => \N__67105\,
            I => \N__67065\
        );

    \I__16205\ : Span4Mux_h
    port map (
            O => \N__67102\,
            I => \N__67065\
        );

    \I__16204\ : Span4Mux_h
    port map (
            O => \N__67095\,
            I => \N__67065\
        );

    \I__16203\ : LocalMux
    port map (
            O => \N__67092\,
            I => \N__67062\
        );

    \I__16202\ : LocalMux
    port map (
            O => \N__67089\,
            I => \N__67057\
        );

    \I__16201\ : Span4Mux_v
    port map (
            O => \N__67086\,
            I => \N__67057\
        );

    \I__16200\ : Span4Mux_h
    port map (
            O => \N__67081\,
            I => \N__67054\
        );

    \I__16199\ : LocalMux
    port map (
            O => \N__67078\,
            I => \N__67051\
        );

    \I__16198\ : Span4Mux_h
    port map (
            O => \N__67075\,
            I => \N__67044\
        );

    \I__16197\ : Span4Mux_h
    port map (
            O => \N__67072\,
            I => \N__67044\
        );

    \I__16196\ : Span4Mux_v
    port map (
            O => \N__67065\,
            I => \N__67044\
        );

    \I__16195\ : Span4Mux_h
    port map (
            O => \N__67062\,
            I => \N__67041\
        );

    \I__16194\ : Span4Mux_v
    port map (
            O => \N__67057\,
            I => \N__67038\
        );

    \I__16193\ : Sp12to4
    port map (
            O => \N__67054\,
            I => \N__67035\
        );

    \I__16192\ : Span4Mux_v
    port map (
            O => \N__67051\,
            I => \N__67030\
        );

    \I__16191\ : Span4Mux_v
    port map (
            O => \N__67044\,
            I => \N__67030\
        );

    \I__16190\ : Odrv4
    port map (
            O => \N__67041\,
            I => \c0.n19111\
        );

    \I__16189\ : Odrv4
    port map (
            O => \N__67038\,
            I => \c0.n19111\
        );

    \I__16188\ : Odrv12
    port map (
            O => \N__67035\,
            I => \c0.n19111\
        );

    \I__16187\ : Odrv4
    port map (
            O => \N__67030\,
            I => \c0.n19111\
        );

    \I__16186\ : CascadeMux
    port map (
            O => \N__67021\,
            I => \N__67017\
        );

    \I__16185\ : CascadeMux
    port map (
            O => \N__67020\,
            I => \N__67014\
        );

    \I__16184\ : InMux
    port map (
            O => \N__67017\,
            I => \N__67011\
        );

    \I__16183\ : InMux
    port map (
            O => \N__67014\,
            I => \N__67008\
        );

    \I__16182\ : LocalMux
    port map (
            O => \N__67011\,
            I => \N__67005\
        );

    \I__16181\ : LocalMux
    port map (
            O => \N__67008\,
            I => \N__67002\
        );

    \I__16180\ : Span4Mux_v
    port map (
            O => \N__67005\,
            I => \N__66999\
        );

    \I__16179\ : Span4Mux_h
    port map (
            O => \N__67002\,
            I => \N__66994\
        );

    \I__16178\ : Span4Mux_v
    port map (
            O => \N__66999\,
            I => \N__66994\
        );

    \I__16177\ : Span4Mux_h
    port map (
            O => \N__66994\,
            I => \N__66991\
        );

    \I__16176\ : Odrv4
    port map (
            O => \N__66991\,
            I => \c0.data_in_frame_29_3\
        );

    \I__16175\ : CascadeMux
    port map (
            O => \N__66988\,
            I => \N__66984\
        );

    \I__16174\ : CascadeMux
    port map (
            O => \N__66987\,
            I => \N__66981\
        );

    \I__16173\ : InMux
    port map (
            O => \N__66984\,
            I => \N__66963\
        );

    \I__16172\ : InMux
    port map (
            O => \N__66981\,
            I => \N__66963\
        );

    \I__16171\ : InMux
    port map (
            O => \N__66980\,
            I => \N__66963\
        );

    \I__16170\ : InMux
    port map (
            O => \N__66979\,
            I => \N__66963\
        );

    \I__16169\ : CascadeMux
    port map (
            O => \N__66978\,
            I => \N__66959\
        );

    \I__16168\ : CascadeMux
    port map (
            O => \N__66977\,
            I => \N__66949\
        );

    \I__16167\ : CascadeMux
    port map (
            O => \N__66976\,
            I => \N__66944\
        );

    \I__16166\ : CascadeMux
    port map (
            O => \N__66975\,
            I => \N__66938\
        );

    \I__16165\ : CascadeMux
    port map (
            O => \N__66974\,
            I => \N__66935\
        );

    \I__16164\ : InMux
    port map (
            O => \N__66973\,
            I => \N__66928\
        );

    \I__16163\ : InMux
    port map (
            O => \N__66972\,
            I => \N__66928\
        );

    \I__16162\ : LocalMux
    port map (
            O => \N__66963\,
            I => \N__66925\
        );

    \I__16161\ : InMux
    port map (
            O => \N__66962\,
            I => \N__66918\
        );

    \I__16160\ : InMux
    port map (
            O => \N__66959\,
            I => \N__66918\
        );

    \I__16159\ : CascadeMux
    port map (
            O => \N__66958\,
            I => \N__66913\
        );

    \I__16158\ : InMux
    port map (
            O => \N__66957\,
            I => \N__66909\
        );

    \I__16157\ : InMux
    port map (
            O => \N__66956\,
            I => \N__66900\
        );

    \I__16156\ : InMux
    port map (
            O => \N__66955\,
            I => \N__66900\
        );

    \I__16155\ : InMux
    port map (
            O => \N__66954\,
            I => \N__66900\
        );

    \I__16154\ : InMux
    port map (
            O => \N__66953\,
            I => \N__66900\
        );

    \I__16153\ : InMux
    port map (
            O => \N__66952\,
            I => \N__66889\
        );

    \I__16152\ : InMux
    port map (
            O => \N__66949\,
            I => \N__66889\
        );

    \I__16151\ : InMux
    port map (
            O => \N__66948\,
            I => \N__66889\
        );

    \I__16150\ : InMux
    port map (
            O => \N__66947\,
            I => \N__66882\
        );

    \I__16149\ : InMux
    port map (
            O => \N__66944\,
            I => \N__66882\
        );

    \I__16148\ : InMux
    port map (
            O => \N__66943\,
            I => \N__66882\
        );

    \I__16147\ : InMux
    port map (
            O => \N__66942\,
            I => \N__66868\
        );

    \I__16146\ : InMux
    port map (
            O => \N__66941\,
            I => \N__66868\
        );

    \I__16145\ : InMux
    port map (
            O => \N__66938\,
            I => \N__66868\
        );

    \I__16144\ : InMux
    port map (
            O => \N__66935\,
            I => \N__66868\
        );

    \I__16143\ : InMux
    port map (
            O => \N__66934\,
            I => \N__66868\
        );

    \I__16142\ : InMux
    port map (
            O => \N__66933\,
            I => \N__66865\
        );

    \I__16141\ : LocalMux
    port map (
            O => \N__66928\,
            I => \N__66860\
        );

    \I__16140\ : Span4Mux_v
    port map (
            O => \N__66925\,
            I => \N__66860\
        );

    \I__16139\ : InMux
    port map (
            O => \N__66924\,
            I => \N__66857\
        );

    \I__16138\ : InMux
    port map (
            O => \N__66923\,
            I => \N__66854\
        );

    \I__16137\ : LocalMux
    port map (
            O => \N__66918\,
            I => \N__66851\
        );

    \I__16136\ : InMux
    port map (
            O => \N__66917\,
            I => \N__66846\
        );

    \I__16135\ : InMux
    port map (
            O => \N__66916\,
            I => \N__66841\
        );

    \I__16134\ : InMux
    port map (
            O => \N__66913\,
            I => \N__66841\
        );

    \I__16133\ : InMux
    port map (
            O => \N__66912\,
            I => \N__66838\
        );

    \I__16132\ : LocalMux
    port map (
            O => \N__66909\,
            I => \N__66835\
        );

    \I__16131\ : LocalMux
    port map (
            O => \N__66900\,
            I => \N__66832\
        );

    \I__16130\ : InMux
    port map (
            O => \N__66899\,
            I => \N__66829\
        );

    \I__16129\ : InMux
    port map (
            O => \N__66898\,
            I => \N__66826\
        );

    \I__16128\ : InMux
    port map (
            O => \N__66897\,
            I => \N__66821\
        );

    \I__16127\ : InMux
    port map (
            O => \N__66896\,
            I => \N__66821\
        );

    \I__16126\ : LocalMux
    port map (
            O => \N__66889\,
            I => \N__66816\
        );

    \I__16125\ : LocalMux
    port map (
            O => \N__66882\,
            I => \N__66816\
        );

    \I__16124\ : InMux
    port map (
            O => \N__66881\,
            I => \N__66809\
        );

    \I__16123\ : InMux
    port map (
            O => \N__66880\,
            I => \N__66809\
        );

    \I__16122\ : InMux
    port map (
            O => \N__66879\,
            I => \N__66809\
        );

    \I__16121\ : LocalMux
    port map (
            O => \N__66868\,
            I => \N__66806\
        );

    \I__16120\ : LocalMux
    port map (
            O => \N__66865\,
            I => \N__66799\
        );

    \I__16119\ : Span4Mux_h
    port map (
            O => \N__66860\,
            I => \N__66799\
        );

    \I__16118\ : LocalMux
    port map (
            O => \N__66857\,
            I => \N__66799\
        );

    \I__16117\ : LocalMux
    port map (
            O => \N__66854\,
            I => \N__66794\
        );

    \I__16116\ : Span4Mux_v
    port map (
            O => \N__66851\,
            I => \N__66794\
        );

    \I__16115\ : CascadeMux
    port map (
            O => \N__66850\,
            I => \N__66791\
        );

    \I__16114\ : InMux
    port map (
            O => \N__66849\,
            I => \N__66788\
        );

    \I__16113\ : LocalMux
    port map (
            O => \N__66846\,
            I => \N__66785\
        );

    \I__16112\ : LocalMux
    port map (
            O => \N__66841\,
            I => \N__66782\
        );

    \I__16111\ : LocalMux
    port map (
            O => \N__66838\,
            I => \N__66777\
        );

    \I__16110\ : Span4Mux_h
    port map (
            O => \N__66835\,
            I => \N__66777\
        );

    \I__16109\ : Span4Mux_v
    port map (
            O => \N__66832\,
            I => \N__66774\
        );

    \I__16108\ : LocalMux
    port map (
            O => \N__66829\,
            I => \N__66771\
        );

    \I__16107\ : LocalMux
    port map (
            O => \N__66826\,
            I => \N__66768\
        );

    \I__16106\ : LocalMux
    port map (
            O => \N__66821\,
            I => \N__66761\
        );

    \I__16105\ : Span4Mux_v
    port map (
            O => \N__66816\,
            I => \N__66761\
        );

    \I__16104\ : LocalMux
    port map (
            O => \N__66809\,
            I => \N__66761\
        );

    \I__16103\ : Span4Mux_v
    port map (
            O => \N__66806\,
            I => \N__66758\
        );

    \I__16102\ : Span4Mux_h
    port map (
            O => \N__66799\,
            I => \N__66755\
        );

    \I__16101\ : Sp12to4
    port map (
            O => \N__66794\,
            I => \N__66751\
        );

    \I__16100\ : InMux
    port map (
            O => \N__66791\,
            I => \N__66748\
        );

    \I__16099\ : LocalMux
    port map (
            O => \N__66788\,
            I => \N__66739\
        );

    \I__16098\ : Span4Mux_v
    port map (
            O => \N__66785\,
            I => \N__66739\
        );

    \I__16097\ : Span4Mux_h
    port map (
            O => \N__66782\,
            I => \N__66739\
        );

    \I__16096\ : Span4Mux_h
    port map (
            O => \N__66777\,
            I => \N__66739\
        );

    \I__16095\ : Span4Mux_h
    port map (
            O => \N__66774\,
            I => \N__66732\
        );

    \I__16094\ : Span4Mux_v
    port map (
            O => \N__66771\,
            I => \N__66732\
        );

    \I__16093\ : Span4Mux_h
    port map (
            O => \N__66768\,
            I => \N__66732\
        );

    \I__16092\ : Span4Mux_v
    port map (
            O => \N__66761\,
            I => \N__66729\
        );

    \I__16091\ : Span4Mux_h
    port map (
            O => \N__66758\,
            I => \N__66724\
        );

    \I__16090\ : Span4Mux_v
    port map (
            O => \N__66755\,
            I => \N__66724\
        );

    \I__16089\ : InMux
    port map (
            O => \N__66754\,
            I => \N__66721\
        );

    \I__16088\ : Span12Mux_v
    port map (
            O => \N__66751\,
            I => \N__66718\
        );

    \I__16087\ : LocalMux
    port map (
            O => \N__66748\,
            I => \N__66711\
        );

    \I__16086\ : Span4Mux_v
    port map (
            O => \N__66739\,
            I => \N__66711\
        );

    \I__16085\ : Span4Mux_h
    port map (
            O => \N__66732\,
            I => \N__66711\
        );

    \I__16084\ : Span4Mux_h
    port map (
            O => \N__66729\,
            I => \N__66708\
        );

    \I__16083\ : Span4Mux_v
    port map (
            O => \N__66724\,
            I => \N__66705\
        );

    \I__16082\ : LocalMux
    port map (
            O => \N__66721\,
            I => \c0.n12_adj_3006\
        );

    \I__16081\ : Odrv12
    port map (
            O => \N__66718\,
            I => \c0.n12_adj_3006\
        );

    \I__16080\ : Odrv4
    port map (
            O => \N__66711\,
            I => \c0.n12_adj_3006\
        );

    \I__16079\ : Odrv4
    port map (
            O => \N__66708\,
            I => \c0.n12_adj_3006\
        );

    \I__16078\ : Odrv4
    port map (
            O => \N__66705\,
            I => \c0.n12_adj_3006\
        );

    \I__16077\ : CascadeMux
    port map (
            O => \N__66694\,
            I => \N__66691\
        );

    \I__16076\ : InMux
    port map (
            O => \N__66691\,
            I => \N__66687\
        );

    \I__16075\ : InMux
    port map (
            O => \N__66690\,
            I => \N__66684\
        );

    \I__16074\ : LocalMux
    port map (
            O => \N__66687\,
            I => \N__66681\
        );

    \I__16073\ : LocalMux
    port map (
            O => \N__66684\,
            I => \N__66676\
        );

    \I__16072\ : Span12Mux_h
    port map (
            O => \N__66681\,
            I => \N__66676\
        );

    \I__16071\ : Odrv12
    port map (
            O => \N__66676\,
            I => \c0.data_in_frame_29_5\
        );

    \I__16070\ : InMux
    port map (
            O => \N__66673\,
            I => \N__66670\
        );

    \I__16069\ : LocalMux
    port map (
            O => \N__66670\,
            I => \N__66667\
        );

    \I__16068\ : Span4Mux_h
    port map (
            O => \N__66667\,
            I => \N__66664\
        );

    \I__16067\ : Odrv4
    port map (
            O => \N__66664\,
            I => \c0.n15_adj_3432\
        );

    \I__16066\ : InMux
    port map (
            O => \N__66661\,
            I => \N__66658\
        );

    \I__16065\ : LocalMux
    port map (
            O => \N__66658\,
            I => \N__66655\
        );

    \I__16064\ : Span4Mux_v
    port map (
            O => \N__66655\,
            I => \N__66652\
        );

    \I__16063\ : Odrv4
    port map (
            O => \N__66652\,
            I => \c0.n20503\
        );

    \I__16062\ : CascadeMux
    port map (
            O => \N__66649\,
            I => \N__66644\
        );

    \I__16061\ : InMux
    port map (
            O => \N__66648\,
            I => \N__66641\
        );

    \I__16060\ : InMux
    port map (
            O => \N__66647\,
            I => \N__66636\
        );

    \I__16059\ : InMux
    port map (
            O => \N__66644\,
            I => \N__66636\
        );

    \I__16058\ : LocalMux
    port map (
            O => \N__66641\,
            I => \N__66633\
        );

    \I__16057\ : LocalMux
    port map (
            O => \N__66636\,
            I => \N__66628\
        );

    \I__16056\ : Span4Mux_h
    port map (
            O => \N__66633\,
            I => \N__66625\
        );

    \I__16055\ : InMux
    port map (
            O => \N__66632\,
            I => \N__66622\
        );

    \I__16054\ : InMux
    port map (
            O => \N__66631\,
            I => \N__66619\
        );

    \I__16053\ : Span12Mux_s10_v
    port map (
            O => \N__66628\,
            I => \N__66616\
        );

    \I__16052\ : Span4Mux_h
    port map (
            O => \N__66625\,
            I => \N__66613\
        );

    \I__16051\ : LocalMux
    port map (
            O => \N__66622\,
            I => data_in_frame_23_1
        );

    \I__16050\ : LocalMux
    port map (
            O => \N__66619\,
            I => data_in_frame_23_1
        );

    \I__16049\ : Odrv12
    port map (
            O => \N__66616\,
            I => data_in_frame_23_1
        );

    \I__16048\ : Odrv4
    port map (
            O => \N__66613\,
            I => data_in_frame_23_1
        );

    \I__16047\ : CascadeMux
    port map (
            O => \N__66604\,
            I => \c0.n20503_cascade_\
        );

    \I__16046\ : InMux
    port map (
            O => \N__66601\,
            I => \N__66598\
        );

    \I__16045\ : LocalMux
    port map (
            O => \N__66598\,
            I => \N__66595\
        );

    \I__16044\ : Span12Mux_h
    port map (
            O => \N__66595\,
            I => \N__66592\
        );

    \I__16043\ : Odrv12
    port map (
            O => \N__66592\,
            I => \c0.n12_adj_3494\
        );

    \I__16042\ : InMux
    port map (
            O => \N__66589\,
            I => \N__66586\
        );

    \I__16041\ : LocalMux
    port map (
            O => \N__66586\,
            I => \N__66583\
        );

    \I__16040\ : Span4Mux_v
    port map (
            O => \N__66583\,
            I => \N__66579\
        );

    \I__16039\ : InMux
    port map (
            O => \N__66582\,
            I => \N__66576\
        );

    \I__16038\ : Odrv4
    port map (
            O => \N__66579\,
            I => \c0.n27_adj_3399\
        );

    \I__16037\ : LocalMux
    port map (
            O => \N__66576\,
            I => \c0.n27_adj_3399\
        );

    \I__16036\ : InMux
    port map (
            O => \N__66571\,
            I => \N__66567\
        );

    \I__16035\ : InMux
    port map (
            O => \N__66570\,
            I => \N__66564\
        );

    \I__16034\ : LocalMux
    port map (
            O => \N__66567\,
            I => \c0.data_in_frame_28_3\
        );

    \I__16033\ : LocalMux
    port map (
            O => \N__66564\,
            I => \c0.data_in_frame_28_3\
        );

    \I__16032\ : CascadeMux
    port map (
            O => \N__66559\,
            I => \c0.n27_adj_3399_cascade_\
        );

    \I__16031\ : InMux
    port map (
            O => \N__66556\,
            I => \N__66553\
        );

    \I__16030\ : LocalMux
    port map (
            O => \N__66553\,
            I => \N__66550\
        );

    \I__16029\ : Span4Mux_h
    port map (
            O => \N__66550\,
            I => \N__66547\
        );

    \I__16028\ : Span4Mux_v
    port map (
            O => \N__66547\,
            I => \N__66542\
        );

    \I__16027\ : InMux
    port map (
            O => \N__66546\,
            I => \N__66537\
        );

    \I__16026\ : InMux
    port map (
            O => \N__66545\,
            I => \N__66537\
        );

    \I__16025\ : Odrv4
    port map (
            O => \N__66542\,
            I => \c0.data_in_frame_26_1\
        );

    \I__16024\ : LocalMux
    port map (
            O => \N__66537\,
            I => \c0.data_in_frame_26_1\
        );

    \I__16023\ : CascadeMux
    port map (
            O => \N__66532\,
            I => \N__66529\
        );

    \I__16022\ : InMux
    port map (
            O => \N__66529\,
            I => \N__66526\
        );

    \I__16021\ : LocalMux
    port map (
            O => \N__66526\,
            I => \N__66523\
        );

    \I__16020\ : Span4Mux_h
    port map (
            O => \N__66523\,
            I => \N__66520\
        );

    \I__16019\ : Span4Mux_h
    port map (
            O => \N__66520\,
            I => \N__66517\
        );

    \I__16018\ : Odrv4
    port map (
            O => \N__66517\,
            I => \c0.n78_adj_3414\
        );

    \I__16017\ : CascadeMux
    port map (
            O => \N__66514\,
            I => \N__66511\
        );

    \I__16016\ : InMux
    port map (
            O => \N__66511\,
            I => \N__66507\
        );

    \I__16015\ : InMux
    port map (
            O => \N__66510\,
            I => \N__66504\
        );

    \I__16014\ : LocalMux
    port map (
            O => \N__66507\,
            I => \N__66501\
        );

    \I__16013\ : LocalMux
    port map (
            O => \N__66504\,
            I => \N__66497\
        );

    \I__16012\ : Span4Mux_h
    port map (
            O => \N__66501\,
            I => \N__66493\
        );

    \I__16011\ : InMux
    port map (
            O => \N__66500\,
            I => \N__66490\
        );

    \I__16010\ : Span4Mux_h
    port map (
            O => \N__66497\,
            I => \N__66487\
        );

    \I__16009\ : InMux
    port map (
            O => \N__66496\,
            I => \N__66484\
        );

    \I__16008\ : Span4Mux_h
    port map (
            O => \N__66493\,
            I => \N__66481\
        );

    \I__16007\ : LocalMux
    port map (
            O => \N__66490\,
            I => \N__66476\
        );

    \I__16006\ : Span4Mux_h
    port map (
            O => \N__66487\,
            I => \N__66476\
        );

    \I__16005\ : LocalMux
    port map (
            O => \N__66484\,
            I => data_in_frame_23_6
        );

    \I__16004\ : Odrv4
    port map (
            O => \N__66481\,
            I => data_in_frame_23_6
        );

    \I__16003\ : Odrv4
    port map (
            O => \N__66476\,
            I => data_in_frame_23_6
        );

    \I__16002\ : InMux
    port map (
            O => \N__66469\,
            I => \N__66466\
        );

    \I__16001\ : LocalMux
    port map (
            O => \N__66466\,
            I => \N__66461\
        );

    \I__16000\ : InMux
    port map (
            O => \N__66465\,
            I => \N__66458\
        );

    \I__15999\ : InMux
    port map (
            O => \N__66464\,
            I => \N__66455\
        );

    \I__15998\ : Span4Mux_v
    port map (
            O => \N__66461\,
            I => \N__66448\
        );

    \I__15997\ : LocalMux
    port map (
            O => \N__66458\,
            I => \N__66448\
        );

    \I__15996\ : LocalMux
    port map (
            O => \N__66455\,
            I => \N__66445\
        );

    \I__15995\ : InMux
    port map (
            O => \N__66454\,
            I => \N__66440\
        );

    \I__15994\ : InMux
    port map (
            O => \N__66453\,
            I => \N__66440\
        );

    \I__15993\ : Span4Mux_h
    port map (
            O => \N__66448\,
            I => \N__66437\
        );

    \I__15992\ : Span12Mux_s10_h
    port map (
            O => \N__66445\,
            I => \N__66434\
        );

    \I__15991\ : LocalMux
    port map (
            O => \N__66440\,
            I => data_in_frame_23_5
        );

    \I__15990\ : Odrv4
    port map (
            O => \N__66437\,
            I => data_in_frame_23_5
        );

    \I__15989\ : Odrv12
    port map (
            O => \N__66434\,
            I => data_in_frame_23_5
        );

    \I__15988\ : InMux
    port map (
            O => \N__66427\,
            I => \N__66424\
        );

    \I__15987\ : LocalMux
    port map (
            O => \N__66424\,
            I => \c0.n19487\
        );

    \I__15986\ : CascadeMux
    port map (
            O => \N__66421\,
            I => \N__66418\
        );

    \I__15985\ : InMux
    port map (
            O => \N__66418\,
            I => \N__66411\
        );

    \I__15984\ : InMux
    port map (
            O => \N__66417\,
            I => \N__66411\
        );

    \I__15983\ : InMux
    port map (
            O => \N__66416\,
            I => \N__66408\
        );

    \I__15982\ : LocalMux
    port map (
            O => \N__66411\,
            I => \N__66405\
        );

    \I__15981\ : LocalMux
    port map (
            O => \N__66408\,
            I => \N__66402\
        );

    \I__15980\ : Span4Mux_h
    port map (
            O => \N__66405\,
            I => \N__66397\
        );

    \I__15979\ : Span4Mux_h
    port map (
            O => \N__66402\,
            I => \N__66397\
        );

    \I__15978\ : Span4Mux_v
    port map (
            O => \N__66397\,
            I => \N__66392\
        );

    \I__15977\ : InMux
    port map (
            O => \N__66396\,
            I => \N__66387\
        );

    \I__15976\ : InMux
    port map (
            O => \N__66395\,
            I => \N__66387\
        );

    \I__15975\ : Odrv4
    port map (
            O => \N__66392\,
            I => data_in_frame_23_7
        );

    \I__15974\ : LocalMux
    port map (
            O => \N__66387\,
            I => data_in_frame_23_7
        );

    \I__15973\ : InMux
    port map (
            O => \N__66382\,
            I => \N__66378\
        );

    \I__15972\ : InMux
    port map (
            O => \N__66381\,
            I => \N__66375\
        );

    \I__15971\ : LocalMux
    port map (
            O => \N__66378\,
            I => \N__66370\
        );

    \I__15970\ : LocalMux
    port map (
            O => \N__66375\,
            I => \N__66370\
        );

    \I__15969\ : Span4Mux_v
    port map (
            O => \N__66370\,
            I => \N__66367\
        );

    \I__15968\ : Span4Mux_h
    port map (
            O => \N__66367\,
            I => \N__66364\
        );

    \I__15967\ : Odrv4
    port map (
            O => \N__66364\,
            I => \c0.n19251\
        );

    \I__15966\ : InMux
    port map (
            O => \N__66361\,
            I => \N__66358\
        );

    \I__15965\ : LocalMux
    port map (
            O => \N__66358\,
            I => \N__66355\
        );

    \I__15964\ : Span4Mux_v
    port map (
            O => \N__66355\,
            I => \N__66351\
        );

    \I__15963\ : InMux
    port map (
            O => \N__66354\,
            I => \N__66348\
        );

    \I__15962\ : Span4Mux_v
    port map (
            O => \N__66351\,
            I => \N__66345\
        );

    \I__15961\ : LocalMux
    port map (
            O => \N__66348\,
            I => \N__66342\
        );

    \I__15960\ : Odrv4
    port map (
            O => \N__66345\,
            I => \c0.n7_adj_3347\
        );

    \I__15959\ : Odrv12
    port map (
            O => \N__66342\,
            I => \c0.n7_adj_3347\
        );

    \I__15958\ : InMux
    port map (
            O => \N__66337\,
            I => \N__66333\
        );

    \I__15957\ : CascadeMux
    port map (
            O => \N__66336\,
            I => \N__66330\
        );

    \I__15956\ : LocalMux
    port map (
            O => \N__66333\,
            I => \N__66327\
        );

    \I__15955\ : InMux
    port map (
            O => \N__66330\,
            I => \N__66323\
        );

    \I__15954\ : Span4Mux_v
    port map (
            O => \N__66327\,
            I => \N__66320\
        );

    \I__15953\ : InMux
    port map (
            O => \N__66326\,
            I => \N__66317\
        );

    \I__15952\ : LocalMux
    port map (
            O => \N__66323\,
            I => \c0.data_in_frame_10_6\
        );

    \I__15951\ : Odrv4
    port map (
            O => \N__66320\,
            I => \c0.data_in_frame_10_6\
        );

    \I__15950\ : LocalMux
    port map (
            O => \N__66317\,
            I => \c0.data_in_frame_10_6\
        );

    \I__15949\ : CascadeMux
    port map (
            O => \N__66310\,
            I => \N__66307\
        );

    \I__15948\ : InMux
    port map (
            O => \N__66307\,
            I => \N__66304\
        );

    \I__15947\ : LocalMux
    port map (
            O => \N__66304\,
            I => \N__66301\
        );

    \I__15946\ : Odrv4
    port map (
            O => \N__66301\,
            I => \c0.n19359\
        );

    \I__15945\ : InMux
    port map (
            O => \N__66298\,
            I => \N__66295\
        );

    \I__15944\ : LocalMux
    port map (
            O => \N__66295\,
            I => \N__66291\
        );

    \I__15943\ : InMux
    port map (
            O => \N__66294\,
            I => \N__66288\
        );

    \I__15942\ : Span4Mux_v
    port map (
            O => \N__66291\,
            I => \N__66281\
        );

    \I__15941\ : LocalMux
    port map (
            O => \N__66288\,
            I => \N__66281\
        );

    \I__15940\ : InMux
    port map (
            O => \N__66287\,
            I => \N__66278\
        );

    \I__15939\ : CascadeMux
    port map (
            O => \N__66286\,
            I => \N__66275\
        );

    \I__15938\ : Span4Mux_h
    port map (
            O => \N__66281\,
            I => \N__66272\
        );

    \I__15937\ : LocalMux
    port map (
            O => \N__66278\,
            I => \N__66269\
        );

    \I__15936\ : InMux
    port map (
            O => \N__66275\,
            I => \N__66266\
        );

    \I__15935\ : Span4Mux_v
    port map (
            O => \N__66272\,
            I => \N__66261\
        );

    \I__15934\ : Span4Mux_v
    port map (
            O => \N__66269\,
            I => \N__66261\
        );

    \I__15933\ : LocalMux
    port map (
            O => \N__66266\,
            I => \c0.data_in_frame_12_6\
        );

    \I__15932\ : Odrv4
    port map (
            O => \N__66261\,
            I => \c0.data_in_frame_12_6\
        );

    \I__15931\ : InMux
    port map (
            O => \N__66256\,
            I => \N__66253\
        );

    \I__15930\ : LocalMux
    port map (
            O => \N__66253\,
            I => \N__66250\
        );

    \I__15929\ : Span4Mux_v
    port map (
            O => \N__66250\,
            I => \N__66247\
        );

    \I__15928\ : Odrv4
    port map (
            O => \N__66247\,
            I => \c0.n22_adj_3535\
        );

    \I__15927\ : InMux
    port map (
            O => \N__66244\,
            I => \N__66240\
        );

    \I__15926\ : InMux
    port map (
            O => \N__66243\,
            I => \N__66236\
        );

    \I__15925\ : LocalMux
    port map (
            O => \N__66240\,
            I => \N__66233\
        );

    \I__15924\ : CascadeMux
    port map (
            O => \N__66239\,
            I => \N__66230\
        );

    \I__15923\ : LocalMux
    port map (
            O => \N__66236\,
            I => \N__66227\
        );

    \I__15922\ : Span4Mux_h
    port map (
            O => \N__66233\,
            I => \N__66224\
        );

    \I__15921\ : InMux
    port map (
            O => \N__66230\,
            I => \N__66221\
        );

    \I__15920\ : Sp12to4
    port map (
            O => \N__66227\,
            I => \N__66216\
        );

    \I__15919\ : Sp12to4
    port map (
            O => \N__66224\,
            I => \N__66216\
        );

    \I__15918\ : LocalMux
    port map (
            O => \N__66221\,
            I => \c0.data_in_frame_20_1\
        );

    \I__15917\ : Odrv12
    port map (
            O => \N__66216\,
            I => \c0.data_in_frame_20_1\
        );

    \I__15916\ : CascadeMux
    port map (
            O => \N__66211\,
            I => \N__66206\
        );

    \I__15915\ : InMux
    port map (
            O => \N__66210\,
            I => \N__66198\
        );

    \I__15914\ : InMux
    port map (
            O => \N__66209\,
            I => \N__66198\
        );

    \I__15913\ : InMux
    port map (
            O => \N__66206\,
            I => \N__66195\
        );

    \I__15912\ : CascadeMux
    port map (
            O => \N__66205\,
            I => \N__66190\
        );

    \I__15911\ : CascadeMux
    port map (
            O => \N__66204\,
            I => \N__66181\
        );

    \I__15910\ : CascadeMux
    port map (
            O => \N__66203\,
            I => \N__66178\
        );

    \I__15909\ : LocalMux
    port map (
            O => \N__66198\,
            I => \N__66172\
        );

    \I__15908\ : LocalMux
    port map (
            O => \N__66195\,
            I => \N__66172\
        );

    \I__15907\ : InMux
    port map (
            O => \N__66194\,
            I => \N__66169\
        );

    \I__15906\ : InMux
    port map (
            O => \N__66193\,
            I => \N__66166\
        );

    \I__15905\ : InMux
    port map (
            O => \N__66190\,
            I => \N__66163\
        );

    \I__15904\ : CascadeMux
    port map (
            O => \N__66189\,
            I => \N__66159\
        );

    \I__15903\ : CascadeMux
    port map (
            O => \N__66188\,
            I => \N__66150\
        );

    \I__15902\ : CascadeMux
    port map (
            O => \N__66187\,
            I => \N__66147\
        );

    \I__15901\ : CascadeMux
    port map (
            O => \N__66186\,
            I => \N__66141\
        );

    \I__15900\ : InMux
    port map (
            O => \N__66185\,
            I => \N__66136\
        );

    \I__15899\ : InMux
    port map (
            O => \N__66184\,
            I => \N__66133\
        );

    \I__15898\ : InMux
    port map (
            O => \N__66181\,
            I => \N__66126\
        );

    \I__15897\ : InMux
    port map (
            O => \N__66178\,
            I => \N__66126\
        );

    \I__15896\ : InMux
    port map (
            O => \N__66177\,
            I => \N__66126\
        );

    \I__15895\ : Span4Mux_v
    port map (
            O => \N__66172\,
            I => \N__66122\
        );

    \I__15894\ : LocalMux
    port map (
            O => \N__66169\,
            I => \N__66117\
        );

    \I__15893\ : LocalMux
    port map (
            O => \N__66166\,
            I => \N__66114\
        );

    \I__15892\ : LocalMux
    port map (
            O => \N__66163\,
            I => \N__66111\
        );

    \I__15891\ : InMux
    port map (
            O => \N__66162\,
            I => \N__66102\
        );

    \I__15890\ : InMux
    port map (
            O => \N__66159\,
            I => \N__66102\
        );

    \I__15889\ : InMux
    port map (
            O => \N__66158\,
            I => \N__66102\
        );

    \I__15888\ : InMux
    port map (
            O => \N__66157\,
            I => \N__66102\
        );

    \I__15887\ : InMux
    port map (
            O => \N__66156\,
            I => \N__66099\
        );

    \I__15886\ : InMux
    port map (
            O => \N__66155\,
            I => \N__66096\
        );

    \I__15885\ : InMux
    port map (
            O => \N__66154\,
            I => \N__66093\
        );

    \I__15884\ : InMux
    port map (
            O => \N__66153\,
            I => \N__66084\
        );

    \I__15883\ : InMux
    port map (
            O => \N__66150\,
            I => \N__66084\
        );

    \I__15882\ : InMux
    port map (
            O => \N__66147\,
            I => \N__66084\
        );

    \I__15881\ : InMux
    port map (
            O => \N__66146\,
            I => \N__66084\
        );

    \I__15880\ : InMux
    port map (
            O => \N__66145\,
            I => \N__66081\
        );

    \I__15879\ : InMux
    port map (
            O => \N__66144\,
            I => \N__66078\
        );

    \I__15878\ : InMux
    port map (
            O => \N__66141\,
            I => \N__66071\
        );

    \I__15877\ : InMux
    port map (
            O => \N__66140\,
            I => \N__66071\
        );

    \I__15876\ : InMux
    port map (
            O => \N__66139\,
            I => \N__66071\
        );

    \I__15875\ : LocalMux
    port map (
            O => \N__66136\,
            I => \N__66068\
        );

    \I__15874\ : LocalMux
    port map (
            O => \N__66133\,
            I => \N__66061\
        );

    \I__15873\ : LocalMux
    port map (
            O => \N__66126\,
            I => \N__66061\
        );

    \I__15872\ : InMux
    port map (
            O => \N__66125\,
            I => \N__66057\
        );

    \I__15871\ : Span4Mux_h
    port map (
            O => \N__66122\,
            I => \N__66054\
        );

    \I__15870\ : InMux
    port map (
            O => \N__66121\,
            I => \N__66051\
        );

    \I__15869\ : CascadeMux
    port map (
            O => \N__66120\,
            I => \N__66047\
        );

    \I__15868\ : Span4Mux_h
    port map (
            O => \N__66117\,
            I => \N__66040\
        );

    \I__15867\ : Span4Mux_h
    port map (
            O => \N__66114\,
            I => \N__66040\
        );

    \I__15866\ : Span4Mux_v
    port map (
            O => \N__66111\,
            I => \N__66033\
        );

    \I__15865\ : LocalMux
    port map (
            O => \N__66102\,
            I => \N__66033\
        );

    \I__15864\ : LocalMux
    port map (
            O => \N__66099\,
            I => \N__66026\
        );

    \I__15863\ : LocalMux
    port map (
            O => \N__66096\,
            I => \N__66026\
        );

    \I__15862\ : LocalMux
    port map (
            O => \N__66093\,
            I => \N__66026\
        );

    \I__15861\ : LocalMux
    port map (
            O => \N__66084\,
            I => \N__66023\
        );

    \I__15860\ : LocalMux
    port map (
            O => \N__66081\,
            I => \N__66020\
        );

    \I__15859\ : LocalMux
    port map (
            O => \N__66078\,
            I => \N__66013\
        );

    \I__15858\ : LocalMux
    port map (
            O => \N__66071\,
            I => \N__66013\
        );

    \I__15857\ : Span4Mux_v
    port map (
            O => \N__66068\,
            I => \N__66013\
        );

    \I__15856\ : InMux
    port map (
            O => \N__66067\,
            I => \N__66008\
        );

    \I__15855\ : CascadeMux
    port map (
            O => \N__66066\,
            I => \N__66004\
        );

    \I__15854\ : Span4Mux_v
    port map (
            O => \N__66061\,
            I => \N__66001\
        );

    \I__15853\ : InMux
    port map (
            O => \N__66060\,
            I => \N__65998\
        );

    \I__15852\ : LocalMux
    port map (
            O => \N__66057\,
            I => \N__65995\
        );

    \I__15851\ : Span4Mux_v
    port map (
            O => \N__66054\,
            I => \N__65992\
        );

    \I__15850\ : LocalMux
    port map (
            O => \N__66051\,
            I => \N__65989\
        );

    \I__15849\ : InMux
    port map (
            O => \N__66050\,
            I => \N__65986\
        );

    \I__15848\ : InMux
    port map (
            O => \N__66047\,
            I => \N__65979\
        );

    \I__15847\ : InMux
    port map (
            O => \N__66046\,
            I => \N__65979\
        );

    \I__15846\ : InMux
    port map (
            O => \N__66045\,
            I => \N__65979\
        );

    \I__15845\ : Span4Mux_h
    port map (
            O => \N__66040\,
            I => \N__65976\
        );

    \I__15844\ : InMux
    port map (
            O => \N__66039\,
            I => \N__65971\
        );

    \I__15843\ : InMux
    port map (
            O => \N__66038\,
            I => \N__65971\
        );

    \I__15842\ : Span4Mux_v
    port map (
            O => \N__66033\,
            I => \N__65968\
        );

    \I__15841\ : Span4Mux_v
    port map (
            O => \N__66026\,
            I => \N__65965\
        );

    \I__15840\ : Span4Mux_v
    port map (
            O => \N__66023\,
            I => \N__65958\
        );

    \I__15839\ : Span4Mux_h
    port map (
            O => \N__66020\,
            I => \N__65958\
        );

    \I__15838\ : Span4Mux_v
    port map (
            O => \N__66013\,
            I => \N__65958\
        );

    \I__15837\ : InMux
    port map (
            O => \N__66012\,
            I => \N__65955\
        );

    \I__15836\ : InMux
    port map (
            O => \N__66011\,
            I => \N__65952\
        );

    \I__15835\ : LocalMux
    port map (
            O => \N__66008\,
            I => \N__65949\
        );

    \I__15834\ : InMux
    port map (
            O => \N__66007\,
            I => \N__65944\
        );

    \I__15833\ : InMux
    port map (
            O => \N__66004\,
            I => \N__65944\
        );

    \I__15832\ : Span4Mux_v
    port map (
            O => \N__66001\,
            I => \N__65941\
        );

    \I__15831\ : LocalMux
    port map (
            O => \N__65998\,
            I => \N__65936\
        );

    \I__15830\ : Span4Mux_h
    port map (
            O => \N__65995\,
            I => \N__65936\
        );

    \I__15829\ : Sp12to4
    port map (
            O => \N__65992\,
            I => \N__65933\
        );

    \I__15828\ : Span4Mux_h
    port map (
            O => \N__65989\,
            I => \N__65930\
        );

    \I__15827\ : LocalMux
    port map (
            O => \N__65986\,
            I => \N__65921\
        );

    \I__15826\ : LocalMux
    port map (
            O => \N__65979\,
            I => \N__65921\
        );

    \I__15825\ : Span4Mux_h
    port map (
            O => \N__65976\,
            I => \N__65921\
        );

    \I__15824\ : LocalMux
    port map (
            O => \N__65971\,
            I => \N__65921\
        );

    \I__15823\ : Span4Mux_h
    port map (
            O => \N__65968\,
            I => \N__65918\
        );

    \I__15822\ : Span4Mux_v
    port map (
            O => \N__65965\,
            I => \N__65913\
        );

    \I__15821\ : Span4Mux_v
    port map (
            O => \N__65958\,
            I => \N__65913\
        );

    \I__15820\ : LocalMux
    port map (
            O => \N__65955\,
            I => \N__65904\
        );

    \I__15819\ : LocalMux
    port map (
            O => \N__65952\,
            I => \N__65904\
        );

    \I__15818\ : Sp12to4
    port map (
            O => \N__65949\,
            I => \N__65904\
        );

    \I__15817\ : LocalMux
    port map (
            O => \N__65944\,
            I => \N__65904\
        );

    \I__15816\ : Span4Mux_h
    port map (
            O => \N__65941\,
            I => \N__65901\
        );

    \I__15815\ : Sp12to4
    port map (
            O => \N__65936\,
            I => \N__65894\
        );

    \I__15814\ : Span12Mux_h
    port map (
            O => \N__65933\,
            I => \N__65894\
        );

    \I__15813\ : Sp12to4
    port map (
            O => \N__65930\,
            I => \N__65894\
        );

    \I__15812\ : Span4Mux_v
    port map (
            O => \N__65921\,
            I => \N__65891\
        );

    \I__15811\ : Span4Mux_v
    port map (
            O => \N__65918\,
            I => \N__65888\
        );

    \I__15810\ : Span4Mux_h
    port map (
            O => \N__65913\,
            I => \N__65885\
        );

    \I__15809\ : Span12Mux_h
    port map (
            O => \N__65904\,
            I => \N__65878\
        );

    \I__15808\ : Sp12to4
    port map (
            O => \N__65901\,
            I => \N__65878\
        );

    \I__15807\ : Span12Mux_v
    port map (
            O => \N__65894\,
            I => \N__65878\
        );

    \I__15806\ : Odrv4
    port map (
            O => \N__65891\,
            I => \c0.n12_adj_3265\
        );

    \I__15805\ : Odrv4
    port map (
            O => \N__65888\,
            I => \c0.n12_adj_3265\
        );

    \I__15804\ : Odrv4
    port map (
            O => \N__65885\,
            I => \c0.n12_adj_3265\
        );

    \I__15803\ : Odrv12
    port map (
            O => \N__65878\,
            I => \c0.n12_adj_3265\
        );

    \I__15802\ : CascadeMux
    port map (
            O => \N__65869\,
            I => \N__65865\
        );

    \I__15801\ : InMux
    port map (
            O => \N__65868\,
            I => \N__65860\
        );

    \I__15800\ : InMux
    port map (
            O => \N__65865\,
            I => \N__65857\
        );

    \I__15799\ : InMux
    port map (
            O => \N__65864\,
            I => \N__65854\
        );

    \I__15798\ : CascadeMux
    port map (
            O => \N__65863\,
            I => \N__65850\
        );

    \I__15797\ : LocalMux
    port map (
            O => \N__65860\,
            I => \N__65846\
        );

    \I__15796\ : LocalMux
    port map (
            O => \N__65857\,
            I => \N__65843\
        );

    \I__15795\ : LocalMux
    port map (
            O => \N__65854\,
            I => \N__65840\
        );

    \I__15794\ : InMux
    port map (
            O => \N__65853\,
            I => \N__65837\
        );

    \I__15793\ : InMux
    port map (
            O => \N__65850\,
            I => \N__65834\
        );

    \I__15792\ : InMux
    port map (
            O => \N__65849\,
            I => \N__65831\
        );

    \I__15791\ : Span4Mux_v
    port map (
            O => \N__65846\,
            I => \N__65828\
        );

    \I__15790\ : Span4Mux_v
    port map (
            O => \N__65843\,
            I => \N__65823\
        );

    \I__15789\ : Span4Mux_v
    port map (
            O => \N__65840\,
            I => \N__65823\
        );

    \I__15788\ : LocalMux
    port map (
            O => \N__65837\,
            I => \N__65818\
        );

    \I__15787\ : LocalMux
    port map (
            O => \N__65834\,
            I => \N__65818\
        );

    \I__15786\ : LocalMux
    port map (
            O => \N__65831\,
            I => \N__65815\
        );

    \I__15785\ : Span4Mux_h
    port map (
            O => \N__65828\,
            I => \N__65812\
        );

    \I__15784\ : Span4Mux_h
    port map (
            O => \N__65823\,
            I => \N__65809\
        );

    \I__15783\ : Span4Mux_v
    port map (
            O => \N__65818\,
            I => \N__65806\
        );

    \I__15782\ : Odrv12
    port map (
            O => \N__65815\,
            I => \c0.data_in_frame_12_3\
        );

    \I__15781\ : Odrv4
    port map (
            O => \N__65812\,
            I => \c0.data_in_frame_12_3\
        );

    \I__15780\ : Odrv4
    port map (
            O => \N__65809\,
            I => \c0.data_in_frame_12_3\
        );

    \I__15779\ : Odrv4
    port map (
            O => \N__65806\,
            I => \c0.data_in_frame_12_3\
        );

    \I__15778\ : InMux
    port map (
            O => \N__65797\,
            I => \N__65792\
        );

    \I__15777\ : InMux
    port map (
            O => \N__65796\,
            I => \N__65789\
        );

    \I__15776\ : InMux
    port map (
            O => \N__65795\,
            I => \N__65786\
        );

    \I__15775\ : LocalMux
    port map (
            O => \N__65792\,
            I => \N__65783\
        );

    \I__15774\ : LocalMux
    port map (
            O => \N__65789\,
            I => \N__65775\
        );

    \I__15773\ : LocalMux
    port map (
            O => \N__65786\,
            I => \N__65775\
        );

    \I__15772\ : Span4Mux_v
    port map (
            O => \N__65783\,
            I => \N__65772\
        );

    \I__15771\ : InMux
    port map (
            O => \N__65782\,
            I => \N__65769\
        );

    \I__15770\ : InMux
    port map (
            O => \N__65781\,
            I => \N__65766\
        );

    \I__15769\ : InMux
    port map (
            O => \N__65780\,
            I => \N__65763\
        );

    \I__15768\ : Span4Mux_v
    port map (
            O => \N__65775\,
            I => \N__65759\
        );

    \I__15767\ : Sp12to4
    port map (
            O => \N__65772\,
            I => \N__65752\
        );

    \I__15766\ : LocalMux
    port map (
            O => \N__65769\,
            I => \N__65752\
        );

    \I__15765\ : LocalMux
    port map (
            O => \N__65766\,
            I => \N__65752\
        );

    \I__15764\ : LocalMux
    port map (
            O => \N__65763\,
            I => \N__65749\
        );

    \I__15763\ : CascadeMux
    port map (
            O => \N__65762\,
            I => \N__65746\
        );

    \I__15762\ : Span4Mux_h
    port map (
            O => \N__65759\,
            I => \N__65743\
        );

    \I__15761\ : Span12Mux_h
    port map (
            O => \N__65752\,
            I => \N__65738\
        );

    \I__15760\ : Sp12to4
    port map (
            O => \N__65749\,
            I => \N__65738\
        );

    \I__15759\ : InMux
    port map (
            O => \N__65746\,
            I => \N__65735\
        );

    \I__15758\ : Span4Mux_v
    port map (
            O => \N__65743\,
            I => \N__65732\
        );

    \I__15757\ : Span12Mux_v
    port map (
            O => \N__65738\,
            I => \N__65729\
        );

    \I__15756\ : LocalMux
    port map (
            O => \N__65735\,
            I => data_in_frame_19_2
        );

    \I__15755\ : Odrv4
    port map (
            O => \N__65732\,
            I => data_in_frame_19_2
        );

    \I__15754\ : Odrv12
    port map (
            O => \N__65729\,
            I => data_in_frame_19_2
        );

    \I__15753\ : InMux
    port map (
            O => \N__65722\,
            I => \N__65719\
        );

    \I__15752\ : LocalMux
    port map (
            O => \N__65719\,
            I => \N__65716\
        );

    \I__15751\ : Span4Mux_h
    port map (
            O => \N__65716\,
            I => \N__65712\
        );

    \I__15750\ : InMux
    port map (
            O => \N__65715\,
            I => \N__65708\
        );

    \I__15749\ : Span4Mux_h
    port map (
            O => \N__65712\,
            I => \N__65705\
        );

    \I__15748\ : InMux
    port map (
            O => \N__65711\,
            I => \N__65702\
        );

    \I__15747\ : LocalMux
    port map (
            O => \N__65708\,
            I => data_in_frame_19_5
        );

    \I__15746\ : Odrv4
    port map (
            O => \N__65705\,
            I => data_in_frame_19_5
        );

    \I__15745\ : LocalMux
    port map (
            O => \N__65702\,
            I => data_in_frame_19_5
        );

    \I__15744\ : InMux
    port map (
            O => \N__65695\,
            I => \N__65690\
        );

    \I__15743\ : InMux
    port map (
            O => \N__65694\,
            I => \N__65687\
        );

    \I__15742\ : InMux
    port map (
            O => \N__65693\,
            I => \N__65684\
        );

    \I__15741\ : LocalMux
    port map (
            O => \N__65690\,
            I => \N__65681\
        );

    \I__15740\ : LocalMux
    port map (
            O => \N__65687\,
            I => \N__65675\
        );

    \I__15739\ : LocalMux
    port map (
            O => \N__65684\,
            I => \N__65675\
        );

    \I__15738\ : Span4Mux_h
    port map (
            O => \N__65681\,
            I => \N__65671\
        );

    \I__15737\ : InMux
    port map (
            O => \N__65680\,
            I => \N__65668\
        );

    \I__15736\ : Span4Mux_h
    port map (
            O => \N__65675\,
            I => \N__65665\
        );

    \I__15735\ : CascadeMux
    port map (
            O => \N__65674\,
            I => \N__65662\
        );

    \I__15734\ : Span4Mux_v
    port map (
            O => \N__65671\,
            I => \N__65658\
        );

    \I__15733\ : LocalMux
    port map (
            O => \N__65668\,
            I => \N__65655\
        );

    \I__15732\ : Span4Mux_h
    port map (
            O => \N__65665\,
            I => \N__65652\
        );

    \I__15731\ : InMux
    port map (
            O => \N__65662\,
            I => \N__65649\
        );

    \I__15730\ : InMux
    port map (
            O => \N__65661\,
            I => \N__65646\
        );

    \I__15729\ : Span4Mux_v
    port map (
            O => \N__65658\,
            I => \N__65643\
        );

    \I__15728\ : Span4Mux_h
    port map (
            O => \N__65655\,
            I => \N__65638\
        );

    \I__15727\ : Span4Mux_v
    port map (
            O => \N__65652\,
            I => \N__65638\
        );

    \I__15726\ : LocalMux
    port map (
            O => \N__65649\,
            I => \N__65635\
        );

    \I__15725\ : LocalMux
    port map (
            O => \N__65646\,
            I => data_in_frame_19_1
        );

    \I__15724\ : Odrv4
    port map (
            O => \N__65643\,
            I => data_in_frame_19_1
        );

    \I__15723\ : Odrv4
    port map (
            O => \N__65638\,
            I => data_in_frame_19_1
        );

    \I__15722\ : Odrv12
    port map (
            O => \N__65635\,
            I => data_in_frame_19_1
        );

    \I__15721\ : InMux
    port map (
            O => \N__65626\,
            I => \N__65623\
        );

    \I__15720\ : LocalMux
    port map (
            O => \N__65623\,
            I => \N__65620\
        );

    \I__15719\ : Span4Mux_h
    port map (
            O => \N__65620\,
            I => \N__65615\
        );

    \I__15718\ : InMux
    port map (
            O => \N__65619\,
            I => \N__65610\
        );

    \I__15717\ : InMux
    port map (
            O => \N__65618\,
            I => \N__65610\
        );

    \I__15716\ : Odrv4
    port map (
            O => \N__65615\,
            I => \c0.n6166\
        );

    \I__15715\ : LocalMux
    port map (
            O => \N__65610\,
            I => \c0.n6166\
        );

    \I__15714\ : InMux
    port map (
            O => \N__65605\,
            I => \N__65602\
        );

    \I__15713\ : LocalMux
    port map (
            O => \N__65602\,
            I => \N__65599\
        );

    \I__15712\ : Span4Mux_h
    port map (
            O => \N__65599\,
            I => \N__65591\
        );

    \I__15711\ : InMux
    port map (
            O => \N__65598\,
            I => \N__65587\
        );

    \I__15710\ : InMux
    port map (
            O => \N__65597\,
            I => \N__65584\
        );

    \I__15709\ : InMux
    port map (
            O => \N__65596\,
            I => \N__65581\
        );

    \I__15708\ : InMux
    port map (
            O => \N__65595\,
            I => \N__65575\
        );

    \I__15707\ : InMux
    port map (
            O => \N__65594\,
            I => \N__65575\
        );

    \I__15706\ : Span4Mux_h
    port map (
            O => \N__65591\,
            I => \N__65572\
        );

    \I__15705\ : InMux
    port map (
            O => \N__65590\,
            I => \N__65569\
        );

    \I__15704\ : LocalMux
    port map (
            O => \N__65587\,
            I => \N__65566\
        );

    \I__15703\ : LocalMux
    port map (
            O => \N__65584\,
            I => \N__65563\
        );

    \I__15702\ : LocalMux
    port map (
            O => \N__65581\,
            I => \N__65560\
        );

    \I__15701\ : InMux
    port map (
            O => \N__65580\,
            I => \N__65557\
        );

    \I__15700\ : LocalMux
    port map (
            O => \N__65575\,
            I => \N__65554\
        );

    \I__15699\ : Sp12to4
    port map (
            O => \N__65572\,
            I => \N__65551\
        );

    \I__15698\ : LocalMux
    port map (
            O => \N__65569\,
            I => \N__65544\
        );

    \I__15697\ : Sp12to4
    port map (
            O => \N__65566\,
            I => \N__65544\
        );

    \I__15696\ : Sp12to4
    port map (
            O => \N__65563\,
            I => \N__65544\
        );

    \I__15695\ : Sp12to4
    port map (
            O => \N__65560\,
            I => \N__65541\
        );

    \I__15694\ : LocalMux
    port map (
            O => \N__65557\,
            I => \N__65532\
        );

    \I__15693\ : Span12Mux_v
    port map (
            O => \N__65554\,
            I => \N__65532\
        );

    \I__15692\ : Span12Mux_v
    port map (
            O => \N__65551\,
            I => \N__65532\
        );

    \I__15691\ : Span12Mux_v
    port map (
            O => \N__65544\,
            I => \N__65532\
        );

    \I__15690\ : Odrv12
    port map (
            O => \N__65541\,
            I => n19130
        );

    \I__15689\ : Odrv12
    port map (
            O => \N__65532\,
            I => n19130
        );

    \I__15688\ : InMux
    port map (
            O => \N__65527\,
            I => \N__65522\
        );

    \I__15687\ : CascadeMux
    port map (
            O => \N__65526\,
            I => \N__65516\
        );

    \I__15686\ : InMux
    port map (
            O => \N__65525\,
            I => \N__65512\
        );

    \I__15685\ : LocalMux
    port map (
            O => \N__65522\,
            I => \N__65509\
        );

    \I__15684\ : InMux
    port map (
            O => \N__65521\,
            I => \N__65504\
        );

    \I__15683\ : InMux
    port map (
            O => \N__65520\,
            I => \N__65504\
        );

    \I__15682\ : InMux
    port map (
            O => \N__65519\,
            I => \N__65499\
        );

    \I__15681\ : InMux
    port map (
            O => \N__65516\,
            I => \N__65499\
        );

    \I__15680\ : InMux
    port map (
            O => \N__65515\,
            I => \N__65496\
        );

    \I__15679\ : LocalMux
    port map (
            O => \N__65512\,
            I => \N__65490\
        );

    \I__15678\ : Span4Mux_h
    port map (
            O => \N__65509\,
            I => \N__65485\
        );

    \I__15677\ : LocalMux
    port map (
            O => \N__65504\,
            I => \N__65485\
        );

    \I__15676\ : LocalMux
    port map (
            O => \N__65499\,
            I => \N__65482\
        );

    \I__15675\ : LocalMux
    port map (
            O => \N__65496\,
            I => \N__65479\
        );

    \I__15674\ : InMux
    port map (
            O => \N__65495\,
            I => \N__65474\
        );

    \I__15673\ : InMux
    port map (
            O => \N__65494\,
            I => \N__65474\
        );

    \I__15672\ : InMux
    port map (
            O => \N__65493\,
            I => \N__65471\
        );

    \I__15671\ : Span4Mux_h
    port map (
            O => \N__65490\,
            I => \N__65466\
        );

    \I__15670\ : Span4Mux_v
    port map (
            O => \N__65485\,
            I => \N__65466\
        );

    \I__15669\ : Span4Mux_h
    port map (
            O => \N__65482\,
            I => \N__65459\
        );

    \I__15668\ : Span4Mux_h
    port map (
            O => \N__65479\,
            I => \N__65459\
        );

    \I__15667\ : LocalMux
    port map (
            O => \N__65474\,
            I => \N__65459\
        );

    \I__15666\ : LocalMux
    port map (
            O => \N__65471\,
            I => data_in_frame_16_2
        );

    \I__15665\ : Odrv4
    port map (
            O => \N__65466\,
            I => data_in_frame_16_2
        );

    \I__15664\ : Odrv4
    port map (
            O => \N__65459\,
            I => data_in_frame_16_2
        );

    \I__15663\ : InMux
    port map (
            O => \N__65452\,
            I => \N__65449\
        );

    \I__15662\ : LocalMux
    port map (
            O => \N__65449\,
            I => \N__65445\
        );

    \I__15661\ : InMux
    port map (
            O => \N__65448\,
            I => \N__65442\
        );

    \I__15660\ : Span4Mux_v
    port map (
            O => \N__65445\,
            I => \N__65439\
        );

    \I__15659\ : LocalMux
    port map (
            O => \N__65442\,
            I => \c0.data_in_frame_28_5\
        );

    \I__15658\ : Odrv4
    port map (
            O => \N__65439\,
            I => \c0.data_in_frame_28_5\
        );

    \I__15657\ : InMux
    port map (
            O => \N__65434\,
            I => \N__65430\
        );

    \I__15656\ : CascadeMux
    port map (
            O => \N__65433\,
            I => \N__65426\
        );

    \I__15655\ : LocalMux
    port map (
            O => \N__65430\,
            I => \N__65423\
        );

    \I__15654\ : InMux
    port map (
            O => \N__65429\,
            I => \N__65420\
        );

    \I__15653\ : InMux
    port map (
            O => \N__65426\,
            I => \N__65417\
        );

    \I__15652\ : Span4Mux_h
    port map (
            O => \N__65423\,
            I => \N__65412\
        );

    \I__15651\ : LocalMux
    port map (
            O => \N__65420\,
            I => \N__65412\
        );

    \I__15650\ : LocalMux
    port map (
            O => \N__65417\,
            I => \c0.n19381\
        );

    \I__15649\ : Odrv4
    port map (
            O => \N__65412\,
            I => \c0.n19381\
        );

    \I__15648\ : InMux
    port map (
            O => \N__65407\,
            I => \N__65403\
        );

    \I__15647\ : InMux
    port map (
            O => \N__65406\,
            I => \N__65400\
        );

    \I__15646\ : LocalMux
    port map (
            O => \N__65403\,
            I => \N__65394\
        );

    \I__15645\ : LocalMux
    port map (
            O => \N__65400\,
            I => \N__65391\
        );

    \I__15644\ : InMux
    port map (
            O => \N__65399\,
            I => \N__65388\
        );

    \I__15643\ : InMux
    port map (
            O => \N__65398\,
            I => \N__65385\
        );

    \I__15642\ : CascadeMux
    port map (
            O => \N__65397\,
            I => \N__65382\
        );

    \I__15641\ : Span4Mux_h
    port map (
            O => \N__65394\,
            I => \N__65379\
        );

    \I__15640\ : Span4Mux_h
    port map (
            O => \N__65391\,
            I => \N__65374\
        );

    \I__15639\ : LocalMux
    port map (
            O => \N__65388\,
            I => \N__65374\
        );

    \I__15638\ : LocalMux
    port map (
            O => \N__65385\,
            I => \N__65371\
        );

    \I__15637\ : InMux
    port map (
            O => \N__65382\,
            I => \N__65368\
        );

    \I__15636\ : Span4Mux_v
    port map (
            O => \N__65379\,
            I => \N__65365\
        );

    \I__15635\ : Span4Mux_v
    port map (
            O => \N__65374\,
            I => \N__65362\
        );

    \I__15634\ : Span4Mux_v
    port map (
            O => \N__65371\,
            I => \N__65359\
        );

    \I__15633\ : LocalMux
    port map (
            O => \N__65368\,
            I => \c0.data_in_frame_7_0\
        );

    \I__15632\ : Odrv4
    port map (
            O => \N__65365\,
            I => \c0.data_in_frame_7_0\
        );

    \I__15631\ : Odrv4
    port map (
            O => \N__65362\,
            I => \c0.data_in_frame_7_0\
        );

    \I__15630\ : Odrv4
    port map (
            O => \N__65359\,
            I => \c0.data_in_frame_7_0\
        );

    \I__15629\ : CascadeMux
    port map (
            O => \N__65350\,
            I => \N__65347\
        );

    \I__15628\ : InMux
    port map (
            O => \N__65347\,
            I => \N__65344\
        );

    \I__15627\ : LocalMux
    port map (
            O => \N__65344\,
            I => \N__65340\
        );

    \I__15626\ : InMux
    port map (
            O => \N__65343\,
            I => \N__65337\
        );

    \I__15625\ : Span4Mux_h
    port map (
            O => \N__65340\,
            I => \N__65334\
        );

    \I__15624\ : LocalMux
    port map (
            O => \N__65337\,
            I => \N__65331\
        );

    \I__15623\ : Odrv4
    port map (
            O => \N__65334\,
            I => \c0.n7_adj_3355\
        );

    \I__15622\ : Odrv12
    port map (
            O => \N__65331\,
            I => \c0.n7_adj_3355\
        );

    \I__15621\ : CascadeMux
    port map (
            O => \N__65326\,
            I => \N__65322\
        );

    \I__15620\ : InMux
    port map (
            O => \N__65325\,
            I => \N__65317\
        );

    \I__15619\ : InMux
    port map (
            O => \N__65322\,
            I => \N__65314\
        );

    \I__15618\ : InMux
    port map (
            O => \N__65321\,
            I => \N__65309\
        );

    \I__15617\ : InMux
    port map (
            O => \N__65320\,
            I => \N__65309\
        );

    \I__15616\ : LocalMux
    port map (
            O => \N__65317\,
            I => \N__65306\
        );

    \I__15615\ : LocalMux
    port map (
            O => \N__65314\,
            I => \c0.data_in_frame_17_5\
        );

    \I__15614\ : LocalMux
    port map (
            O => \N__65309\,
            I => \c0.data_in_frame_17_5\
        );

    \I__15613\ : Odrv4
    port map (
            O => \N__65306\,
            I => \c0.data_in_frame_17_5\
        );

    \I__15612\ : InMux
    port map (
            O => \N__65299\,
            I => \N__65293\
        );

    \I__15611\ : InMux
    port map (
            O => \N__65298\,
            I => \N__65293\
        );

    \I__15610\ : LocalMux
    port map (
            O => \N__65293\,
            I => \N__65289\
        );

    \I__15609\ : InMux
    port map (
            O => \N__65292\,
            I => \N__65286\
        );

    \I__15608\ : Odrv4
    port map (
            O => \N__65289\,
            I => \c0.n11590\
        );

    \I__15607\ : LocalMux
    port map (
            O => \N__65286\,
            I => \c0.n11590\
        );

    \I__15606\ : CascadeMux
    port map (
            O => \N__65281\,
            I => \N__65278\
        );

    \I__15605\ : InMux
    port map (
            O => \N__65278\,
            I => \N__65275\
        );

    \I__15604\ : LocalMux
    port map (
            O => \N__65275\,
            I => \N__65272\
        );

    \I__15603\ : Span4Mux_v
    port map (
            O => \N__65272\,
            I => \N__65269\
        );

    \I__15602\ : Span4Mux_h
    port map (
            O => \N__65269\,
            I => \N__65266\
        );

    \I__15601\ : Odrv4
    port map (
            O => \N__65266\,
            I => \c0.n14_adj_3449\
        );

    \I__15600\ : InMux
    port map (
            O => \N__65263\,
            I => \N__65253\
        );

    \I__15599\ : InMux
    port map (
            O => \N__65262\,
            I => \N__65253\
        );

    \I__15598\ : InMux
    port map (
            O => \N__65261\,
            I => \N__65250\
        );

    \I__15597\ : InMux
    port map (
            O => \N__65260\,
            I => \N__65243\
        );

    \I__15596\ : InMux
    port map (
            O => \N__65259\,
            I => \N__65235\
        );

    \I__15595\ : CascadeMux
    port map (
            O => \N__65258\,
            I => \N__65231\
        );

    \I__15594\ : LocalMux
    port map (
            O => \N__65253\,
            I => \N__65227\
        );

    \I__15593\ : LocalMux
    port map (
            O => \N__65250\,
            I => \N__65223\
        );

    \I__15592\ : InMux
    port map (
            O => \N__65249\,
            I => \N__65218\
        );

    \I__15591\ : InMux
    port map (
            O => \N__65248\,
            I => \N__65218\
        );

    \I__15590\ : InMux
    port map (
            O => \N__65247\,
            I => \N__65212\
        );

    \I__15589\ : InMux
    port map (
            O => \N__65246\,
            I => \N__65212\
        );

    \I__15588\ : LocalMux
    port map (
            O => \N__65243\,
            I => \N__65209\
        );

    \I__15587\ : InMux
    port map (
            O => \N__65242\,
            I => \N__65206\
        );

    \I__15586\ : InMux
    port map (
            O => \N__65241\,
            I => \N__65203\
        );

    \I__15585\ : InMux
    port map (
            O => \N__65240\,
            I => \N__65199\
        );

    \I__15584\ : InMux
    port map (
            O => \N__65239\,
            I => \N__65195\
        );

    \I__15583\ : InMux
    port map (
            O => \N__65238\,
            I => \N__65192\
        );

    \I__15582\ : LocalMux
    port map (
            O => \N__65235\,
            I => \N__65186\
        );

    \I__15581\ : InMux
    port map (
            O => \N__65234\,
            I => \N__65179\
        );

    \I__15580\ : InMux
    port map (
            O => \N__65231\,
            I => \N__65179\
        );

    \I__15579\ : InMux
    port map (
            O => \N__65230\,
            I => \N__65179\
        );

    \I__15578\ : Span4Mux_h
    port map (
            O => \N__65227\,
            I => \N__65176\
        );

    \I__15577\ : InMux
    port map (
            O => \N__65226\,
            I => \N__65173\
        );

    \I__15576\ : Span4Mux_v
    port map (
            O => \N__65223\,
            I => \N__65169\
        );

    \I__15575\ : LocalMux
    port map (
            O => \N__65218\,
            I => \N__65166\
        );

    \I__15574\ : InMux
    port map (
            O => \N__65217\,
            I => \N__65163\
        );

    \I__15573\ : LocalMux
    port map (
            O => \N__65212\,
            I => \N__65160\
        );

    \I__15572\ : Span4Mux_h
    port map (
            O => \N__65209\,
            I => \N__65155\
        );

    \I__15571\ : LocalMux
    port map (
            O => \N__65206\,
            I => \N__65155\
        );

    \I__15570\ : LocalMux
    port map (
            O => \N__65203\,
            I => \N__65152\
        );

    \I__15569\ : InMux
    port map (
            O => \N__65202\,
            I => \N__65149\
        );

    \I__15568\ : LocalMux
    port map (
            O => \N__65199\,
            I => \N__65144\
        );

    \I__15567\ : InMux
    port map (
            O => \N__65198\,
            I => \N__65141\
        );

    \I__15566\ : LocalMux
    port map (
            O => \N__65195\,
            I => \N__65136\
        );

    \I__15565\ : LocalMux
    port map (
            O => \N__65192\,
            I => \N__65136\
        );

    \I__15564\ : InMux
    port map (
            O => \N__65191\,
            I => \N__65129\
        );

    \I__15563\ : InMux
    port map (
            O => \N__65190\,
            I => \N__65129\
        );

    \I__15562\ : InMux
    port map (
            O => \N__65189\,
            I => \N__65129\
        );

    \I__15561\ : Span4Mux_v
    port map (
            O => \N__65186\,
            I => \N__65124\
        );

    \I__15560\ : LocalMux
    port map (
            O => \N__65179\,
            I => \N__65124\
        );

    \I__15559\ : Span4Mux_v
    port map (
            O => \N__65176\,
            I => \N__65119\
        );

    \I__15558\ : LocalMux
    port map (
            O => \N__65173\,
            I => \N__65119\
        );

    \I__15557\ : InMux
    port map (
            O => \N__65172\,
            I => \N__65114\
        );

    \I__15556\ : Span4Mux_h
    port map (
            O => \N__65169\,
            I => \N__65109\
        );

    \I__15555\ : Span4Mux_h
    port map (
            O => \N__65166\,
            I => \N__65109\
        );

    \I__15554\ : LocalMux
    port map (
            O => \N__65163\,
            I => \N__65104\
        );

    \I__15553\ : Span4Mux_h
    port map (
            O => \N__65160\,
            I => \N__65104\
        );

    \I__15552\ : Span4Mux_v
    port map (
            O => \N__65155\,
            I => \N__65101\
        );

    \I__15551\ : Span4Mux_v
    port map (
            O => \N__65152\,
            I => \N__65098\
        );

    \I__15550\ : LocalMux
    port map (
            O => \N__65149\,
            I => \N__65095\
        );

    \I__15549\ : InMux
    port map (
            O => \N__65148\,
            I => \N__65091\
        );

    \I__15548\ : InMux
    port map (
            O => \N__65147\,
            I => \N__65088\
        );

    \I__15547\ : Span4Mux_v
    port map (
            O => \N__65144\,
            I => \N__65085\
        );

    \I__15546\ : LocalMux
    port map (
            O => \N__65141\,
            I => \N__65082\
        );

    \I__15545\ : Span4Mux_v
    port map (
            O => \N__65136\,
            I => \N__65079\
        );

    \I__15544\ : LocalMux
    port map (
            O => \N__65129\,
            I => \N__65074\
        );

    \I__15543\ : Span4Mux_v
    port map (
            O => \N__65124\,
            I => \N__65074\
        );

    \I__15542\ : Span4Mux_h
    port map (
            O => \N__65119\,
            I => \N__65071\
        );

    \I__15541\ : InMux
    port map (
            O => \N__65118\,
            I => \N__65064\
        );

    \I__15540\ : InMux
    port map (
            O => \N__65117\,
            I => \N__65064\
        );

    \I__15539\ : LocalMux
    port map (
            O => \N__65114\,
            I => \N__65057\
        );

    \I__15538\ : Span4Mux_h
    port map (
            O => \N__65109\,
            I => \N__65057\
        );

    \I__15537\ : Span4Mux_h
    port map (
            O => \N__65104\,
            I => \N__65057\
        );

    \I__15536\ : Sp12to4
    port map (
            O => \N__65101\,
            I => \N__65052\
        );

    \I__15535\ : Sp12to4
    port map (
            O => \N__65098\,
            I => \N__65052\
        );

    \I__15534\ : Span4Mux_v
    port map (
            O => \N__65095\,
            I => \N__65049\
        );

    \I__15533\ : InMux
    port map (
            O => \N__65094\,
            I => \N__65046\
        );

    \I__15532\ : LocalMux
    port map (
            O => \N__65091\,
            I => \N__65037\
        );

    \I__15531\ : LocalMux
    port map (
            O => \N__65088\,
            I => \N__65037\
        );

    \I__15530\ : Span4Mux_h
    port map (
            O => \N__65085\,
            I => \N__65037\
        );

    \I__15529\ : Span4Mux_v
    port map (
            O => \N__65082\,
            I => \N__65037\
        );

    \I__15528\ : Span4Mux_v
    port map (
            O => \N__65079\,
            I => \N__65034\
        );

    \I__15527\ : Span4Mux_v
    port map (
            O => \N__65074\,
            I => \N__65031\
        );

    \I__15526\ : Sp12to4
    port map (
            O => \N__65071\,
            I => \N__65028\
        );

    \I__15525\ : InMux
    port map (
            O => \N__65070\,
            I => \N__65025\
        );

    \I__15524\ : InMux
    port map (
            O => \N__65069\,
            I => \N__65022\
        );

    \I__15523\ : LocalMux
    port map (
            O => \N__65064\,
            I => \N__65019\
        );

    \I__15522\ : Sp12to4
    port map (
            O => \N__65057\,
            I => \N__65014\
        );

    \I__15521\ : Span12Mux_h
    port map (
            O => \N__65052\,
            I => \N__65014\
        );

    \I__15520\ : Span4Mux_h
    port map (
            O => \N__65049\,
            I => \N__65011\
        );

    \I__15519\ : LocalMux
    port map (
            O => \N__65046\,
            I => \N__65000\
        );

    \I__15518\ : Sp12to4
    port map (
            O => \N__65037\,
            I => \N__65000\
        );

    \I__15517\ : Sp12to4
    port map (
            O => \N__65034\,
            I => \N__65000\
        );

    \I__15516\ : Sp12to4
    port map (
            O => \N__65031\,
            I => \N__65000\
        );

    \I__15515\ : Span12Mux_v
    port map (
            O => \N__65028\,
            I => \N__65000\
        );

    \I__15514\ : LocalMux
    port map (
            O => \N__65025\,
            I => \N__64991\
        );

    \I__15513\ : LocalMux
    port map (
            O => \N__65022\,
            I => \N__64991\
        );

    \I__15512\ : Span12Mux_h
    port map (
            O => \N__65019\,
            I => \N__64991\
        );

    \I__15511\ : Span12Mux_v
    port map (
            O => \N__65014\,
            I => \N__64991\
        );

    \I__15510\ : Odrv4
    port map (
            O => \N__65011\,
            I => rx_data_0
        );

    \I__15509\ : Odrv12
    port map (
            O => \N__65000\,
            I => rx_data_0
        );

    \I__15508\ : Odrv12
    port map (
            O => \N__64991\,
            I => rx_data_0
        );

    \I__15507\ : InMux
    port map (
            O => \N__64984\,
            I => \N__64980\
        );

    \I__15506\ : InMux
    port map (
            O => \N__64983\,
            I => \N__64976\
        );

    \I__15505\ : LocalMux
    port map (
            O => \N__64980\,
            I => \N__64973\
        );

    \I__15504\ : InMux
    port map (
            O => \N__64979\,
            I => \N__64969\
        );

    \I__15503\ : LocalMux
    port map (
            O => \N__64976\,
            I => \N__64966\
        );

    \I__15502\ : Span4Mux_v
    port map (
            O => \N__64973\,
            I => \N__64963\
        );

    \I__15501\ : InMux
    port map (
            O => \N__64972\,
            I => \N__64960\
        );

    \I__15500\ : LocalMux
    port map (
            O => \N__64969\,
            I => \c0.data_in_frame_15_1\
        );

    \I__15499\ : Odrv12
    port map (
            O => \N__64966\,
            I => \c0.data_in_frame_15_1\
        );

    \I__15498\ : Odrv4
    port map (
            O => \N__64963\,
            I => \c0.data_in_frame_15_1\
        );

    \I__15497\ : LocalMux
    port map (
            O => \N__64960\,
            I => \c0.data_in_frame_15_1\
        );

    \I__15496\ : InMux
    port map (
            O => \N__64951\,
            I => \N__64946\
        );

    \I__15495\ : InMux
    port map (
            O => \N__64950\,
            I => \N__64943\
        );

    \I__15494\ : InMux
    port map (
            O => \N__64949\,
            I => \N__64939\
        );

    \I__15493\ : LocalMux
    port map (
            O => \N__64946\,
            I => \N__64936\
        );

    \I__15492\ : LocalMux
    port map (
            O => \N__64943\,
            I => \N__64933\
        );

    \I__15491\ : CascadeMux
    port map (
            O => \N__64942\,
            I => \N__64930\
        );

    \I__15490\ : LocalMux
    port map (
            O => \N__64939\,
            I => \N__64927\
        );

    \I__15489\ : Span4Mux_h
    port map (
            O => \N__64936\,
            I => \N__64924\
        );

    \I__15488\ : Span4Mux_v
    port map (
            O => \N__64933\,
            I => \N__64921\
        );

    \I__15487\ : InMux
    port map (
            O => \N__64930\,
            I => \N__64917\
        );

    \I__15486\ : Span4Mux_h
    port map (
            O => \N__64927\,
            I => \N__64910\
        );

    \I__15485\ : Span4Mux_v
    port map (
            O => \N__64924\,
            I => \N__64910\
        );

    \I__15484\ : Span4Mux_v
    port map (
            O => \N__64921\,
            I => \N__64910\
        );

    \I__15483\ : InMux
    port map (
            O => \N__64920\,
            I => \N__64907\
        );

    \I__15482\ : LocalMux
    port map (
            O => \N__64917\,
            I => \c0.data_in_frame_14_7\
        );

    \I__15481\ : Odrv4
    port map (
            O => \N__64910\,
            I => \c0.data_in_frame_14_7\
        );

    \I__15480\ : LocalMux
    port map (
            O => \N__64907\,
            I => \c0.data_in_frame_14_7\
        );

    \I__15479\ : InMux
    port map (
            O => \N__64900\,
            I => \N__64896\
        );

    \I__15478\ : InMux
    port map (
            O => \N__64899\,
            I => \N__64893\
        );

    \I__15477\ : LocalMux
    port map (
            O => \N__64896\,
            I => \N__64889\
        );

    \I__15476\ : LocalMux
    port map (
            O => \N__64893\,
            I => \N__64883\
        );

    \I__15475\ : InMux
    port map (
            O => \N__64892\,
            I => \N__64880\
        );

    \I__15474\ : Span4Mux_h
    port map (
            O => \N__64889\,
            I => \N__64877\
        );

    \I__15473\ : InMux
    port map (
            O => \N__64888\,
            I => \N__64874\
        );

    \I__15472\ : CascadeMux
    port map (
            O => \N__64887\,
            I => \N__64871\
        );

    \I__15471\ : InMux
    port map (
            O => \N__64886\,
            I => \N__64868\
        );

    \I__15470\ : Span4Mux_v
    port map (
            O => \N__64883\,
            I => \N__64865\
        );

    \I__15469\ : LocalMux
    port map (
            O => \N__64880\,
            I => \N__64860\
        );

    \I__15468\ : Span4Mux_v
    port map (
            O => \N__64877\,
            I => \N__64860\
        );

    \I__15467\ : LocalMux
    port map (
            O => \N__64874\,
            I => \N__64857\
        );

    \I__15466\ : InMux
    port map (
            O => \N__64871\,
            I => \N__64854\
        );

    \I__15465\ : LocalMux
    port map (
            O => \N__64868\,
            I => \N__64849\
        );

    \I__15464\ : Span4Mux_h
    port map (
            O => \N__64865\,
            I => \N__64849\
        );

    \I__15463\ : Span4Mux_h
    port map (
            O => \N__64860\,
            I => \N__64846\
        );

    \I__15462\ : Span12Mux_h
    port map (
            O => \N__64857\,
            I => \N__64843\
        );

    \I__15461\ : LocalMux
    port map (
            O => \N__64854\,
            I => \c0.data_in_frame_14_6\
        );

    \I__15460\ : Odrv4
    port map (
            O => \N__64849\,
            I => \c0.data_in_frame_14_6\
        );

    \I__15459\ : Odrv4
    port map (
            O => \N__64846\,
            I => \c0.data_in_frame_14_6\
        );

    \I__15458\ : Odrv12
    port map (
            O => \N__64843\,
            I => \c0.data_in_frame_14_6\
        );

    \I__15457\ : InMux
    port map (
            O => \N__64834\,
            I => \N__64827\
        );

    \I__15456\ : InMux
    port map (
            O => \N__64833\,
            I => \N__64822\
        );

    \I__15455\ : InMux
    port map (
            O => \N__64832\,
            I => \N__64822\
        );

    \I__15454\ : CascadeMux
    port map (
            O => \N__64831\,
            I => \N__64818\
        );

    \I__15453\ : InMux
    port map (
            O => \N__64830\,
            I => \N__64815\
        );

    \I__15452\ : LocalMux
    port map (
            O => \N__64827\,
            I => \N__64812\
        );

    \I__15451\ : LocalMux
    port map (
            O => \N__64822\,
            I => \N__64809\
        );

    \I__15450\ : CascadeMux
    port map (
            O => \N__64821\,
            I => \N__64806\
        );

    \I__15449\ : InMux
    port map (
            O => \N__64818\,
            I => \N__64803\
        );

    \I__15448\ : LocalMux
    port map (
            O => \N__64815\,
            I => \N__64800\
        );

    \I__15447\ : Span4Mux_v
    port map (
            O => \N__64812\,
            I => \N__64795\
        );

    \I__15446\ : Span4Mux_v
    port map (
            O => \N__64809\,
            I => \N__64795\
        );

    \I__15445\ : InMux
    port map (
            O => \N__64806\,
            I => \N__64792\
        );

    \I__15444\ : LocalMux
    port map (
            O => \N__64803\,
            I => \N__64789\
        );

    \I__15443\ : Span4Mux_v
    port map (
            O => \N__64800\,
            I => \N__64786\
        );

    \I__15442\ : Sp12to4
    port map (
            O => \N__64795\,
            I => \N__64781\
        );

    \I__15441\ : LocalMux
    port map (
            O => \N__64792\,
            I => \N__64781\
        );

    \I__15440\ : Span4Mux_h
    port map (
            O => \N__64789\,
            I => \N__64776\
        );

    \I__15439\ : Span4Mux_h
    port map (
            O => \N__64786\,
            I => \N__64776\
        );

    \I__15438\ : Odrv12
    port map (
            O => \N__64781\,
            I => \c0.n19554\
        );

    \I__15437\ : Odrv4
    port map (
            O => \N__64776\,
            I => \c0.n19554\
        );

    \I__15436\ : InMux
    port map (
            O => \N__64771\,
            I => \N__64764\
        );

    \I__15435\ : InMux
    port map (
            O => \N__64770\,
            I => \N__64764\
        );

    \I__15434\ : InMux
    port map (
            O => \N__64769\,
            I => \N__64761\
        );

    \I__15433\ : LocalMux
    port map (
            O => \N__64764\,
            I => \N__64757\
        );

    \I__15432\ : LocalMux
    port map (
            O => \N__64761\,
            I => \N__64754\
        );

    \I__15431\ : CascadeMux
    port map (
            O => \N__64760\,
            I => \N__64751\
        );

    \I__15430\ : Span4Mux_v
    port map (
            O => \N__64757\,
            I => \N__64748\
        );

    \I__15429\ : Span4Mux_v
    port map (
            O => \N__64754\,
            I => \N__64745\
        );

    \I__15428\ : InMux
    port map (
            O => \N__64751\,
            I => \N__64742\
        );

    \I__15427\ : Span4Mux_v
    port map (
            O => \N__64748\,
            I => \N__64739\
        );

    \I__15426\ : Span4Mux_v
    port map (
            O => \N__64745\,
            I => \N__64736\
        );

    \I__15425\ : LocalMux
    port map (
            O => \N__64742\,
            I => \N__64731\
        );

    \I__15424\ : Span4Mux_h
    port map (
            O => \N__64739\,
            I => \N__64731\
        );

    \I__15423\ : Span4Mux_v
    port map (
            O => \N__64736\,
            I => \N__64728\
        );

    \I__15422\ : Odrv4
    port map (
            O => \N__64731\,
            I => \c0.data_in_frame_17_4\
        );

    \I__15421\ : Odrv4
    port map (
            O => \N__64728\,
            I => \c0.data_in_frame_17_4\
        );

    \I__15420\ : CascadeMux
    port map (
            O => \N__64723\,
            I => \N__64720\
        );

    \I__15419\ : InMux
    port map (
            O => \N__64720\,
            I => \N__64717\
        );

    \I__15418\ : LocalMux
    port map (
            O => \N__64717\,
            I => \N__64714\
        );

    \I__15417\ : Sp12to4
    port map (
            O => \N__64714\,
            I => \N__64711\
        );

    \I__15416\ : Odrv12
    port map (
            O => \N__64711\,
            I => \c0.n18_adj_3235\
        );

    \I__15415\ : CascadeMux
    port map (
            O => \N__64708\,
            I => \N__64704\
        );

    \I__15414\ : InMux
    port map (
            O => \N__64707\,
            I => \N__64700\
        );

    \I__15413\ : InMux
    port map (
            O => \N__64704\,
            I => \N__64696\
        );

    \I__15412\ : InMux
    port map (
            O => \N__64703\,
            I => \N__64693\
        );

    \I__15411\ : LocalMux
    port map (
            O => \N__64700\,
            I => \N__64690\
        );

    \I__15410\ : InMux
    port map (
            O => \N__64699\,
            I => \N__64687\
        );

    \I__15409\ : LocalMux
    port map (
            O => \N__64696\,
            I => \N__64684\
        );

    \I__15408\ : LocalMux
    port map (
            O => \N__64693\,
            I => \N__64680\
        );

    \I__15407\ : Span4Mux_v
    port map (
            O => \N__64690\,
            I => \N__64675\
        );

    \I__15406\ : LocalMux
    port map (
            O => \N__64687\,
            I => \N__64675\
        );

    \I__15405\ : Span4Mux_h
    port map (
            O => \N__64684\,
            I => \N__64672\
        );

    \I__15404\ : CascadeMux
    port map (
            O => \N__64683\,
            I => \N__64669\
        );

    \I__15403\ : Span4Mux_v
    port map (
            O => \N__64680\,
            I => \N__64666\
        );

    \I__15402\ : Span4Mux_v
    port map (
            O => \N__64675\,
            I => \N__64661\
        );

    \I__15401\ : Span4Mux_v
    port map (
            O => \N__64672\,
            I => \N__64661\
        );

    \I__15400\ : InMux
    port map (
            O => \N__64669\,
            I => \N__64658\
        );

    \I__15399\ : Span4Mux_v
    port map (
            O => \N__64666\,
            I => \N__64655\
        );

    \I__15398\ : Span4Mux_v
    port map (
            O => \N__64661\,
            I => \N__64652\
        );

    \I__15397\ : LocalMux
    port map (
            O => \N__64658\,
            I => \c0.data_in_frame_15_3\
        );

    \I__15396\ : Odrv4
    port map (
            O => \N__64655\,
            I => \c0.data_in_frame_15_3\
        );

    \I__15395\ : Odrv4
    port map (
            O => \N__64652\,
            I => \c0.data_in_frame_15_3\
        );

    \I__15394\ : InMux
    port map (
            O => \N__64645\,
            I => \N__64642\
        );

    \I__15393\ : LocalMux
    port map (
            O => \N__64642\,
            I => \N__64639\
        );

    \I__15392\ : Span4Mux_v
    port map (
            O => \N__64639\,
            I => \N__64636\
        );

    \I__15391\ : Odrv4
    port map (
            O => \N__64636\,
            I => \c0.n10_adj_3483\
        );

    \I__15390\ : InMux
    port map (
            O => \N__64633\,
            I => \N__64629\
        );

    \I__15389\ : InMux
    port map (
            O => \N__64632\,
            I => \N__64625\
        );

    \I__15388\ : LocalMux
    port map (
            O => \N__64629\,
            I => \N__64620\
        );

    \I__15387\ : InMux
    port map (
            O => \N__64628\,
            I => \N__64617\
        );

    \I__15386\ : LocalMux
    port map (
            O => \N__64625\,
            I => \N__64614\
        );

    \I__15385\ : InMux
    port map (
            O => \N__64624\,
            I => \N__64609\
        );

    \I__15384\ : InMux
    port map (
            O => \N__64623\,
            I => \N__64609\
        );

    \I__15383\ : Span4Mux_v
    port map (
            O => \N__64620\,
            I => \N__64603\
        );

    \I__15382\ : LocalMux
    port map (
            O => \N__64617\,
            I => \N__64603\
        );

    \I__15381\ : Span4Mux_v
    port map (
            O => \N__64614\,
            I => \N__64598\
        );

    \I__15380\ : LocalMux
    port map (
            O => \N__64609\,
            I => \N__64598\
        );

    \I__15379\ : InMux
    port map (
            O => \N__64608\,
            I => \N__64595\
        );

    \I__15378\ : Span4Mux_h
    port map (
            O => \N__64603\,
            I => \N__64590\
        );

    \I__15377\ : Span4Mux_v
    port map (
            O => \N__64598\,
            I => \N__64590\
        );

    \I__15376\ : LocalMux
    port map (
            O => \N__64595\,
            I => \c0.n18420\
        );

    \I__15375\ : Odrv4
    port map (
            O => \N__64590\,
            I => \c0.n18420\
        );

    \I__15374\ : InMux
    port map (
            O => \N__64585\,
            I => \N__64579\
        );

    \I__15373\ : InMux
    port map (
            O => \N__64584\,
            I => \N__64574\
        );

    \I__15372\ : InMux
    port map (
            O => \N__64583\,
            I => \N__64569\
        );

    \I__15371\ : InMux
    port map (
            O => \N__64582\,
            I => \N__64569\
        );

    \I__15370\ : LocalMux
    port map (
            O => \N__64579\,
            I => \N__64566\
        );

    \I__15369\ : CascadeMux
    port map (
            O => \N__64578\,
            I => \N__64561\
        );

    \I__15368\ : InMux
    port map (
            O => \N__64577\,
            I => \N__64558\
        );

    \I__15367\ : LocalMux
    port map (
            O => \N__64574\,
            I => \N__64555\
        );

    \I__15366\ : LocalMux
    port map (
            O => \N__64569\,
            I => \N__64552\
        );

    \I__15365\ : Span4Mux_v
    port map (
            O => \N__64566\,
            I => \N__64543\
        );

    \I__15364\ : InMux
    port map (
            O => \N__64565\,
            I => \N__64535\
        );

    \I__15363\ : InMux
    port map (
            O => \N__64564\,
            I => \N__64535\
        );

    \I__15362\ : InMux
    port map (
            O => \N__64561\,
            I => \N__64535\
        );

    \I__15361\ : LocalMux
    port map (
            O => \N__64558\,
            I => \N__64530\
        );

    \I__15360\ : Span4Mux_v
    port map (
            O => \N__64555\,
            I => \N__64530\
        );

    \I__15359\ : Span4Mux_v
    port map (
            O => \N__64552\,
            I => \N__64527\
        );

    \I__15358\ : InMux
    port map (
            O => \N__64551\,
            I => \N__64524\
        );

    \I__15357\ : InMux
    port map (
            O => \N__64550\,
            I => \N__64519\
        );

    \I__15356\ : InMux
    port map (
            O => \N__64549\,
            I => \N__64519\
        );

    \I__15355\ : InMux
    port map (
            O => \N__64548\,
            I => \N__64512\
        );

    \I__15354\ : InMux
    port map (
            O => \N__64547\,
            I => \N__64512\
        );

    \I__15353\ : InMux
    port map (
            O => \N__64546\,
            I => \N__64512\
        );

    \I__15352\ : Span4Mux_h
    port map (
            O => \N__64543\,
            I => \N__64509\
        );

    \I__15351\ : InMux
    port map (
            O => \N__64542\,
            I => \N__64506\
        );

    \I__15350\ : LocalMux
    port map (
            O => \N__64535\,
            I => \N__64503\
        );

    \I__15349\ : Span4Mux_v
    port map (
            O => \N__64530\,
            I => \N__64499\
        );

    \I__15348\ : Span4Mux_v
    port map (
            O => \N__64527\,
            I => \N__64496\
        );

    \I__15347\ : LocalMux
    port map (
            O => \N__64524\,
            I => \N__64493\
        );

    \I__15346\ : LocalMux
    port map (
            O => \N__64519\,
            I => \N__64486\
        );

    \I__15345\ : LocalMux
    port map (
            O => \N__64512\,
            I => \N__64486\
        );

    \I__15344\ : Span4Mux_h
    port map (
            O => \N__64509\,
            I => \N__64486\
        );

    \I__15343\ : LocalMux
    port map (
            O => \N__64506\,
            I => \N__64481\
        );

    \I__15342\ : Span12Mux_h
    port map (
            O => \N__64503\,
            I => \N__64481\
        );

    \I__15341\ : InMux
    port map (
            O => \N__64502\,
            I => \N__64478\
        );

    \I__15340\ : Span4Mux_h
    port map (
            O => \N__64499\,
            I => \N__64475\
        );

    \I__15339\ : Span4Mux_v
    port map (
            O => \N__64496\,
            I => \N__64472\
        );

    \I__15338\ : Span4Mux_h
    port map (
            O => \N__64493\,
            I => \N__64467\
        );

    \I__15337\ : Span4Mux_v
    port map (
            O => \N__64486\,
            I => \N__64467\
        );

    \I__15336\ : Span12Mux_v
    port map (
            O => \N__64481\,
            I => \N__64464\
        );

    \I__15335\ : LocalMux
    port map (
            O => \N__64478\,
            I => \c0.n19131\
        );

    \I__15334\ : Odrv4
    port map (
            O => \N__64475\,
            I => \c0.n19131\
        );

    \I__15333\ : Odrv4
    port map (
            O => \N__64472\,
            I => \c0.n19131\
        );

    \I__15332\ : Odrv4
    port map (
            O => \N__64467\,
            I => \c0.n19131\
        );

    \I__15331\ : Odrv12
    port map (
            O => \N__64464\,
            I => \c0.n19131\
        );

    \I__15330\ : CascadeMux
    port map (
            O => \N__64453\,
            I => \N__64450\
        );

    \I__15329\ : InMux
    port map (
            O => \N__64450\,
            I => \N__64446\
        );

    \I__15328\ : InMux
    port map (
            O => \N__64449\,
            I => \N__64443\
        );

    \I__15327\ : LocalMux
    port map (
            O => \N__64446\,
            I => \N__64439\
        );

    \I__15326\ : LocalMux
    port map (
            O => \N__64443\,
            I => \N__64435\
        );

    \I__15325\ : InMux
    port map (
            O => \N__64442\,
            I => \N__64432\
        );

    \I__15324\ : Span12Mux_h
    port map (
            O => \N__64439\,
            I => \N__64429\
        );

    \I__15323\ : InMux
    port map (
            O => \N__64438\,
            I => \N__64426\
        );

    \I__15322\ : Span4Mux_h
    port map (
            O => \N__64435\,
            I => \N__64423\
        );

    \I__15321\ : LocalMux
    port map (
            O => \N__64432\,
            I => \c0.data_in_frame_11_7\
        );

    \I__15320\ : Odrv12
    port map (
            O => \N__64429\,
            I => \c0.data_in_frame_11_7\
        );

    \I__15319\ : LocalMux
    port map (
            O => \N__64426\,
            I => \c0.data_in_frame_11_7\
        );

    \I__15318\ : Odrv4
    port map (
            O => \N__64423\,
            I => \c0.data_in_frame_11_7\
        );

    \I__15317\ : InMux
    port map (
            O => \N__64414\,
            I => \N__64406\
        );

    \I__15316\ : InMux
    port map (
            O => \N__64413\,
            I => \N__64401\
        );

    \I__15315\ : InMux
    port map (
            O => \N__64412\,
            I => \N__64401\
        );

    \I__15314\ : InMux
    port map (
            O => \N__64411\,
            I => \N__64398\
        );

    \I__15313\ : InMux
    port map (
            O => \N__64410\,
            I => \N__64394\
        );

    \I__15312\ : InMux
    port map (
            O => \N__64409\,
            I => \N__64390\
        );

    \I__15311\ : LocalMux
    port map (
            O => \N__64406\,
            I => \N__64379\
        );

    \I__15310\ : LocalMux
    port map (
            O => \N__64401\,
            I => \N__64379\
        );

    \I__15309\ : LocalMux
    port map (
            O => \N__64398\,
            I => \N__64379\
        );

    \I__15308\ : InMux
    port map (
            O => \N__64397\,
            I => \N__64376\
        );

    \I__15307\ : LocalMux
    port map (
            O => \N__64394\,
            I => \N__64373\
        );

    \I__15306\ : InMux
    port map (
            O => \N__64393\,
            I => \N__64370\
        );

    \I__15305\ : LocalMux
    port map (
            O => \N__64390\,
            I => \N__64367\
        );

    \I__15304\ : CascadeMux
    port map (
            O => \N__64389\,
            I => \N__64363\
        );

    \I__15303\ : InMux
    port map (
            O => \N__64388\,
            I => \N__64355\
        );

    \I__15302\ : InMux
    port map (
            O => \N__64387\,
            I => \N__64355\
        );

    \I__15301\ : InMux
    port map (
            O => \N__64386\,
            I => \N__64355\
        );

    \I__15300\ : Span4Mux_h
    port map (
            O => \N__64379\,
            I => \N__64352\
        );

    \I__15299\ : LocalMux
    port map (
            O => \N__64376\,
            I => \N__64349\
        );

    \I__15298\ : Span4Mux_v
    port map (
            O => \N__64373\,
            I => \N__64346\
        );

    \I__15297\ : LocalMux
    port map (
            O => \N__64370\,
            I => \N__64341\
        );

    \I__15296\ : Span4Mux_v
    port map (
            O => \N__64367\,
            I => \N__64337\
        );

    \I__15295\ : InMux
    port map (
            O => \N__64366\,
            I => \N__64330\
        );

    \I__15294\ : InMux
    port map (
            O => \N__64363\,
            I => \N__64330\
        );

    \I__15293\ : InMux
    port map (
            O => \N__64362\,
            I => \N__64330\
        );

    \I__15292\ : LocalMux
    port map (
            O => \N__64355\,
            I => \N__64327\
        );

    \I__15291\ : Span4Mux_v
    port map (
            O => \N__64352\,
            I => \N__64322\
        );

    \I__15290\ : Span4Mux_v
    port map (
            O => \N__64349\,
            I => \N__64322\
        );

    \I__15289\ : Span4Mux_h
    port map (
            O => \N__64346\,
            I => \N__64319\
        );

    \I__15288\ : InMux
    port map (
            O => \N__64345\,
            I => \N__64314\
        );

    \I__15287\ : InMux
    port map (
            O => \N__64344\,
            I => \N__64314\
        );

    \I__15286\ : Span4Mux_v
    port map (
            O => \N__64341\,
            I => \N__64311\
        );

    \I__15285\ : InMux
    port map (
            O => \N__64340\,
            I => \N__64308\
        );

    \I__15284\ : Span4Mux_h
    port map (
            O => \N__64337\,
            I => \N__64305\
        );

    \I__15283\ : LocalMux
    port map (
            O => \N__64330\,
            I => \N__64302\
        );

    \I__15282\ : Sp12to4
    port map (
            O => \N__64327\,
            I => \N__64299\
        );

    \I__15281\ : Sp12to4
    port map (
            O => \N__64322\,
            I => \N__64296\
        );

    \I__15280\ : Sp12to4
    port map (
            O => \N__64319\,
            I => \N__64293\
        );

    \I__15279\ : LocalMux
    port map (
            O => \N__64314\,
            I => \N__64290\
        );

    \I__15278\ : Sp12to4
    port map (
            O => \N__64311\,
            I => \N__64287\
        );

    \I__15277\ : LocalMux
    port map (
            O => \N__64308\,
            I => \N__64284\
        );

    \I__15276\ : Span4Mux_v
    port map (
            O => \N__64305\,
            I => \N__64279\
        );

    \I__15275\ : Span4Mux_v
    port map (
            O => \N__64302\,
            I => \N__64279\
        );

    \I__15274\ : Span12Mux_v
    port map (
            O => \N__64299\,
            I => \N__64272\
        );

    \I__15273\ : Span12Mux_v
    port map (
            O => \N__64296\,
            I => \N__64272\
        );

    \I__15272\ : Span12Mux_v
    port map (
            O => \N__64293\,
            I => \N__64272\
        );

    \I__15271\ : Span12Mux_s8_v
    port map (
            O => \N__64290\,
            I => \N__64267\
        );

    \I__15270\ : Span12Mux_h
    port map (
            O => \N__64287\,
            I => \N__64267\
        );

    \I__15269\ : Span4Mux_v
    port map (
            O => \N__64284\,
            I => \N__64264\
        );

    \I__15268\ : Odrv4
    port map (
            O => \N__64279\,
            I => \c0.n15489\
        );

    \I__15267\ : Odrv12
    port map (
            O => \N__64272\,
            I => \c0.n15489\
        );

    \I__15266\ : Odrv12
    port map (
            O => \N__64267\,
            I => \c0.n15489\
        );

    \I__15265\ : Odrv4
    port map (
            O => \N__64264\,
            I => \c0.n15489\
        );

    \I__15264\ : InMux
    port map (
            O => \N__64255\,
            I => \N__64239\
        );

    \I__15263\ : InMux
    port map (
            O => \N__64254\,
            I => \N__64228\
        );

    \I__15262\ : InMux
    port map (
            O => \N__64253\,
            I => \N__64228\
        );

    \I__15261\ : InMux
    port map (
            O => \N__64252\,
            I => \N__64228\
        );

    \I__15260\ : InMux
    port map (
            O => \N__64251\,
            I => \N__64228\
        );

    \I__15259\ : InMux
    port map (
            O => \N__64250\,
            I => \N__64225\
        );

    \I__15258\ : CascadeMux
    port map (
            O => \N__64249\,
            I => \N__64222\
        );

    \I__15257\ : InMux
    port map (
            O => \N__64248\,
            I => \N__64217\
        );

    \I__15256\ : InMux
    port map (
            O => \N__64247\,
            I => \N__64210\
        );

    \I__15255\ : InMux
    port map (
            O => \N__64246\,
            I => \N__64210\
        );

    \I__15254\ : InMux
    port map (
            O => \N__64245\,
            I => \N__64210\
        );

    \I__15253\ : InMux
    port map (
            O => \N__64244\,
            I => \N__64203\
        );

    \I__15252\ : InMux
    port map (
            O => \N__64243\,
            I => \N__64203\
        );

    \I__15251\ : InMux
    port map (
            O => \N__64242\,
            I => \N__64203\
        );

    \I__15250\ : LocalMux
    port map (
            O => \N__64239\,
            I => \N__64200\
        );

    \I__15249\ : InMux
    port map (
            O => \N__64238\,
            I => \N__64193\
        );

    \I__15248\ : InMux
    port map (
            O => \N__64237\,
            I => \N__64193\
        );

    \I__15247\ : LocalMux
    port map (
            O => \N__64228\,
            I => \N__64188\
        );

    \I__15246\ : LocalMux
    port map (
            O => \N__64225\,
            I => \N__64188\
        );

    \I__15245\ : InMux
    port map (
            O => \N__64222\,
            I => \N__64185\
        );

    \I__15244\ : InMux
    port map (
            O => \N__64221\,
            I => \N__64180\
        );

    \I__15243\ : InMux
    port map (
            O => \N__64220\,
            I => \N__64177\
        );

    \I__15242\ : LocalMux
    port map (
            O => \N__64217\,
            I => \N__64174\
        );

    \I__15241\ : LocalMux
    port map (
            O => \N__64210\,
            I => \N__64167\
        );

    \I__15240\ : LocalMux
    port map (
            O => \N__64203\,
            I => \N__64167\
        );

    \I__15239\ : Span4Mux_v
    port map (
            O => \N__64200\,
            I => \N__64167\
        );

    \I__15238\ : InMux
    port map (
            O => \N__64199\,
            I => \N__64164\
        );

    \I__15237\ : InMux
    port map (
            O => \N__64198\,
            I => \N__64161\
        );

    \I__15236\ : LocalMux
    port map (
            O => \N__64193\,
            I => \N__64158\
        );

    \I__15235\ : Span4Mux_v
    port map (
            O => \N__64188\,
            I => \N__64153\
        );

    \I__15234\ : LocalMux
    port map (
            O => \N__64185\,
            I => \N__64153\
        );

    \I__15233\ : InMux
    port map (
            O => \N__64184\,
            I => \N__64148\
        );

    \I__15232\ : InMux
    port map (
            O => \N__64183\,
            I => \N__64148\
        );

    \I__15231\ : LocalMux
    port map (
            O => \N__64180\,
            I => \N__64145\
        );

    \I__15230\ : LocalMux
    port map (
            O => \N__64177\,
            I => \N__64140\
        );

    \I__15229\ : Span4Mux_v
    port map (
            O => \N__64174\,
            I => \N__64140\
        );

    \I__15228\ : Span4Mux_v
    port map (
            O => \N__64167\,
            I => \N__64137\
        );

    \I__15227\ : LocalMux
    port map (
            O => \N__64164\,
            I => \N__64133\
        );

    \I__15226\ : LocalMux
    port map (
            O => \N__64161\,
            I => \N__64130\
        );

    \I__15225\ : Span4Mux_v
    port map (
            O => \N__64158\,
            I => \N__64127\
        );

    \I__15224\ : Span4Mux_h
    port map (
            O => \N__64153\,
            I => \N__64124\
        );

    \I__15223\ : LocalMux
    port map (
            O => \N__64148\,
            I => \N__64121\
        );

    \I__15222\ : Span4Mux_h
    port map (
            O => \N__64145\,
            I => \N__64114\
        );

    \I__15221\ : Span4Mux_v
    port map (
            O => \N__64140\,
            I => \N__64114\
        );

    \I__15220\ : Span4Mux_h
    port map (
            O => \N__64137\,
            I => \N__64114\
        );

    \I__15219\ : InMux
    port map (
            O => \N__64136\,
            I => \N__64110\
        );

    \I__15218\ : Span4Mux_v
    port map (
            O => \N__64133\,
            I => \N__64107\
        );

    \I__15217\ : Span4Mux_h
    port map (
            O => \N__64130\,
            I => \N__64104\
        );

    \I__15216\ : Span4Mux_h
    port map (
            O => \N__64127\,
            I => \N__64101\
        );

    \I__15215\ : Sp12to4
    port map (
            O => \N__64124\,
            I => \N__64096\
        );

    \I__15214\ : Span12Mux_s10_v
    port map (
            O => \N__64121\,
            I => \N__64096\
        );

    \I__15213\ : Span4Mux_v
    port map (
            O => \N__64114\,
            I => \N__64093\
        );

    \I__15212\ : InMux
    port map (
            O => \N__64113\,
            I => \N__64090\
        );

    \I__15211\ : LocalMux
    port map (
            O => \N__64110\,
            I => \N__64087\
        );

    \I__15210\ : Span4Mux_h
    port map (
            O => \N__64107\,
            I => \N__64084\
        );

    \I__15209\ : Sp12to4
    port map (
            O => \N__64104\,
            I => \N__64081\
        );

    \I__15208\ : Span4Mux_v
    port map (
            O => \N__64101\,
            I => \N__64078\
        );

    \I__15207\ : Span12Mux_v
    port map (
            O => \N__64096\,
            I => \N__64075\
        );

    \I__15206\ : Span4Mux_v
    port map (
            O => \N__64093\,
            I => \N__64072\
        );

    \I__15205\ : LocalMux
    port map (
            O => \N__64090\,
            I => \c0.n19140\
        );

    \I__15204\ : Odrv12
    port map (
            O => \N__64087\,
            I => \c0.n19140\
        );

    \I__15203\ : Odrv4
    port map (
            O => \N__64084\,
            I => \c0.n19140\
        );

    \I__15202\ : Odrv12
    port map (
            O => \N__64081\,
            I => \c0.n19140\
        );

    \I__15201\ : Odrv4
    port map (
            O => \N__64078\,
            I => \c0.n19140\
        );

    \I__15200\ : Odrv12
    port map (
            O => \N__64075\,
            I => \c0.n19140\
        );

    \I__15199\ : Odrv4
    port map (
            O => \N__64072\,
            I => \c0.n19140\
        );

    \I__15198\ : InMux
    port map (
            O => \N__64057\,
            I => \N__64053\
        );

    \I__15197\ : InMux
    port map (
            O => \N__64056\,
            I => \N__64050\
        );

    \I__15196\ : LocalMux
    port map (
            O => \N__64053\,
            I => \N__64046\
        );

    \I__15195\ : LocalMux
    port map (
            O => \N__64050\,
            I => \N__64043\
        );

    \I__15194\ : CascadeMux
    port map (
            O => \N__64049\,
            I => \N__64040\
        );

    \I__15193\ : Span4Mux_v
    port map (
            O => \N__64046\,
            I => \N__64036\
        );

    \I__15192\ : Span4Mux_h
    port map (
            O => \N__64043\,
            I => \N__64033\
        );

    \I__15191\ : InMux
    port map (
            O => \N__64040\,
            I => \N__64028\
        );

    \I__15190\ : InMux
    port map (
            O => \N__64039\,
            I => \N__64028\
        );

    \I__15189\ : Odrv4
    port map (
            O => \N__64036\,
            I => \c0.data_in_frame_15_5\
        );

    \I__15188\ : Odrv4
    port map (
            O => \N__64033\,
            I => \c0.data_in_frame_15_5\
        );

    \I__15187\ : LocalMux
    port map (
            O => \N__64028\,
            I => \c0.data_in_frame_15_5\
        );

    \I__15186\ : CascadeMux
    port map (
            O => \N__64021\,
            I => \c0.n9_adj_3552_cascade_\
        );

    \I__15185\ : CascadeMux
    port map (
            O => \N__64018\,
            I => \N__64015\
        );

    \I__15184\ : InMux
    port map (
            O => \N__64015\,
            I => \N__64010\
        );

    \I__15183\ : CascadeMux
    port map (
            O => \N__64014\,
            I => \N__64007\
        );

    \I__15182\ : InMux
    port map (
            O => \N__64013\,
            I => \N__64004\
        );

    \I__15181\ : LocalMux
    port map (
            O => \N__64010\,
            I => \N__63999\
        );

    \I__15180\ : InMux
    port map (
            O => \N__64007\,
            I => \N__63996\
        );

    \I__15179\ : LocalMux
    port map (
            O => \N__64004\,
            I => \N__63991\
        );

    \I__15178\ : InMux
    port map (
            O => \N__64003\,
            I => \N__63988\
        );

    \I__15177\ : InMux
    port map (
            O => \N__64002\,
            I => \N__63985\
        );

    \I__15176\ : Span4Mux_v
    port map (
            O => \N__63999\,
            I => \N__63982\
        );

    \I__15175\ : LocalMux
    port map (
            O => \N__63996\,
            I => \N__63979\
        );

    \I__15174\ : InMux
    port map (
            O => \N__63995\,
            I => \N__63974\
        );

    \I__15173\ : InMux
    port map (
            O => \N__63994\,
            I => \N__63974\
        );

    \I__15172\ : Span12Mux_h
    port map (
            O => \N__63991\,
            I => \N__63971\
        );

    \I__15171\ : LocalMux
    port map (
            O => \N__63988\,
            I => \N__63968\
        );

    \I__15170\ : LocalMux
    port map (
            O => \N__63985\,
            I => data_in_frame_18_3
        );

    \I__15169\ : Odrv4
    port map (
            O => \N__63982\,
            I => data_in_frame_18_3
        );

    \I__15168\ : Odrv4
    port map (
            O => \N__63979\,
            I => data_in_frame_18_3
        );

    \I__15167\ : LocalMux
    port map (
            O => \N__63974\,
            I => data_in_frame_18_3
        );

    \I__15166\ : Odrv12
    port map (
            O => \N__63971\,
            I => data_in_frame_18_3
        );

    \I__15165\ : Odrv4
    port map (
            O => \N__63968\,
            I => data_in_frame_18_3
        );

    \I__15164\ : InMux
    port map (
            O => \N__63955\,
            I => \N__63952\
        );

    \I__15163\ : LocalMux
    port map (
            O => \N__63952\,
            I => \N__63949\
        );

    \I__15162\ : Span4Mux_v
    port map (
            O => \N__63949\,
            I => \N__63945\
        );

    \I__15161\ : InMux
    port map (
            O => \N__63948\,
            I => \N__63940\
        );

    \I__15160\ : Span4Mux_h
    port map (
            O => \N__63945\,
            I => \N__63934\
        );

    \I__15159\ : InMux
    port map (
            O => \N__63944\,
            I => \N__63931\
        );

    \I__15158\ : InMux
    port map (
            O => \N__63943\,
            I => \N__63928\
        );

    \I__15157\ : LocalMux
    port map (
            O => \N__63940\,
            I => \N__63925\
        );

    \I__15156\ : InMux
    port map (
            O => \N__63939\,
            I => \N__63922\
        );

    \I__15155\ : InMux
    port map (
            O => \N__63938\,
            I => \N__63919\
        );

    \I__15154\ : InMux
    port map (
            O => \N__63937\,
            I => \N__63916\
        );

    \I__15153\ : Span4Mux_h
    port map (
            O => \N__63934\,
            I => \N__63910\
        );

    \I__15152\ : LocalMux
    port map (
            O => \N__63931\,
            I => \N__63910\
        );

    \I__15151\ : LocalMux
    port map (
            O => \N__63928\,
            I => \N__63907\
        );

    \I__15150\ : Span4Mux_h
    port map (
            O => \N__63925\,
            I => \N__63900\
        );

    \I__15149\ : LocalMux
    port map (
            O => \N__63922\,
            I => \N__63900\
        );

    \I__15148\ : LocalMux
    port map (
            O => \N__63919\,
            I => \N__63900\
        );

    \I__15147\ : LocalMux
    port map (
            O => \N__63916\,
            I => \N__63897\
        );

    \I__15146\ : InMux
    port map (
            O => \N__63915\,
            I => \N__63894\
        );

    \I__15145\ : Span4Mux_v
    port map (
            O => \N__63910\,
            I => \N__63891\
        );

    \I__15144\ : Span4Mux_h
    port map (
            O => \N__63907\,
            I => \N__63888\
        );

    \I__15143\ : Span4Mux_v
    port map (
            O => \N__63900\,
            I => \N__63885\
        );

    \I__15142\ : Span4Mux_v
    port map (
            O => \N__63897\,
            I => \N__63880\
        );

    \I__15141\ : LocalMux
    port map (
            O => \N__63894\,
            I => \N__63880\
        );

    \I__15140\ : Odrv4
    port map (
            O => \N__63891\,
            I => n19129
        );

    \I__15139\ : Odrv4
    port map (
            O => \N__63888\,
            I => n19129
        );

    \I__15138\ : Odrv4
    port map (
            O => \N__63885\,
            I => n19129
        );

    \I__15137\ : Odrv4
    port map (
            O => \N__63880\,
            I => n19129
        );

    \I__15136\ : InMux
    port map (
            O => \N__63871\,
            I => \N__63865\
        );

    \I__15135\ : InMux
    port map (
            O => \N__63870\,
            I => \N__63865\
        );

    \I__15134\ : LocalMux
    port map (
            O => \N__63865\,
            I => data_in_frame_18_4
        );

    \I__15133\ : InMux
    port map (
            O => \N__63862\,
            I => \N__63858\
        );

    \I__15132\ : InMux
    port map (
            O => \N__63861\,
            I => \N__63855\
        );

    \I__15131\ : LocalMux
    port map (
            O => \N__63858\,
            I => \N__63850\
        );

    \I__15130\ : LocalMux
    port map (
            O => \N__63855\,
            I => \N__63847\
        );

    \I__15129\ : InMux
    port map (
            O => \N__63854\,
            I => \N__63844\
        );

    \I__15128\ : CascadeMux
    port map (
            O => \N__63853\,
            I => \N__63840\
        );

    \I__15127\ : Span4Mux_v
    port map (
            O => \N__63850\,
            I => \N__63837\
        );

    \I__15126\ : Span4Mux_h
    port map (
            O => \N__63847\,
            I => \N__63834\
        );

    \I__15125\ : LocalMux
    port map (
            O => \N__63844\,
            I => \N__63831\
        );

    \I__15124\ : InMux
    port map (
            O => \N__63843\,
            I => \N__63828\
        );

    \I__15123\ : InMux
    port map (
            O => \N__63840\,
            I => \N__63825\
        );

    \I__15122\ : Span4Mux_v
    port map (
            O => \N__63837\,
            I => \N__63822\
        );

    \I__15121\ : Span4Mux_h
    port map (
            O => \N__63834\,
            I => \N__63819\
        );

    \I__15120\ : Span12Mux_h
    port map (
            O => \N__63831\,
            I => \N__63814\
        );

    \I__15119\ : LocalMux
    port map (
            O => \N__63828\,
            I => \N__63814\
        );

    \I__15118\ : LocalMux
    port map (
            O => \N__63825\,
            I => \c0.data_in_frame_12_1\
        );

    \I__15117\ : Odrv4
    port map (
            O => \N__63822\,
            I => \c0.data_in_frame_12_1\
        );

    \I__15116\ : Odrv4
    port map (
            O => \N__63819\,
            I => \c0.data_in_frame_12_1\
        );

    \I__15115\ : Odrv12
    port map (
            O => \N__63814\,
            I => \c0.data_in_frame_12_1\
        );

    \I__15114\ : InMux
    port map (
            O => \N__63805\,
            I => \N__63802\
        );

    \I__15113\ : LocalMux
    port map (
            O => \N__63802\,
            I => \c0.n7_adj_3000\
        );

    \I__15112\ : CascadeMux
    port map (
            O => \N__63799\,
            I => \N__63796\
        );

    \I__15111\ : InMux
    port map (
            O => \N__63796\,
            I => \N__63791\
        );

    \I__15110\ : InMux
    port map (
            O => \N__63795\,
            I => \N__63786\
        );

    \I__15109\ : InMux
    port map (
            O => \N__63794\,
            I => \N__63786\
        );

    \I__15108\ : LocalMux
    port map (
            O => \N__63791\,
            I => \c0.n19430\
        );

    \I__15107\ : LocalMux
    port map (
            O => \N__63786\,
            I => \c0.n19430\
        );

    \I__15106\ : CascadeMux
    port map (
            O => \N__63781\,
            I => \c0.n7_adj_3000_cascade_\
        );

    \I__15105\ : InMux
    port map (
            O => \N__63778\,
            I => \N__63771\
        );

    \I__15104\ : CascadeMux
    port map (
            O => \N__63777\,
            I => \N__63768\
        );

    \I__15103\ : InMux
    port map (
            O => \N__63776\,
            I => \N__63762\
        );

    \I__15102\ : InMux
    port map (
            O => \N__63775\,
            I => \N__63759\
        );

    \I__15101\ : InMux
    port map (
            O => \N__63774\,
            I => \N__63756\
        );

    \I__15100\ : LocalMux
    port map (
            O => \N__63771\,
            I => \N__63753\
        );

    \I__15099\ : InMux
    port map (
            O => \N__63768\,
            I => \N__63748\
        );

    \I__15098\ : InMux
    port map (
            O => \N__63767\,
            I => \N__63748\
        );

    \I__15097\ : InMux
    port map (
            O => \N__63766\,
            I => \N__63743\
        );

    \I__15096\ : InMux
    port map (
            O => \N__63765\,
            I => \N__63743\
        );

    \I__15095\ : LocalMux
    port map (
            O => \N__63762\,
            I => \N__63736\
        );

    \I__15094\ : LocalMux
    port map (
            O => \N__63759\,
            I => \N__63736\
        );

    \I__15093\ : LocalMux
    port map (
            O => \N__63756\,
            I => \N__63733\
        );

    \I__15092\ : Span4Mux_h
    port map (
            O => \N__63753\,
            I => \N__63728\
        );

    \I__15091\ : LocalMux
    port map (
            O => \N__63748\,
            I => \N__63728\
        );

    \I__15090\ : LocalMux
    port map (
            O => \N__63743\,
            I => \N__63725\
        );

    \I__15089\ : InMux
    port map (
            O => \N__63742\,
            I => \N__63720\
        );

    \I__15088\ : InMux
    port map (
            O => \N__63741\,
            I => \N__63720\
        );

    \I__15087\ : Sp12to4
    port map (
            O => \N__63736\,
            I => \N__63715\
        );

    \I__15086\ : Span12Mux_h
    port map (
            O => \N__63733\,
            I => \N__63715\
        );

    \I__15085\ : Span4Mux_h
    port map (
            O => \N__63728\,
            I => \N__63712\
        );

    \I__15084\ : Span12Mux_v
    port map (
            O => \N__63725\,
            I => \N__63709\
        );

    \I__15083\ : LocalMux
    port map (
            O => \N__63720\,
            I => data_in_frame_16_3
        );

    \I__15082\ : Odrv12
    port map (
            O => \N__63715\,
            I => data_in_frame_16_3
        );

    \I__15081\ : Odrv4
    port map (
            O => \N__63712\,
            I => data_in_frame_16_3
        );

    \I__15080\ : Odrv12
    port map (
            O => \N__63709\,
            I => data_in_frame_16_3
        );

    \I__15079\ : CascadeMux
    port map (
            O => \N__63700\,
            I => \N__63697\
        );

    \I__15078\ : InMux
    port map (
            O => \N__63697\,
            I => \N__63694\
        );

    \I__15077\ : LocalMux
    port map (
            O => \N__63694\,
            I => \N__63691\
        );

    \I__15076\ : Odrv4
    port map (
            O => \N__63691\,
            I => \c0.n6\
        );

    \I__15075\ : CascadeMux
    port map (
            O => \N__63688\,
            I => \N__63684\
        );

    \I__15074\ : InMux
    port map (
            O => \N__63687\,
            I => \N__63680\
        );

    \I__15073\ : InMux
    port map (
            O => \N__63684\,
            I => \N__63673\
        );

    \I__15072\ : InMux
    port map (
            O => \N__63683\,
            I => \N__63673\
        );

    \I__15071\ : LocalMux
    port map (
            O => \N__63680\,
            I => \N__63670\
        );

    \I__15070\ : InMux
    port map (
            O => \N__63679\,
            I => \N__63665\
        );

    \I__15069\ : InMux
    port map (
            O => \N__63678\,
            I => \N__63665\
        );

    \I__15068\ : LocalMux
    port map (
            O => \N__63673\,
            I => \N__63658\
        );

    \I__15067\ : Span4Mux_v
    port map (
            O => \N__63670\,
            I => \N__63658\
        );

    \I__15066\ : LocalMux
    port map (
            O => \N__63665\,
            I => \N__63658\
        );

    \I__15065\ : Span4Mux_h
    port map (
            O => \N__63658\,
            I => \N__63655\
        );

    \I__15064\ : Odrv4
    port map (
            O => \N__63655\,
            I => \c0.n19187\
        );

    \I__15063\ : CascadeMux
    port map (
            O => \N__63652\,
            I => \N__63648\
        );

    \I__15062\ : InMux
    port map (
            O => \N__63651\,
            I => \N__63643\
        );

    \I__15061\ : InMux
    port map (
            O => \N__63648\,
            I => \N__63640\
        );

    \I__15060\ : InMux
    port map (
            O => \N__63647\,
            I => \N__63637\
        );

    \I__15059\ : InMux
    port map (
            O => \N__63646\,
            I => \N__63634\
        );

    \I__15058\ : LocalMux
    port map (
            O => \N__63643\,
            I => \N__63631\
        );

    \I__15057\ : LocalMux
    port map (
            O => \N__63640\,
            I => \N__63622\
        );

    \I__15056\ : LocalMux
    port map (
            O => \N__63637\,
            I => \N__63622\
        );

    \I__15055\ : LocalMux
    port map (
            O => \N__63634\,
            I => \N__63619\
        );

    \I__15054\ : Span4Mux_v
    port map (
            O => \N__63631\,
            I => \N__63616\
        );

    \I__15053\ : InMux
    port map (
            O => \N__63630\,
            I => \N__63611\
        );

    \I__15052\ : InMux
    port map (
            O => \N__63629\,
            I => \N__63611\
        );

    \I__15051\ : InMux
    port map (
            O => \N__63628\,
            I => \N__63608\
        );

    \I__15050\ : InMux
    port map (
            O => \N__63627\,
            I => \N__63605\
        );

    \I__15049\ : Span4Mux_v
    port map (
            O => \N__63622\,
            I => \N__63602\
        );

    \I__15048\ : Span4Mux_v
    port map (
            O => \N__63619\,
            I => \N__63597\
        );

    \I__15047\ : Span4Mux_h
    port map (
            O => \N__63616\,
            I => \N__63597\
        );

    \I__15046\ : LocalMux
    port map (
            O => \N__63611\,
            I => \N__63590\
        );

    \I__15045\ : LocalMux
    port map (
            O => \N__63608\,
            I => \N__63590\
        );

    \I__15044\ : LocalMux
    port map (
            O => \N__63605\,
            I => \N__63590\
        );

    \I__15043\ : Odrv4
    port map (
            O => \N__63602\,
            I => \c0.n46_adj_3443\
        );

    \I__15042\ : Odrv4
    port map (
            O => \N__63597\,
            I => \c0.n46_adj_3443\
        );

    \I__15041\ : Odrv12
    port map (
            O => \N__63590\,
            I => \c0.n46_adj_3443\
        );

    \I__15040\ : CascadeMux
    port map (
            O => \N__63583\,
            I => \N__63580\
        );

    \I__15039\ : InMux
    port map (
            O => \N__63580\,
            I => \N__63577\
        );

    \I__15038\ : LocalMux
    port map (
            O => \N__63577\,
            I => \N__63570\
        );

    \I__15037\ : InMux
    port map (
            O => \N__63576\,
            I => \N__63567\
        );

    \I__15036\ : CascadeMux
    port map (
            O => \N__63575\,
            I => \N__63564\
        );

    \I__15035\ : InMux
    port map (
            O => \N__63574\,
            I => \N__63561\
        );

    \I__15034\ : CascadeMux
    port map (
            O => \N__63573\,
            I => \N__63557\
        );

    \I__15033\ : Span4Mux_v
    port map (
            O => \N__63570\,
            I => \N__63552\
        );

    \I__15032\ : LocalMux
    port map (
            O => \N__63567\,
            I => \N__63552\
        );

    \I__15031\ : InMux
    port map (
            O => \N__63564\,
            I => \N__63549\
        );

    \I__15030\ : LocalMux
    port map (
            O => \N__63561\,
            I => \N__63546\
        );

    \I__15029\ : InMux
    port map (
            O => \N__63560\,
            I => \N__63543\
        );

    \I__15028\ : InMux
    port map (
            O => \N__63557\,
            I => \N__63540\
        );

    \I__15027\ : Span4Mux_v
    port map (
            O => \N__63552\,
            I => \N__63535\
        );

    \I__15026\ : LocalMux
    port map (
            O => \N__63549\,
            I => \N__63535\
        );

    \I__15025\ : Span4Mux_v
    port map (
            O => \N__63546\,
            I => \N__63529\
        );

    \I__15024\ : LocalMux
    port map (
            O => \N__63543\,
            I => \N__63529\
        );

    \I__15023\ : LocalMux
    port map (
            O => \N__63540\,
            I => \N__63526\
        );

    \I__15022\ : Span4Mux_h
    port map (
            O => \N__63535\,
            I => \N__63523\
        );

    \I__15021\ : CascadeMux
    port map (
            O => \N__63534\,
            I => \N__63520\
        );

    \I__15020\ : Sp12to4
    port map (
            O => \N__63529\,
            I => \N__63517\
        );

    \I__15019\ : Span4Mux_h
    port map (
            O => \N__63526\,
            I => \N__63512\
        );

    \I__15018\ : Span4Mux_h
    port map (
            O => \N__63523\,
            I => \N__63512\
        );

    \I__15017\ : InMux
    port map (
            O => \N__63520\,
            I => \N__63509\
        );

    \I__15016\ : Span12Mux_h
    port map (
            O => \N__63517\,
            I => \N__63506\
        );

    \I__15015\ : Span4Mux_v
    port map (
            O => \N__63512\,
            I => \N__63503\
        );

    \I__15014\ : LocalMux
    port map (
            O => \N__63509\,
            I => \c0.data_in_frame_15_0\
        );

    \I__15013\ : Odrv12
    port map (
            O => \N__63506\,
            I => \c0.data_in_frame_15_0\
        );

    \I__15012\ : Odrv4
    port map (
            O => \N__63503\,
            I => \c0.data_in_frame_15_0\
        );

    \I__15011\ : InMux
    port map (
            O => \N__63496\,
            I => \N__63489\
        );

    \I__15010\ : InMux
    port map (
            O => \N__63495\,
            I => \N__63489\
        );

    \I__15009\ : InMux
    port map (
            O => \N__63494\,
            I => \N__63486\
        );

    \I__15008\ : LocalMux
    port map (
            O => \N__63489\,
            I => \N__63482\
        );

    \I__15007\ : LocalMux
    port map (
            O => \N__63486\,
            I => \N__63479\
        );

    \I__15006\ : InMux
    port map (
            O => \N__63485\,
            I => \N__63476\
        );

    \I__15005\ : Span4Mux_v
    port map (
            O => \N__63482\,
            I => \N__63473\
        );

    \I__15004\ : Span4Mux_v
    port map (
            O => \N__63479\,
            I => \N__63468\
        );

    \I__15003\ : LocalMux
    port map (
            O => \N__63476\,
            I => \N__63468\
        );

    \I__15002\ : Sp12to4
    port map (
            O => \N__63473\,
            I => \N__63465\
        );

    \I__15001\ : Span4Mux_h
    port map (
            O => \N__63468\,
            I => \N__63462\
        );

    \I__15000\ : Odrv12
    port map (
            O => \N__63465\,
            I => \c0.n40_adj_3413\
        );

    \I__14999\ : Odrv4
    port map (
            O => \N__63462\,
            I => \c0.n40_adj_3413\
        );

    \I__14998\ : CascadeMux
    port map (
            O => \N__63457\,
            I => \N__63452\
        );

    \I__14997\ : CascadeMux
    port map (
            O => \N__63456\,
            I => \N__63449\
        );

    \I__14996\ : InMux
    port map (
            O => \N__63455\,
            I => \N__63446\
        );

    \I__14995\ : InMux
    port map (
            O => \N__63452\,
            I => \N__63441\
        );

    \I__14994\ : InMux
    port map (
            O => \N__63449\,
            I => \N__63441\
        );

    \I__14993\ : LocalMux
    port map (
            O => \N__63446\,
            I => \N__63438\
        );

    \I__14992\ : LocalMux
    port map (
            O => \N__63441\,
            I => \N__63435\
        );

    \I__14991\ : Sp12to4
    port map (
            O => \N__63438\,
            I => \N__63432\
        );

    \I__14990\ : Span4Mux_h
    port map (
            O => \N__63435\,
            I => \N__63429\
        );

    \I__14989\ : Span12Mux_v
    port map (
            O => \N__63432\,
            I => \N__63426\
        );

    \I__14988\ : Span4Mux_v
    port map (
            O => \N__63429\,
            I => \N__63423\
        );

    \I__14987\ : Odrv12
    port map (
            O => \N__63426\,
            I => \c0.n45_adj_3138\
        );

    \I__14986\ : Odrv4
    port map (
            O => \N__63423\,
            I => \c0.n45_adj_3138\
        );

    \I__14985\ : InMux
    port map (
            O => \N__63418\,
            I => \N__63409\
        );

    \I__14984\ : InMux
    port map (
            O => \N__63417\,
            I => \N__63404\
        );

    \I__14983\ : InMux
    port map (
            O => \N__63416\,
            I => \N__63404\
        );

    \I__14982\ : InMux
    port map (
            O => \N__63415\,
            I => \N__63399\
        );

    \I__14981\ : InMux
    port map (
            O => \N__63414\,
            I => \N__63399\
        );

    \I__14980\ : InMux
    port map (
            O => \N__63413\,
            I => \N__63396\
        );

    \I__14979\ : InMux
    port map (
            O => \N__63412\,
            I => \N__63391\
        );

    \I__14978\ : LocalMux
    port map (
            O => \N__63409\,
            I => \N__63386\
        );

    \I__14977\ : LocalMux
    port map (
            O => \N__63404\,
            I => \N__63381\
        );

    \I__14976\ : LocalMux
    port map (
            O => \N__63399\,
            I => \N__63381\
        );

    \I__14975\ : LocalMux
    port map (
            O => \N__63396\,
            I => \N__63374\
        );

    \I__14974\ : InMux
    port map (
            O => \N__63395\,
            I => \N__63371\
        );

    \I__14973\ : InMux
    port map (
            O => \N__63394\,
            I => \N__63368\
        );

    \I__14972\ : LocalMux
    port map (
            O => \N__63391\,
            I => \N__63365\
        );

    \I__14971\ : CascadeMux
    port map (
            O => \N__63390\,
            I => \N__63362\
        );

    \I__14970\ : CascadeMux
    port map (
            O => \N__63389\,
            I => \N__63359\
        );

    \I__14969\ : Span4Mux_v
    port map (
            O => \N__63386\,
            I => \N__63348\
        );

    \I__14968\ : Span4Mux_v
    port map (
            O => \N__63381\,
            I => \N__63348\
        );

    \I__14967\ : InMux
    port map (
            O => \N__63380\,
            I => \N__63343\
        );

    \I__14966\ : InMux
    port map (
            O => \N__63379\,
            I => \N__63343\
        );

    \I__14965\ : InMux
    port map (
            O => \N__63378\,
            I => \N__63340\
        );

    \I__14964\ : InMux
    port map (
            O => \N__63377\,
            I => \N__63337\
        );

    \I__14963\ : Span4Mux_h
    port map (
            O => \N__63374\,
            I => \N__63334\
        );

    \I__14962\ : LocalMux
    port map (
            O => \N__63371\,
            I => \N__63331\
        );

    \I__14961\ : LocalMux
    port map (
            O => \N__63368\,
            I => \N__63328\
        );

    \I__14960\ : Span4Mux_v
    port map (
            O => \N__63365\,
            I => \N__63325\
        );

    \I__14959\ : InMux
    port map (
            O => \N__63362\,
            I => \N__63318\
        );

    \I__14958\ : InMux
    port map (
            O => \N__63359\,
            I => \N__63318\
        );

    \I__14957\ : InMux
    port map (
            O => \N__63358\,
            I => \N__63318\
        );

    \I__14956\ : InMux
    port map (
            O => \N__63357\,
            I => \N__63315\
        );

    \I__14955\ : InMux
    port map (
            O => \N__63356\,
            I => \N__63312\
        );

    \I__14954\ : InMux
    port map (
            O => \N__63355\,
            I => \N__63305\
        );

    \I__14953\ : InMux
    port map (
            O => \N__63354\,
            I => \N__63305\
        );

    \I__14952\ : InMux
    port map (
            O => \N__63353\,
            I => \N__63305\
        );

    \I__14951\ : Span4Mux_h
    port map (
            O => \N__63348\,
            I => \N__63300\
        );

    \I__14950\ : LocalMux
    port map (
            O => \N__63343\,
            I => \N__63300\
        );

    \I__14949\ : LocalMux
    port map (
            O => \N__63340\,
            I => \N__63295\
        );

    \I__14948\ : LocalMux
    port map (
            O => \N__63337\,
            I => \N__63295\
        );

    \I__14947\ : Span4Mux_h
    port map (
            O => \N__63334\,
            I => \N__63292\
        );

    \I__14946\ : Span4Mux_h
    port map (
            O => \N__63331\,
            I => \N__63287\
        );

    \I__14945\ : Span4Mux_h
    port map (
            O => \N__63328\,
            I => \N__63287\
        );

    \I__14944\ : Sp12to4
    port map (
            O => \N__63325\,
            I => \N__63282\
        );

    \I__14943\ : LocalMux
    port map (
            O => \N__63318\,
            I => \N__63282\
        );

    \I__14942\ : LocalMux
    port map (
            O => \N__63315\,
            I => \N__63273\
        );

    \I__14941\ : LocalMux
    port map (
            O => \N__63312\,
            I => \N__63273\
        );

    \I__14940\ : LocalMux
    port map (
            O => \N__63305\,
            I => \N__63273\
        );

    \I__14939\ : Span4Mux_v
    port map (
            O => \N__63300\,
            I => \N__63270\
        );

    \I__14938\ : Span12Mux_h
    port map (
            O => \N__63295\,
            I => \N__63265\
        );

    \I__14937\ : Sp12to4
    port map (
            O => \N__63292\,
            I => \N__63265\
        );

    \I__14936\ : Sp12to4
    port map (
            O => \N__63287\,
            I => \N__63260\
        );

    \I__14935\ : Span12Mux_h
    port map (
            O => \N__63282\,
            I => \N__63260\
        );

    \I__14934\ : InMux
    port map (
            O => \N__63281\,
            I => \N__63257\
        );

    \I__14933\ : InMux
    port map (
            O => \N__63280\,
            I => \N__63254\
        );

    \I__14932\ : Span4Mux_v
    port map (
            O => \N__63273\,
            I => \N__63251\
        );

    \I__14931\ : Sp12to4
    port map (
            O => \N__63270\,
            I => \N__63246\
        );

    \I__14930\ : Span12Mux_v
    port map (
            O => \N__63265\,
            I => \N__63246\
        );

    \I__14929\ : Span12Mux_v
    port map (
            O => \N__63260\,
            I => \N__63243\
        );

    \I__14928\ : LocalMux
    port map (
            O => \N__63257\,
            I => \c0.n19115\
        );

    \I__14927\ : LocalMux
    port map (
            O => \N__63254\,
            I => \c0.n19115\
        );

    \I__14926\ : Odrv4
    port map (
            O => \N__63251\,
            I => \c0.n19115\
        );

    \I__14925\ : Odrv12
    port map (
            O => \N__63246\,
            I => \c0.n19115\
        );

    \I__14924\ : Odrv12
    port map (
            O => \N__63243\,
            I => \c0.n19115\
        );

    \I__14923\ : InMux
    port map (
            O => \N__63232\,
            I => \N__63228\
        );

    \I__14922\ : InMux
    port map (
            O => \N__63231\,
            I => \N__63225\
        );

    \I__14921\ : LocalMux
    port map (
            O => \N__63228\,
            I => \N__63219\
        );

    \I__14920\ : LocalMux
    port map (
            O => \N__63225\,
            I => \N__63219\
        );

    \I__14919\ : InMux
    port map (
            O => \N__63224\,
            I => \N__63215\
        );

    \I__14918\ : Span4Mux_h
    port map (
            O => \N__63219\,
            I => \N__63212\
        );

    \I__14917\ : InMux
    port map (
            O => \N__63218\,
            I => \N__63209\
        );

    \I__14916\ : LocalMux
    port map (
            O => \N__63215\,
            I => \c0.data_in_frame_9_3\
        );

    \I__14915\ : Odrv4
    port map (
            O => \N__63212\,
            I => \c0.data_in_frame_9_3\
        );

    \I__14914\ : LocalMux
    port map (
            O => \N__63209\,
            I => \c0.data_in_frame_9_3\
        );

    \I__14913\ : InMux
    port map (
            O => \N__63202\,
            I => \N__63198\
        );

    \I__14912\ : InMux
    port map (
            O => \N__63201\,
            I => \N__63194\
        );

    \I__14911\ : LocalMux
    port map (
            O => \N__63198\,
            I => \N__63191\
        );

    \I__14910\ : InMux
    port map (
            O => \N__63197\,
            I => \N__63188\
        );

    \I__14909\ : LocalMux
    port map (
            O => \N__63194\,
            I => \c0.data_in_frame_11_5\
        );

    \I__14908\ : Odrv12
    port map (
            O => \N__63191\,
            I => \c0.data_in_frame_11_5\
        );

    \I__14907\ : LocalMux
    port map (
            O => \N__63188\,
            I => \c0.data_in_frame_11_5\
        );

    \I__14906\ : InMux
    port map (
            O => \N__63181\,
            I => \N__63175\
        );

    \I__14905\ : InMux
    port map (
            O => \N__63180\,
            I => \N__63175\
        );

    \I__14904\ : LocalMux
    port map (
            O => \N__63175\,
            I => \N__63172\
        );

    \I__14903\ : Span12Mux_h
    port map (
            O => \N__63172\,
            I => \N__63169\
        );

    \I__14902\ : Odrv12
    port map (
            O => \N__63169\,
            I => \c0.n5_adj_3043\
        );

    \I__14901\ : CascadeMux
    port map (
            O => \N__63166\,
            I => \N__63163\
        );

    \I__14900\ : InMux
    port map (
            O => \N__63163\,
            I => \N__63159\
        );

    \I__14899\ : InMux
    port map (
            O => \N__63162\,
            I => \N__63156\
        );

    \I__14898\ : LocalMux
    port map (
            O => \N__63159\,
            I => \N__63150\
        );

    \I__14897\ : LocalMux
    port map (
            O => \N__63156\,
            I => \N__63150\
        );

    \I__14896\ : InMux
    port map (
            O => \N__63155\,
            I => \N__63145\
        );

    \I__14895\ : Span4Mux_v
    port map (
            O => \N__63150\,
            I => \N__63142\
        );

    \I__14894\ : CascadeMux
    port map (
            O => \N__63149\,
            I => \N__63139\
        );

    \I__14893\ : CascadeMux
    port map (
            O => \N__63148\,
            I => \N__63136\
        );

    \I__14892\ : LocalMux
    port map (
            O => \N__63145\,
            I => \N__63132\
        );

    \I__14891\ : Span4Mux_h
    port map (
            O => \N__63142\,
            I => \N__63129\
        );

    \I__14890\ : InMux
    port map (
            O => \N__63139\,
            I => \N__63124\
        );

    \I__14889\ : InMux
    port map (
            O => \N__63136\,
            I => \N__63124\
        );

    \I__14888\ : InMux
    port map (
            O => \N__63135\,
            I => \N__63121\
        );

    \I__14887\ : Span12Mux_v
    port map (
            O => \N__63132\,
            I => \N__63118\
        );

    \I__14886\ : Odrv4
    port map (
            O => \N__63129\,
            I => \c0.data_in_frame_7_1\
        );

    \I__14885\ : LocalMux
    port map (
            O => \N__63124\,
            I => \c0.data_in_frame_7_1\
        );

    \I__14884\ : LocalMux
    port map (
            O => \N__63121\,
            I => \c0.data_in_frame_7_1\
        );

    \I__14883\ : Odrv12
    port map (
            O => \N__63118\,
            I => \c0.data_in_frame_7_1\
        );

    \I__14882\ : InMux
    port map (
            O => \N__63109\,
            I => \N__63106\
        );

    \I__14881\ : LocalMux
    port map (
            O => \N__63106\,
            I => \N__63101\
        );

    \I__14880\ : InMux
    port map (
            O => \N__63105\,
            I => \N__63096\
        );

    \I__14879\ : InMux
    port map (
            O => \N__63104\,
            I => \N__63093\
        );

    \I__14878\ : Span4Mux_h
    port map (
            O => \N__63101\,
            I => \N__63090\
        );

    \I__14877\ : InMux
    port map (
            O => \N__63100\,
            I => \N__63087\
        );

    \I__14876\ : InMux
    port map (
            O => \N__63099\,
            I => \N__63084\
        );

    \I__14875\ : LocalMux
    port map (
            O => \N__63096\,
            I => \N__63081\
        );

    \I__14874\ : LocalMux
    port map (
            O => \N__63093\,
            I => \c0.data_in_frame_9_0\
        );

    \I__14873\ : Odrv4
    port map (
            O => \N__63090\,
            I => \c0.data_in_frame_9_0\
        );

    \I__14872\ : LocalMux
    port map (
            O => \N__63087\,
            I => \c0.data_in_frame_9_0\
        );

    \I__14871\ : LocalMux
    port map (
            O => \N__63084\,
            I => \c0.data_in_frame_9_0\
        );

    \I__14870\ : Odrv12
    port map (
            O => \N__63081\,
            I => \c0.data_in_frame_9_0\
        );

    \I__14869\ : CascadeMux
    port map (
            O => \N__63070\,
            I => \N__63067\
        );

    \I__14868\ : InMux
    port map (
            O => \N__63067\,
            I => \N__63062\
        );

    \I__14867\ : InMux
    port map (
            O => \N__63066\,
            I => \N__63057\
        );

    \I__14866\ : InMux
    port map (
            O => \N__63065\,
            I => \N__63057\
        );

    \I__14865\ : LocalMux
    port map (
            O => \N__63062\,
            I => \N__63054\
        );

    \I__14864\ : LocalMux
    port map (
            O => \N__63057\,
            I => \c0.data_in_frame_11_3\
        );

    \I__14863\ : Odrv12
    port map (
            O => \N__63054\,
            I => \c0.data_in_frame_11_3\
        );

    \I__14862\ : InMux
    port map (
            O => \N__63049\,
            I => \N__63045\
        );

    \I__14861\ : CascadeMux
    port map (
            O => \N__63048\,
            I => \N__63041\
        );

    \I__14860\ : LocalMux
    port map (
            O => \N__63045\,
            I => \N__63038\
        );

    \I__14859\ : InMux
    port map (
            O => \N__63044\,
            I => \N__63035\
        );

    \I__14858\ : InMux
    port map (
            O => \N__63041\,
            I => \N__63031\
        );

    \I__14857\ : Span4Mux_v
    port map (
            O => \N__63038\,
            I => \N__63028\
        );

    \I__14856\ : LocalMux
    port map (
            O => \N__63035\,
            I => \N__63025\
        );

    \I__14855\ : InMux
    port map (
            O => \N__63034\,
            I => \N__63022\
        );

    \I__14854\ : LocalMux
    port map (
            O => \N__63031\,
            I => \c0.data_in_frame_13_4\
        );

    \I__14853\ : Odrv4
    port map (
            O => \N__63028\,
            I => \c0.data_in_frame_13_4\
        );

    \I__14852\ : Odrv4
    port map (
            O => \N__63025\,
            I => \c0.data_in_frame_13_4\
        );

    \I__14851\ : LocalMux
    port map (
            O => \N__63022\,
            I => \c0.data_in_frame_13_4\
        );

    \I__14850\ : CascadeMux
    port map (
            O => \N__63013\,
            I => \N__63010\
        );

    \I__14849\ : InMux
    port map (
            O => \N__63010\,
            I => \N__63007\
        );

    \I__14848\ : LocalMux
    port map (
            O => \N__63007\,
            I => \N__63004\
        );

    \I__14847\ : Span4Mux_v
    port map (
            O => \N__63004\,
            I => \N__63001\
        );

    \I__14846\ : Span4Mux_h
    port map (
            O => \N__63001\,
            I => \N__62998\
        );

    \I__14845\ : Odrv4
    port map (
            O => \N__62998\,
            I => \c0.n11_adj_3492\
        );

    \I__14844\ : CascadeMux
    port map (
            O => \N__62995\,
            I => \c0.n11_adj_3492_cascade_\
        );

    \I__14843\ : InMux
    port map (
            O => \N__62992\,
            I => \N__62989\
        );

    \I__14842\ : LocalMux
    port map (
            O => \N__62989\,
            I => \N__62985\
        );

    \I__14841\ : InMux
    port map (
            O => \N__62988\,
            I => \N__62982\
        );

    \I__14840\ : Span4Mux_v
    port map (
            O => \N__62985\,
            I => \N__62976\
        );

    \I__14839\ : LocalMux
    port map (
            O => \N__62982\,
            I => \N__62976\
        );

    \I__14838\ : InMux
    port map (
            O => \N__62981\,
            I => \N__62973\
        );

    \I__14837\ : Span4Mux_h
    port map (
            O => \N__62976\,
            I => \N__62970\
        );

    \I__14836\ : LocalMux
    port map (
            O => \N__62973\,
            I => \N__62965\
        );

    \I__14835\ : Span4Mux_h
    port map (
            O => \N__62970\,
            I => \N__62962\
        );

    \I__14834\ : InMux
    port map (
            O => \N__62969\,
            I => \N__62957\
        );

    \I__14833\ : InMux
    port map (
            O => \N__62968\,
            I => \N__62957\
        );

    \I__14832\ : Odrv4
    port map (
            O => \N__62965\,
            I => data_in_frame_16_0
        );

    \I__14831\ : Odrv4
    port map (
            O => \N__62962\,
            I => data_in_frame_16_0
        );

    \I__14830\ : LocalMux
    port map (
            O => \N__62957\,
            I => data_in_frame_16_0
        );

    \I__14829\ : InMux
    port map (
            O => \N__62950\,
            I => \N__62947\
        );

    \I__14828\ : LocalMux
    port map (
            O => \N__62947\,
            I => \N__62944\
        );

    \I__14827\ : Span4Mux_h
    port map (
            O => \N__62944\,
            I => \N__62941\
        );

    \I__14826\ : Span4Mux_v
    port map (
            O => \N__62941\,
            I => \N__62938\
        );

    \I__14825\ : Odrv4
    port map (
            O => \N__62938\,
            I => \c0.n20_adj_3527\
        );

    \I__14824\ : InMux
    port map (
            O => \N__62935\,
            I => \N__62931\
        );

    \I__14823\ : CascadeMux
    port map (
            O => \N__62934\,
            I => \N__62928\
        );

    \I__14822\ : LocalMux
    port map (
            O => \N__62931\,
            I => \N__62923\
        );

    \I__14821\ : InMux
    port map (
            O => \N__62928\,
            I => \N__62916\
        );

    \I__14820\ : InMux
    port map (
            O => \N__62927\,
            I => \N__62916\
        );

    \I__14819\ : InMux
    port map (
            O => \N__62926\,
            I => \N__62916\
        );

    \I__14818\ : Odrv4
    port map (
            O => \N__62923\,
            I => \c0.data_in_frame_11_1\
        );

    \I__14817\ : LocalMux
    port map (
            O => \N__62916\,
            I => \c0.data_in_frame_11_1\
        );

    \I__14816\ : InMux
    port map (
            O => \N__62911\,
            I => \N__62908\
        );

    \I__14815\ : LocalMux
    port map (
            O => \N__62908\,
            I => \N__62905\
        );

    \I__14814\ : Span4Mux_h
    port map (
            O => \N__62905\,
            I => \N__62901\
        );

    \I__14813\ : InMux
    port map (
            O => \N__62904\,
            I => \N__62898\
        );

    \I__14812\ : Span4Mux_h
    port map (
            O => \N__62901\,
            I => \N__62895\
        );

    \I__14811\ : LocalMux
    port map (
            O => \N__62898\,
            I => \c0.n19229\
        );

    \I__14810\ : Odrv4
    port map (
            O => \N__62895\,
            I => \c0.n19229\
        );

    \I__14809\ : InMux
    port map (
            O => \N__62890\,
            I => \N__62886\
        );

    \I__14808\ : InMux
    port map (
            O => \N__62889\,
            I => \N__62882\
        );

    \I__14807\ : LocalMux
    port map (
            O => \N__62886\,
            I => \N__62879\
        );

    \I__14806\ : CascadeMux
    port map (
            O => \N__62885\,
            I => \N__62875\
        );

    \I__14805\ : LocalMux
    port map (
            O => \N__62882\,
            I => \N__62872\
        );

    \I__14804\ : Span4Mux_v
    port map (
            O => \N__62879\,
            I => \N__62869\
        );

    \I__14803\ : CascadeMux
    port map (
            O => \N__62878\,
            I => \N__62866\
        );

    \I__14802\ : InMux
    port map (
            O => \N__62875\,
            I => \N__62863\
        );

    \I__14801\ : Span4Mux_v
    port map (
            O => \N__62872\,
            I => \N__62858\
        );

    \I__14800\ : Span4Mux_h
    port map (
            O => \N__62869\,
            I => \N__62858\
        );

    \I__14799\ : InMux
    port map (
            O => \N__62866\,
            I => \N__62855\
        );

    \I__14798\ : LocalMux
    port map (
            O => \N__62863\,
            I => \c0.data_in_frame_11_2\
        );

    \I__14797\ : Odrv4
    port map (
            O => \N__62858\,
            I => \c0.data_in_frame_11_2\
        );

    \I__14796\ : LocalMux
    port map (
            O => \N__62855\,
            I => \c0.data_in_frame_11_2\
        );

    \I__14795\ : InMux
    port map (
            O => \N__62848\,
            I => \N__62839\
        );

    \I__14794\ : InMux
    port map (
            O => \N__62847\,
            I => \N__62839\
        );

    \I__14793\ : InMux
    port map (
            O => \N__62846\,
            I => \N__62834\
        );

    \I__14792\ : InMux
    port map (
            O => \N__62845\,
            I => \N__62831\
        );

    \I__14791\ : InMux
    port map (
            O => \N__62844\,
            I => \N__62827\
        );

    \I__14790\ : LocalMux
    port map (
            O => \N__62839\,
            I => \N__62824\
        );

    \I__14789\ : InMux
    port map (
            O => \N__62838\,
            I => \N__62819\
        );

    \I__14788\ : InMux
    port map (
            O => \N__62837\,
            I => \N__62819\
        );

    \I__14787\ : LocalMux
    port map (
            O => \N__62834\,
            I => \N__62816\
        );

    \I__14786\ : LocalMux
    port map (
            O => \N__62831\,
            I => \N__62813\
        );

    \I__14785\ : InMux
    port map (
            O => \N__62830\,
            I => \N__62807\
        );

    \I__14784\ : LocalMux
    port map (
            O => \N__62827\,
            I => \N__62804\
        );

    \I__14783\ : Span4Mux_v
    port map (
            O => \N__62824\,
            I => \N__62798\
        );

    \I__14782\ : LocalMux
    port map (
            O => \N__62819\,
            I => \N__62795\
        );

    \I__14781\ : Span4Mux_v
    port map (
            O => \N__62816\,
            I => \N__62788\
        );

    \I__14780\ : Span4Mux_v
    port map (
            O => \N__62813\,
            I => \N__62788\
        );

    \I__14779\ : InMux
    port map (
            O => \N__62812\,
            I => \N__62785\
        );

    \I__14778\ : InMux
    port map (
            O => \N__62811\,
            I => \N__62782\
        );

    \I__14777\ : InMux
    port map (
            O => \N__62810\,
            I => \N__62779\
        );

    \I__14776\ : LocalMux
    port map (
            O => \N__62807\,
            I => \N__62774\
        );

    \I__14775\ : Span4Mux_v
    port map (
            O => \N__62804\,
            I => \N__62774\
        );

    \I__14774\ : InMux
    port map (
            O => \N__62803\,
            I => \N__62771\
        );

    \I__14773\ : InMux
    port map (
            O => \N__62802\,
            I => \N__62766\
        );

    \I__14772\ : InMux
    port map (
            O => \N__62801\,
            I => \N__62766\
        );

    \I__14771\ : Sp12to4
    port map (
            O => \N__62798\,
            I => \N__62763\
        );

    \I__14770\ : Sp12to4
    port map (
            O => \N__62795\,
            I => \N__62760\
        );

    \I__14769\ : InMux
    port map (
            O => \N__62794\,
            I => \N__62755\
        );

    \I__14768\ : InMux
    port map (
            O => \N__62793\,
            I => \N__62755\
        );

    \I__14767\ : Sp12to4
    port map (
            O => \N__62788\,
            I => \N__62752\
        );

    \I__14766\ : LocalMux
    port map (
            O => \N__62785\,
            I => \N__62743\
        );

    \I__14765\ : LocalMux
    port map (
            O => \N__62782\,
            I => \N__62743\
        );

    \I__14764\ : LocalMux
    port map (
            O => \N__62779\,
            I => \N__62743\
        );

    \I__14763\ : Sp12to4
    port map (
            O => \N__62774\,
            I => \N__62743\
        );

    \I__14762\ : LocalMux
    port map (
            O => \N__62771\,
            I => \N__62734\
        );

    \I__14761\ : LocalMux
    port map (
            O => \N__62766\,
            I => \N__62734\
        );

    \I__14760\ : Span12Mux_h
    port map (
            O => \N__62763\,
            I => \N__62734\
        );

    \I__14759\ : Span12Mux_s11_v
    port map (
            O => \N__62760\,
            I => \N__62734\
        );

    \I__14758\ : LocalMux
    port map (
            O => \N__62755\,
            I => \c0.n19134\
        );

    \I__14757\ : Odrv12
    port map (
            O => \N__62752\,
            I => \c0.n19134\
        );

    \I__14756\ : Odrv12
    port map (
            O => \N__62743\,
            I => \c0.n19134\
        );

    \I__14755\ : Odrv12
    port map (
            O => \N__62734\,
            I => \c0.n19134\
        );

    \I__14754\ : CascadeMux
    port map (
            O => \N__62725\,
            I => \N__62721\
        );

    \I__14753\ : CascadeMux
    port map (
            O => \N__62724\,
            I => \N__62717\
        );

    \I__14752\ : InMux
    port map (
            O => \N__62721\,
            I => \N__62713\
        );

    \I__14751\ : InMux
    port map (
            O => \N__62720\,
            I => \N__62710\
        );

    \I__14750\ : InMux
    port map (
            O => \N__62717\,
            I => \N__62705\
        );

    \I__14749\ : InMux
    port map (
            O => \N__62716\,
            I => \N__62705\
        );

    \I__14748\ : LocalMux
    port map (
            O => \N__62713\,
            I => \c0.data_in_frame_10_7\
        );

    \I__14747\ : LocalMux
    port map (
            O => \N__62710\,
            I => \c0.data_in_frame_10_7\
        );

    \I__14746\ : LocalMux
    port map (
            O => \N__62705\,
            I => \c0.data_in_frame_10_7\
        );

    \I__14745\ : CascadeMux
    port map (
            O => \N__62698\,
            I => \N__62695\
        );

    \I__14744\ : InMux
    port map (
            O => \N__62695\,
            I => \N__62692\
        );

    \I__14743\ : LocalMux
    port map (
            O => \N__62692\,
            I => \N__62689\
        );

    \I__14742\ : Span4Mux_h
    port map (
            O => \N__62689\,
            I => \N__62686\
        );

    \I__14741\ : Odrv4
    port map (
            O => \N__62686\,
            I => \c0.n6_adj_3037\
        );

    \I__14740\ : InMux
    port map (
            O => \N__62683\,
            I => \N__62676\
        );

    \I__14739\ : InMux
    port map (
            O => \N__62682\,
            I => \N__62673\
        );

    \I__14738\ : CascadeMux
    port map (
            O => \N__62681\,
            I => \N__62670\
        );

    \I__14737\ : InMux
    port map (
            O => \N__62680\,
            I => \N__62667\
        );

    \I__14736\ : InMux
    port map (
            O => \N__62679\,
            I => \N__62664\
        );

    \I__14735\ : LocalMux
    port map (
            O => \N__62676\,
            I => \N__62659\
        );

    \I__14734\ : LocalMux
    port map (
            O => \N__62673\,
            I => \N__62659\
        );

    \I__14733\ : InMux
    port map (
            O => \N__62670\,
            I => \N__62655\
        );

    \I__14732\ : LocalMux
    port map (
            O => \N__62667\,
            I => \N__62650\
        );

    \I__14731\ : LocalMux
    port map (
            O => \N__62664\,
            I => \N__62650\
        );

    \I__14730\ : Span12Mux_v
    port map (
            O => \N__62659\,
            I => \N__62647\
        );

    \I__14729\ : InMux
    port map (
            O => \N__62658\,
            I => \N__62644\
        );

    \I__14728\ : LocalMux
    port map (
            O => \N__62655\,
            I => \c0.data_in_frame_5_7\
        );

    \I__14727\ : Odrv12
    port map (
            O => \N__62650\,
            I => \c0.data_in_frame_5_7\
        );

    \I__14726\ : Odrv12
    port map (
            O => \N__62647\,
            I => \c0.data_in_frame_5_7\
        );

    \I__14725\ : LocalMux
    port map (
            O => \N__62644\,
            I => \c0.data_in_frame_5_7\
        );

    \I__14724\ : InMux
    port map (
            O => \N__62635\,
            I => \N__62632\
        );

    \I__14723\ : LocalMux
    port map (
            O => \N__62632\,
            I => \c0.n4_adj_3036\
        );

    \I__14722\ : CascadeMux
    port map (
            O => \N__62629\,
            I => \c0.n6_adj_3037_cascade_\
        );

    \I__14721\ : CascadeMux
    port map (
            O => \N__62626\,
            I => \N__62621\
        );

    \I__14720\ : InMux
    port map (
            O => \N__62625\,
            I => \N__62615\
        );

    \I__14719\ : InMux
    port map (
            O => \N__62624\,
            I => \N__62612\
        );

    \I__14718\ : InMux
    port map (
            O => \N__62621\,
            I => \N__62609\
        );

    \I__14717\ : InMux
    port map (
            O => \N__62620\,
            I => \N__62606\
        );

    \I__14716\ : InMux
    port map (
            O => \N__62619\,
            I => \N__62601\
        );

    \I__14715\ : InMux
    port map (
            O => \N__62618\,
            I => \N__62601\
        );

    \I__14714\ : LocalMux
    port map (
            O => \N__62615\,
            I => \N__62596\
        );

    \I__14713\ : LocalMux
    port map (
            O => \N__62612\,
            I => \N__62596\
        );

    \I__14712\ : LocalMux
    port map (
            O => \N__62609\,
            I => \c0.data_in_frame_3_5\
        );

    \I__14711\ : LocalMux
    port map (
            O => \N__62606\,
            I => \c0.data_in_frame_3_5\
        );

    \I__14710\ : LocalMux
    port map (
            O => \N__62601\,
            I => \c0.data_in_frame_3_5\
        );

    \I__14709\ : Odrv4
    port map (
            O => \N__62596\,
            I => \c0.data_in_frame_3_5\
        );

    \I__14708\ : InMux
    port map (
            O => \N__62587\,
            I => \N__62584\
        );

    \I__14707\ : LocalMux
    port map (
            O => \N__62584\,
            I => \N__62579\
        );

    \I__14706\ : InMux
    port map (
            O => \N__62583\,
            I => \N__62576\
        );

    \I__14705\ : InMux
    port map (
            O => \N__62582\,
            I => \N__62573\
        );

    \I__14704\ : Span4Mux_h
    port map (
            O => \N__62579\,
            I => \N__62570\
        );

    \I__14703\ : LocalMux
    port map (
            O => \N__62576\,
            I => \N__62567\
        );

    \I__14702\ : LocalMux
    port map (
            O => \N__62573\,
            I => \N__62564\
        );

    \I__14701\ : Span4Mux_h
    port map (
            O => \N__62570\,
            I => \N__62561\
        );

    \I__14700\ : Span4Mux_h
    port map (
            O => \N__62567\,
            I => \N__62556\
        );

    \I__14699\ : Span4Mux_h
    port map (
            O => \N__62564\,
            I => \N__62556\
        );

    \I__14698\ : Odrv4
    port map (
            O => \N__62561\,
            I => \c0.n19560\
        );

    \I__14697\ : Odrv4
    port map (
            O => \N__62556\,
            I => \c0.n19560\
        );

    \I__14696\ : CascadeMux
    port map (
            O => \N__62551\,
            I => \N__62548\
        );

    \I__14695\ : InMux
    port map (
            O => \N__62548\,
            I => \N__62545\
        );

    \I__14694\ : LocalMux
    port map (
            O => \N__62545\,
            I => \N__62541\
        );

    \I__14693\ : CascadeMux
    port map (
            O => \N__62544\,
            I => \N__62538\
        );

    \I__14692\ : Span4Mux_v
    port map (
            O => \N__62541\,
            I => \N__62535\
        );

    \I__14691\ : InMux
    port map (
            O => \N__62538\,
            I => \N__62532\
        );

    \I__14690\ : Odrv4
    port map (
            O => \N__62535\,
            I => \c0.data_out_frame_0__7__N_1540\
        );

    \I__14689\ : LocalMux
    port map (
            O => \N__62532\,
            I => \c0.data_out_frame_0__7__N_1540\
        );

    \I__14688\ : InMux
    port map (
            O => \N__62527\,
            I => \N__62524\
        );

    \I__14687\ : LocalMux
    port map (
            O => \N__62524\,
            I => \N__62519\
        );

    \I__14686\ : InMux
    port map (
            O => \N__62523\,
            I => \N__62516\
        );

    \I__14685\ : CascadeMux
    port map (
            O => \N__62522\,
            I => \N__62513\
        );

    \I__14684\ : Span4Mux_v
    port map (
            O => \N__62519\,
            I => \N__62507\
        );

    \I__14683\ : LocalMux
    port map (
            O => \N__62516\,
            I => \N__62507\
        );

    \I__14682\ : InMux
    port map (
            O => \N__62513\,
            I => \N__62502\
        );

    \I__14681\ : InMux
    port map (
            O => \N__62512\,
            I => \N__62502\
        );

    \I__14680\ : Odrv4
    port map (
            O => \N__62507\,
            I => \c0.data_in_frame_6_6\
        );

    \I__14679\ : LocalMux
    port map (
            O => \N__62502\,
            I => \c0.data_in_frame_6_6\
        );

    \I__14678\ : InMux
    port map (
            O => \N__62497\,
            I => \N__62492\
        );

    \I__14677\ : CascadeMux
    port map (
            O => \N__62496\,
            I => \N__62489\
        );

    \I__14676\ : InMux
    port map (
            O => \N__62495\,
            I => \N__62486\
        );

    \I__14675\ : LocalMux
    port map (
            O => \N__62492\,
            I => \N__62483\
        );

    \I__14674\ : InMux
    port map (
            O => \N__62489\,
            I => \N__62480\
        );

    \I__14673\ : LocalMux
    port map (
            O => \N__62486\,
            I => \N__62477\
        );

    \I__14672\ : Span4Mux_v
    port map (
            O => \N__62483\,
            I => \N__62474\
        );

    \I__14671\ : LocalMux
    port map (
            O => \N__62480\,
            I => \c0.n19258\
        );

    \I__14670\ : Odrv4
    port map (
            O => \N__62477\,
            I => \c0.n19258\
        );

    \I__14669\ : Odrv4
    port map (
            O => \N__62474\,
            I => \c0.n19258\
        );

    \I__14668\ : InMux
    port map (
            O => \N__62467\,
            I => \N__62461\
        );

    \I__14667\ : InMux
    port map (
            O => \N__62466\,
            I => \N__62456\
        );

    \I__14666\ : InMux
    port map (
            O => \N__62465\,
            I => \N__62456\
        );

    \I__14665\ : CascadeMux
    port map (
            O => \N__62464\,
            I => \N__62453\
        );

    \I__14664\ : LocalMux
    port map (
            O => \N__62461\,
            I => \N__62448\
        );

    \I__14663\ : LocalMux
    port map (
            O => \N__62456\,
            I => \N__62448\
        );

    \I__14662\ : InMux
    port map (
            O => \N__62453\,
            I => \N__62444\
        );

    \I__14661\ : Span4Mux_v
    port map (
            O => \N__62448\,
            I => \N__62441\
        );

    \I__14660\ : InMux
    port map (
            O => \N__62447\,
            I => \N__62437\
        );

    \I__14659\ : LocalMux
    port map (
            O => \N__62444\,
            I => \N__62434\
        );

    \I__14658\ : Span4Mux_h
    port map (
            O => \N__62441\,
            I => \N__62431\
        );

    \I__14657\ : InMux
    port map (
            O => \N__62440\,
            I => \N__62428\
        );

    \I__14656\ : LocalMux
    port map (
            O => \N__62437\,
            I => \c0.data_in_frame_8_0\
        );

    \I__14655\ : Odrv4
    port map (
            O => \N__62434\,
            I => \c0.data_in_frame_8_0\
        );

    \I__14654\ : Odrv4
    port map (
            O => \N__62431\,
            I => \c0.data_in_frame_8_0\
        );

    \I__14653\ : LocalMux
    port map (
            O => \N__62428\,
            I => \c0.data_in_frame_8_0\
        );

    \I__14652\ : InMux
    port map (
            O => \N__62419\,
            I => \N__62415\
        );

    \I__14651\ : InMux
    port map (
            O => \N__62418\,
            I => \N__62412\
        );

    \I__14650\ : LocalMux
    port map (
            O => \N__62415\,
            I => \N__62406\
        );

    \I__14649\ : LocalMux
    port map (
            O => \N__62412\,
            I => \N__62403\
        );

    \I__14648\ : InMux
    port map (
            O => \N__62411\,
            I => \N__62400\
        );

    \I__14647\ : CascadeMux
    port map (
            O => \N__62410\,
            I => \N__62396\
        );

    \I__14646\ : InMux
    port map (
            O => \N__62409\,
            I => \N__62393\
        );

    \I__14645\ : Span4Mux_v
    port map (
            O => \N__62406\,
            I => \N__62386\
        );

    \I__14644\ : Span4Mux_v
    port map (
            O => \N__62403\,
            I => \N__62386\
        );

    \I__14643\ : LocalMux
    port map (
            O => \N__62400\,
            I => \N__62386\
        );

    \I__14642\ : InMux
    port map (
            O => \N__62399\,
            I => \N__62383\
        );

    \I__14641\ : InMux
    port map (
            O => \N__62396\,
            I => \N__62379\
        );

    \I__14640\ : LocalMux
    port map (
            O => \N__62393\,
            I => \N__62374\
        );

    \I__14639\ : Span4Mux_h
    port map (
            O => \N__62386\,
            I => \N__62374\
        );

    \I__14638\ : LocalMux
    port map (
            O => \N__62383\,
            I => \N__62371\
        );

    \I__14637\ : InMux
    port map (
            O => \N__62382\,
            I => \N__62368\
        );

    \I__14636\ : LocalMux
    port map (
            O => \N__62379\,
            I => \c0.data_in_frame_7_7\
        );

    \I__14635\ : Odrv4
    port map (
            O => \N__62374\,
            I => \c0.data_in_frame_7_7\
        );

    \I__14634\ : Odrv4
    port map (
            O => \N__62371\,
            I => \c0.data_in_frame_7_7\
        );

    \I__14633\ : LocalMux
    port map (
            O => \N__62368\,
            I => \c0.data_in_frame_7_7\
        );

    \I__14632\ : CascadeMux
    port map (
            O => \N__62359\,
            I => \N__62356\
        );

    \I__14631\ : InMux
    port map (
            O => \N__62356\,
            I => \N__62350\
        );

    \I__14630\ : InMux
    port map (
            O => \N__62355\,
            I => \N__62347\
        );

    \I__14629\ : InMux
    port map (
            O => \N__62354\,
            I => \N__62344\
        );

    \I__14628\ : InMux
    port map (
            O => \N__62353\,
            I => \N__62340\
        );

    \I__14627\ : LocalMux
    port map (
            O => \N__62350\,
            I => \N__62335\
        );

    \I__14626\ : LocalMux
    port map (
            O => \N__62347\,
            I => \N__62335\
        );

    \I__14625\ : LocalMux
    port map (
            O => \N__62344\,
            I => \N__62332\
        );

    \I__14624\ : InMux
    port map (
            O => \N__62343\,
            I => \N__62329\
        );

    \I__14623\ : LocalMux
    port map (
            O => \N__62340\,
            I => \c0.data_in_frame_5_6\
        );

    \I__14622\ : Odrv4
    port map (
            O => \N__62335\,
            I => \c0.data_in_frame_5_6\
        );

    \I__14621\ : Odrv4
    port map (
            O => \N__62332\,
            I => \c0.data_in_frame_5_6\
        );

    \I__14620\ : LocalMux
    port map (
            O => \N__62329\,
            I => \c0.data_in_frame_5_6\
        );

    \I__14619\ : InMux
    port map (
            O => \N__62320\,
            I => \N__62317\
        );

    \I__14618\ : LocalMux
    port map (
            O => \N__62317\,
            I => \c0.n8_adj_3020\
        );

    \I__14617\ : CascadeMux
    port map (
            O => \N__62314\,
            I => \N__62310\
        );

    \I__14616\ : CascadeMux
    port map (
            O => \N__62313\,
            I => \N__62304\
        );

    \I__14615\ : InMux
    port map (
            O => \N__62310\,
            I => \N__62301\
        );

    \I__14614\ : CascadeMux
    port map (
            O => \N__62309\,
            I => \N__62298\
        );

    \I__14613\ : InMux
    port map (
            O => \N__62308\,
            I => \N__62293\
        );

    \I__14612\ : InMux
    port map (
            O => \N__62307\,
            I => \N__62293\
        );

    \I__14611\ : InMux
    port map (
            O => \N__62304\,
            I => \N__62290\
        );

    \I__14610\ : LocalMux
    port map (
            O => \N__62301\,
            I => \N__62287\
        );

    \I__14609\ : InMux
    port map (
            O => \N__62298\,
            I => \N__62284\
        );

    \I__14608\ : LocalMux
    port map (
            O => \N__62293\,
            I => \N__62281\
        );

    \I__14607\ : LocalMux
    port map (
            O => \N__62290\,
            I => \N__62278\
        );

    \I__14606\ : Span4Mux_v
    port map (
            O => \N__62287\,
            I => \N__62275\
        );

    \I__14605\ : LocalMux
    port map (
            O => \N__62284\,
            I => \N__62270\
        );

    \I__14604\ : Span4Mux_v
    port map (
            O => \N__62281\,
            I => \N__62270\
        );

    \I__14603\ : Span4Mux_h
    port map (
            O => \N__62278\,
            I => \N__62267\
        );

    \I__14602\ : Span4Mux_h
    port map (
            O => \N__62275\,
            I => \N__62264\
        );

    \I__14601\ : Odrv4
    port map (
            O => \N__62270\,
            I => \c0.data_in_frame_13_3\
        );

    \I__14600\ : Odrv4
    port map (
            O => \N__62267\,
            I => \c0.data_in_frame_13_3\
        );

    \I__14599\ : Odrv4
    port map (
            O => \N__62264\,
            I => \c0.data_in_frame_13_3\
        );

    \I__14598\ : InMux
    port map (
            O => \N__62257\,
            I => \N__62251\
        );

    \I__14597\ : InMux
    port map (
            O => \N__62256\,
            I => \N__62247\
        );

    \I__14596\ : InMux
    port map (
            O => \N__62255\,
            I => \N__62244\
        );

    \I__14595\ : CascadeMux
    port map (
            O => \N__62254\,
            I => \N__62241\
        );

    \I__14594\ : LocalMux
    port map (
            O => \N__62251\,
            I => \N__62238\
        );

    \I__14593\ : InMux
    port map (
            O => \N__62250\,
            I => \N__62235\
        );

    \I__14592\ : LocalMux
    port map (
            O => \N__62247\,
            I => \N__62232\
        );

    \I__14591\ : LocalMux
    port map (
            O => \N__62244\,
            I => \N__62229\
        );

    \I__14590\ : InMux
    port map (
            O => \N__62241\,
            I => \N__62226\
        );

    \I__14589\ : Span4Mux_v
    port map (
            O => \N__62238\,
            I => \N__62223\
        );

    \I__14588\ : LocalMux
    port map (
            O => \N__62235\,
            I => \N__62218\
        );

    \I__14587\ : Span4Mux_h
    port map (
            O => \N__62232\,
            I => \N__62218\
        );

    \I__14586\ : Span12Mux_v
    port map (
            O => \N__62229\,
            I => \N__62215\
        );

    \I__14585\ : LocalMux
    port map (
            O => \N__62226\,
            I => \c0.data_in_frame_9_2\
        );

    \I__14584\ : Odrv4
    port map (
            O => \N__62223\,
            I => \c0.data_in_frame_9_2\
        );

    \I__14583\ : Odrv4
    port map (
            O => \N__62218\,
            I => \c0.data_in_frame_9_2\
        );

    \I__14582\ : Odrv12
    port map (
            O => \N__62215\,
            I => \c0.data_in_frame_9_2\
        );

    \I__14581\ : InMux
    port map (
            O => \N__62206\,
            I => \N__62203\
        );

    \I__14580\ : LocalMux
    port map (
            O => \N__62203\,
            I => \N__62200\
        );

    \I__14579\ : Span4Mux_h
    port map (
            O => \N__62200\,
            I => \N__62194\
        );

    \I__14578\ : InMux
    port map (
            O => \N__62199\,
            I => \N__62187\
        );

    \I__14577\ : InMux
    port map (
            O => \N__62198\,
            I => \N__62187\
        );

    \I__14576\ : InMux
    port map (
            O => \N__62197\,
            I => \N__62187\
        );

    \I__14575\ : Odrv4
    port map (
            O => \N__62194\,
            I => \c0.n20095\
        );

    \I__14574\ : LocalMux
    port map (
            O => \N__62187\,
            I => \c0.n20095\
        );

    \I__14573\ : InMux
    port map (
            O => \N__62182\,
            I => \N__62177\
        );

    \I__14572\ : InMux
    port map (
            O => \N__62181\,
            I => \N__62173\
        );

    \I__14571\ : InMux
    port map (
            O => \N__62180\,
            I => \N__62169\
        );

    \I__14570\ : LocalMux
    port map (
            O => \N__62177\,
            I => \N__62166\
        );

    \I__14569\ : InMux
    port map (
            O => \N__62176\,
            I => \N__62160\
        );

    \I__14568\ : LocalMux
    port map (
            O => \N__62173\,
            I => \N__62157\
        );

    \I__14567\ : InMux
    port map (
            O => \N__62172\,
            I => \N__62153\
        );

    \I__14566\ : LocalMux
    port map (
            O => \N__62169\,
            I => \N__62148\
        );

    \I__14565\ : Span4Mux_v
    port map (
            O => \N__62166\,
            I => \N__62148\
        );

    \I__14564\ : InMux
    port map (
            O => \N__62165\,
            I => \N__62145\
        );

    \I__14563\ : InMux
    port map (
            O => \N__62164\,
            I => \N__62140\
        );

    \I__14562\ : InMux
    port map (
            O => \N__62163\,
            I => \N__62140\
        );

    \I__14561\ : LocalMux
    port map (
            O => \N__62160\,
            I => \N__62135\
        );

    \I__14560\ : Span4Mux_v
    port map (
            O => \N__62157\,
            I => \N__62135\
        );

    \I__14559\ : InMux
    port map (
            O => \N__62156\,
            I => \N__62132\
        );

    \I__14558\ : LocalMux
    port map (
            O => \N__62153\,
            I => \N__62123\
        );

    \I__14557\ : Span4Mux_h
    port map (
            O => \N__62148\,
            I => \N__62118\
        );

    \I__14556\ : LocalMux
    port map (
            O => \N__62145\,
            I => \N__62118\
        );

    \I__14555\ : LocalMux
    port map (
            O => \N__62140\,
            I => \N__62111\
        );

    \I__14554\ : Span4Mux_h
    port map (
            O => \N__62135\,
            I => \N__62111\
        );

    \I__14553\ : LocalMux
    port map (
            O => \N__62132\,
            I => \N__62111\
        );

    \I__14552\ : InMux
    port map (
            O => \N__62131\,
            I => \N__62108\
        );

    \I__14551\ : InMux
    port map (
            O => \N__62130\,
            I => \N__62105\
        );

    \I__14550\ : InMux
    port map (
            O => \N__62129\,
            I => \N__62100\
        );

    \I__14549\ : InMux
    port map (
            O => \N__62128\,
            I => \N__62100\
        );

    \I__14548\ : InMux
    port map (
            O => \N__62127\,
            I => \N__62095\
        );

    \I__14547\ : InMux
    port map (
            O => \N__62126\,
            I => \N__62095\
        );

    \I__14546\ : Odrv4
    port map (
            O => \N__62123\,
            I => data_in_frame_0_3
        );

    \I__14545\ : Odrv4
    port map (
            O => \N__62118\,
            I => data_in_frame_0_3
        );

    \I__14544\ : Odrv4
    port map (
            O => \N__62111\,
            I => data_in_frame_0_3
        );

    \I__14543\ : LocalMux
    port map (
            O => \N__62108\,
            I => data_in_frame_0_3
        );

    \I__14542\ : LocalMux
    port map (
            O => \N__62105\,
            I => data_in_frame_0_3
        );

    \I__14541\ : LocalMux
    port map (
            O => \N__62100\,
            I => data_in_frame_0_3
        );

    \I__14540\ : LocalMux
    port map (
            O => \N__62095\,
            I => data_in_frame_0_3
        );

    \I__14539\ : CascadeMux
    port map (
            O => \N__62080\,
            I => \N__62077\
        );

    \I__14538\ : InMux
    port map (
            O => \N__62077\,
            I => \N__62073\
        );

    \I__14537\ : InMux
    port map (
            O => \N__62076\,
            I => \N__62070\
        );

    \I__14536\ : LocalMux
    port map (
            O => \N__62073\,
            I => \N__62067\
        );

    \I__14535\ : LocalMux
    port map (
            O => \N__62070\,
            I => \c0.n5240\
        );

    \I__14534\ : Odrv12
    port map (
            O => \N__62067\,
            I => \c0.n5240\
        );

    \I__14533\ : CascadeMux
    port map (
            O => \N__62062\,
            I => \c0.n7_cascade_\
        );

    \I__14532\ : InMux
    port map (
            O => \N__62059\,
            I => \N__62053\
        );

    \I__14531\ : InMux
    port map (
            O => \N__62058\,
            I => \N__62053\
        );

    \I__14530\ : LocalMux
    port map (
            O => \N__62053\,
            I => \N__62050\
        );

    \I__14529\ : Span4Mux_v
    port map (
            O => \N__62050\,
            I => \N__62045\
        );

    \I__14528\ : CascadeMux
    port map (
            O => \N__62049\,
            I => \N__62042\
        );

    \I__14527\ : CascadeMux
    port map (
            O => \N__62048\,
            I => \N__62036\
        );

    \I__14526\ : Span4Mux_h
    port map (
            O => \N__62045\,
            I => \N__62031\
        );

    \I__14525\ : InMux
    port map (
            O => \N__62042\,
            I => \N__62027\
        );

    \I__14524\ : InMux
    port map (
            O => \N__62041\,
            I => \N__62024\
        );

    \I__14523\ : InMux
    port map (
            O => \N__62040\,
            I => \N__62019\
        );

    \I__14522\ : InMux
    port map (
            O => \N__62039\,
            I => \N__62019\
        );

    \I__14521\ : InMux
    port map (
            O => \N__62036\,
            I => \N__62013\
        );

    \I__14520\ : InMux
    port map (
            O => \N__62035\,
            I => \N__62013\
        );

    \I__14519\ : InMux
    port map (
            O => \N__62034\,
            I => \N__62010\
        );

    \I__14518\ : Span4Mux_v
    port map (
            O => \N__62031\,
            I => \N__62006\
        );

    \I__14517\ : InMux
    port map (
            O => \N__62030\,
            I => \N__62003\
        );

    \I__14516\ : LocalMux
    port map (
            O => \N__62027\,
            I => \N__61997\
        );

    \I__14515\ : LocalMux
    port map (
            O => \N__62024\,
            I => \N__61997\
        );

    \I__14514\ : LocalMux
    port map (
            O => \N__62019\,
            I => \N__61994\
        );

    \I__14513\ : InMux
    port map (
            O => \N__62018\,
            I => \N__61991\
        );

    \I__14512\ : LocalMux
    port map (
            O => \N__62013\,
            I => \N__61988\
        );

    \I__14511\ : LocalMux
    port map (
            O => \N__62010\,
            I => \N__61984\
        );

    \I__14510\ : InMux
    port map (
            O => \N__62009\,
            I => \N__61981\
        );

    \I__14509\ : Span4Mux_h
    port map (
            O => \N__62006\,
            I => \N__61976\
        );

    \I__14508\ : LocalMux
    port map (
            O => \N__62003\,
            I => \N__61976\
        );

    \I__14507\ : CascadeMux
    port map (
            O => \N__62002\,
            I => \N__61973\
        );

    \I__14506\ : Span4Mux_v
    port map (
            O => \N__61997\,
            I => \N__61968\
        );

    \I__14505\ : Span4Mux_v
    port map (
            O => \N__61994\,
            I => \N__61968\
        );

    \I__14504\ : LocalMux
    port map (
            O => \N__61991\,
            I => \N__61965\
        );

    \I__14503\ : Span4Mux_v
    port map (
            O => \N__61988\,
            I => \N__61962\
        );

    \I__14502\ : CascadeMux
    port map (
            O => \N__61987\,
            I => \N__61959\
        );

    \I__14501\ : Span4Mux_v
    port map (
            O => \N__61984\,
            I => \N__61956\
        );

    \I__14500\ : LocalMux
    port map (
            O => \N__61981\,
            I => \N__61951\
        );

    \I__14499\ : Span4Mux_v
    port map (
            O => \N__61976\,
            I => \N__61948\
        );

    \I__14498\ : InMux
    port map (
            O => \N__61973\,
            I => \N__61945\
        );

    \I__14497\ : Span4Mux_h
    port map (
            O => \N__61968\,
            I => \N__61942\
        );

    \I__14496\ : Span4Mux_v
    port map (
            O => \N__61965\,
            I => \N__61937\
        );

    \I__14495\ : Span4Mux_h
    port map (
            O => \N__61962\,
            I => \N__61937\
        );

    \I__14494\ : InMux
    port map (
            O => \N__61959\,
            I => \N__61934\
        );

    \I__14493\ : Sp12to4
    port map (
            O => \N__61956\,
            I => \N__61931\
        );

    \I__14492\ : InMux
    port map (
            O => \N__61955\,
            I => \N__61928\
        );

    \I__14491\ : InMux
    port map (
            O => \N__61954\,
            I => \N__61924\
        );

    \I__14490\ : Span4Mux_v
    port map (
            O => \N__61951\,
            I => \N__61921\
        );

    \I__14489\ : Span4Mux_h
    port map (
            O => \N__61948\,
            I => \N__61916\
        );

    \I__14488\ : LocalMux
    port map (
            O => \N__61945\,
            I => \N__61916\
        );

    \I__14487\ : Span4Mux_h
    port map (
            O => \N__61942\,
            I => \N__61911\
        );

    \I__14486\ : Span4Mux_v
    port map (
            O => \N__61937\,
            I => \N__61911\
        );

    \I__14485\ : LocalMux
    port map (
            O => \N__61934\,
            I => \N__61904\
        );

    \I__14484\ : Span12Mux_h
    port map (
            O => \N__61931\,
            I => \N__61904\
        );

    \I__14483\ : LocalMux
    port map (
            O => \N__61928\,
            I => \N__61904\
        );

    \I__14482\ : InMux
    port map (
            O => \N__61927\,
            I => \N__61901\
        );

    \I__14481\ : LocalMux
    port map (
            O => \N__61924\,
            I => \N__61898\
        );

    \I__14480\ : Span4Mux_h
    port map (
            O => \N__61921\,
            I => \N__61893\
        );

    \I__14479\ : Span4Mux_h
    port map (
            O => \N__61916\,
            I => \N__61893\
        );

    \I__14478\ : Sp12to4
    port map (
            O => \N__61911\,
            I => \N__61888\
        );

    \I__14477\ : Span12Mux_v
    port map (
            O => \N__61904\,
            I => \N__61888\
        );

    \I__14476\ : LocalMux
    port map (
            O => \N__61901\,
            I => \c0.n9_adj_3038\
        );

    \I__14475\ : Odrv4
    port map (
            O => \N__61898\,
            I => \c0.n9_adj_3038\
        );

    \I__14474\ : Odrv4
    port map (
            O => \N__61893\,
            I => \c0.n9_adj_3038\
        );

    \I__14473\ : Odrv12
    port map (
            O => \N__61888\,
            I => \c0.n9_adj_3038\
        );

    \I__14472\ : InMux
    port map (
            O => \N__61879\,
            I => \N__61875\
        );

    \I__14471\ : InMux
    port map (
            O => \N__61878\,
            I => \N__61868\
        );

    \I__14470\ : LocalMux
    port map (
            O => \N__61875\,
            I => \N__61865\
        );

    \I__14469\ : InMux
    port map (
            O => \N__61874\,
            I => \N__61862\
        );

    \I__14468\ : InMux
    port map (
            O => \N__61873\,
            I => \N__61857\
        );

    \I__14467\ : InMux
    port map (
            O => \N__61872\,
            I => \N__61852\
        );

    \I__14466\ : InMux
    port map (
            O => \N__61871\,
            I => \N__61852\
        );

    \I__14465\ : LocalMux
    port map (
            O => \N__61868\,
            I => \N__61847\
        );

    \I__14464\ : Span4Mux_h
    port map (
            O => \N__61865\,
            I => \N__61847\
        );

    \I__14463\ : LocalMux
    port map (
            O => \N__61862\,
            I => \N__61844\
        );

    \I__14462\ : CascadeMux
    port map (
            O => \N__61861\,
            I => \N__61841\
        );

    \I__14461\ : InMux
    port map (
            O => \N__61860\,
            I => \N__61838\
        );

    \I__14460\ : LocalMux
    port map (
            O => \N__61857\,
            I => \N__61833\
        );

    \I__14459\ : LocalMux
    port map (
            O => \N__61852\,
            I => \N__61833\
        );

    \I__14458\ : Span4Mux_v
    port map (
            O => \N__61847\,
            I => \N__61830\
        );

    \I__14457\ : Span4Mux_h
    port map (
            O => \N__61844\,
            I => \N__61827\
        );

    \I__14456\ : InMux
    port map (
            O => \N__61841\,
            I => \N__61823\
        );

    \I__14455\ : LocalMux
    port map (
            O => \N__61838\,
            I => \N__61820\
        );

    \I__14454\ : Span4Mux_v
    port map (
            O => \N__61833\,
            I => \N__61813\
        );

    \I__14453\ : Span4Mux_h
    port map (
            O => \N__61830\,
            I => \N__61813\
        );

    \I__14452\ : Span4Mux_h
    port map (
            O => \N__61827\,
            I => \N__61813\
        );

    \I__14451\ : InMux
    port map (
            O => \N__61826\,
            I => \N__61810\
        );

    \I__14450\ : LocalMux
    port map (
            O => \N__61823\,
            I => \c0.data_in_frame_6_7\
        );

    \I__14449\ : Odrv12
    port map (
            O => \N__61820\,
            I => \c0.data_in_frame_6_7\
        );

    \I__14448\ : Odrv4
    port map (
            O => \N__61813\,
            I => \c0.data_in_frame_6_7\
        );

    \I__14447\ : LocalMux
    port map (
            O => \N__61810\,
            I => \c0.data_in_frame_6_7\
        );

    \I__14446\ : InMux
    port map (
            O => \N__61801\,
            I => \N__61798\
        );

    \I__14445\ : LocalMux
    port map (
            O => \N__61798\,
            I => \N__61791\
        );

    \I__14444\ : InMux
    port map (
            O => \N__61797\,
            I => \N__61786\
        );

    \I__14443\ : InMux
    port map (
            O => \N__61796\,
            I => \N__61786\
        );

    \I__14442\ : InMux
    port map (
            O => \N__61795\,
            I => \N__61781\
        );

    \I__14441\ : InMux
    port map (
            O => \N__61794\,
            I => \N__61781\
        );

    \I__14440\ : Span4Mux_v
    port map (
            O => \N__61791\,
            I => \N__61774\
        );

    \I__14439\ : LocalMux
    port map (
            O => \N__61786\,
            I => \N__61769\
        );

    \I__14438\ : LocalMux
    port map (
            O => \N__61781\,
            I => \N__61769\
        );

    \I__14437\ : InMux
    port map (
            O => \N__61780\,
            I => \N__61761\
        );

    \I__14436\ : InMux
    port map (
            O => \N__61779\,
            I => \N__61761\
        );

    \I__14435\ : CascadeMux
    port map (
            O => \N__61778\,
            I => \N__61749\
        );

    \I__14434\ : CascadeMux
    port map (
            O => \N__61777\,
            I => \N__61746\
        );

    \I__14433\ : Span4Mux_h
    port map (
            O => \N__61774\,
            I => \N__61739\
        );

    \I__14432\ : Span4Mux_v
    port map (
            O => \N__61769\,
            I => \N__61739\
        );

    \I__14431\ : InMux
    port map (
            O => \N__61768\,
            I => \N__61732\
        );

    \I__14430\ : InMux
    port map (
            O => \N__61767\,
            I => \N__61732\
        );

    \I__14429\ : InMux
    port map (
            O => \N__61766\,
            I => \N__61732\
        );

    \I__14428\ : LocalMux
    port map (
            O => \N__61761\,
            I => \N__61727\
        );

    \I__14427\ : InMux
    port map (
            O => \N__61760\,
            I => \N__61716\
        );

    \I__14426\ : InMux
    port map (
            O => \N__61759\,
            I => \N__61716\
        );

    \I__14425\ : InMux
    port map (
            O => \N__61758\,
            I => \N__61716\
        );

    \I__14424\ : InMux
    port map (
            O => \N__61757\,
            I => \N__61713\
        );

    \I__14423\ : InMux
    port map (
            O => \N__61756\,
            I => \N__61702\
        );

    \I__14422\ : InMux
    port map (
            O => \N__61755\,
            I => \N__61702\
        );

    \I__14421\ : InMux
    port map (
            O => \N__61754\,
            I => \N__61702\
        );

    \I__14420\ : InMux
    port map (
            O => \N__61753\,
            I => \N__61702\
        );

    \I__14419\ : InMux
    port map (
            O => \N__61752\,
            I => \N__61702\
        );

    \I__14418\ : InMux
    port map (
            O => \N__61749\,
            I => \N__61693\
        );

    \I__14417\ : InMux
    port map (
            O => \N__61746\,
            I => \N__61693\
        );

    \I__14416\ : InMux
    port map (
            O => \N__61745\,
            I => \N__61693\
        );

    \I__14415\ : InMux
    port map (
            O => \N__61744\,
            I => \N__61693\
        );

    \I__14414\ : Span4Mux_h
    port map (
            O => \N__61739\,
            I => \N__61678\
        );

    \I__14413\ : LocalMux
    port map (
            O => \N__61732\,
            I => \N__61678\
        );

    \I__14412\ : InMux
    port map (
            O => \N__61731\,
            I => \N__61674\
        );

    \I__14411\ : InMux
    port map (
            O => \N__61730\,
            I => \N__61667\
        );

    \I__14410\ : Span4Mux_v
    port map (
            O => \N__61727\,
            I => \N__61664\
        );

    \I__14409\ : InMux
    port map (
            O => \N__61726\,
            I => \N__61659\
        );

    \I__14408\ : InMux
    port map (
            O => \N__61725\,
            I => \N__61659\
        );

    \I__14407\ : InMux
    port map (
            O => \N__61724\,
            I => \N__61654\
        );

    \I__14406\ : InMux
    port map (
            O => \N__61723\,
            I => \N__61654\
        );

    \I__14405\ : LocalMux
    port map (
            O => \N__61716\,
            I => \N__61651\
        );

    \I__14404\ : LocalMux
    port map (
            O => \N__61713\,
            I => \N__61644\
        );

    \I__14403\ : LocalMux
    port map (
            O => \N__61702\,
            I => \N__61644\
        );

    \I__14402\ : LocalMux
    port map (
            O => \N__61693\,
            I => \N__61644\
        );

    \I__14401\ : InMux
    port map (
            O => \N__61692\,
            I => \N__61635\
        );

    \I__14400\ : InMux
    port map (
            O => \N__61691\,
            I => \N__61635\
        );

    \I__14399\ : InMux
    port map (
            O => \N__61690\,
            I => \N__61635\
        );

    \I__14398\ : InMux
    port map (
            O => \N__61689\,
            I => \N__61635\
        );

    \I__14397\ : InMux
    port map (
            O => \N__61688\,
            I => \N__61632\
        );

    \I__14396\ : InMux
    port map (
            O => \N__61687\,
            I => \N__61627\
        );

    \I__14395\ : InMux
    port map (
            O => \N__61686\,
            I => \N__61627\
        );

    \I__14394\ : InMux
    port map (
            O => \N__61685\,
            I => \N__61624\
        );

    \I__14393\ : InMux
    port map (
            O => \N__61684\,
            I => \N__61619\
        );

    \I__14392\ : InMux
    port map (
            O => \N__61683\,
            I => \N__61619\
        );

    \I__14391\ : Span4Mux_h
    port map (
            O => \N__61678\,
            I => \N__61616\
        );

    \I__14390\ : InMux
    port map (
            O => \N__61677\,
            I => \N__61612\
        );

    \I__14389\ : LocalMux
    port map (
            O => \N__61674\,
            I => \N__61609\
        );

    \I__14388\ : InMux
    port map (
            O => \N__61673\,
            I => \N__61600\
        );

    \I__14387\ : InMux
    port map (
            O => \N__61672\,
            I => \N__61600\
        );

    \I__14386\ : InMux
    port map (
            O => \N__61671\,
            I => \N__61600\
        );

    \I__14385\ : InMux
    port map (
            O => \N__61670\,
            I => \N__61600\
        );

    \I__14384\ : LocalMux
    port map (
            O => \N__61667\,
            I => \N__61584\
        );

    \I__14383\ : Span4Mux_h
    port map (
            O => \N__61664\,
            I => \N__61584\
        );

    \I__14382\ : LocalMux
    port map (
            O => \N__61659\,
            I => \N__61584\
        );

    \I__14381\ : LocalMux
    port map (
            O => \N__61654\,
            I => \N__61584\
        );

    \I__14380\ : Span4Mux_v
    port map (
            O => \N__61651\,
            I => \N__61577\
        );

    \I__14379\ : Span4Mux_v
    port map (
            O => \N__61644\,
            I => \N__61577\
        );

    \I__14378\ : LocalMux
    port map (
            O => \N__61635\,
            I => \N__61577\
        );

    \I__14377\ : LocalMux
    port map (
            O => \N__61632\,
            I => \N__61572\
        );

    \I__14376\ : LocalMux
    port map (
            O => \N__61627\,
            I => \N__61572\
        );

    \I__14375\ : LocalMux
    port map (
            O => \N__61624\,
            I => \N__61567\
        );

    \I__14374\ : LocalMux
    port map (
            O => \N__61619\,
            I => \N__61567\
        );

    \I__14373\ : Span4Mux_v
    port map (
            O => \N__61616\,
            I => \N__61564\
        );

    \I__14372\ : InMux
    port map (
            O => \N__61615\,
            I => \N__61561\
        );

    \I__14371\ : LocalMux
    port map (
            O => \N__61612\,
            I => \N__61553\
        );

    \I__14370\ : Span4Mux_v
    port map (
            O => \N__61609\,
            I => \N__61553\
        );

    \I__14369\ : LocalMux
    port map (
            O => \N__61600\,
            I => \N__61553\
        );

    \I__14368\ : CascadeMux
    port map (
            O => \N__61599\,
            I => \N__61546\
        );

    \I__14367\ : InMux
    port map (
            O => \N__61598\,
            I => \N__61543\
        );

    \I__14366\ : InMux
    port map (
            O => \N__61597\,
            I => \N__61538\
        );

    \I__14365\ : InMux
    port map (
            O => \N__61596\,
            I => \N__61538\
        );

    \I__14364\ : InMux
    port map (
            O => \N__61595\,
            I => \N__61531\
        );

    \I__14363\ : InMux
    port map (
            O => \N__61594\,
            I => \N__61531\
        );

    \I__14362\ : InMux
    port map (
            O => \N__61593\,
            I => \N__61531\
        );

    \I__14361\ : Span4Mux_v
    port map (
            O => \N__61584\,
            I => \N__61522\
        );

    \I__14360\ : Span4Mux_h
    port map (
            O => \N__61577\,
            I => \N__61522\
        );

    \I__14359\ : Span4Mux_v
    port map (
            O => \N__61572\,
            I => \N__61522\
        );

    \I__14358\ : Span4Mux_v
    port map (
            O => \N__61567\,
            I => \N__61522\
        );

    \I__14357\ : Sp12to4
    port map (
            O => \N__61564\,
            I => \N__61519\
        );

    \I__14356\ : LocalMux
    port map (
            O => \N__61561\,
            I => \N__61516\
        );

    \I__14355\ : InMux
    port map (
            O => \N__61560\,
            I => \N__61513\
        );

    \I__14354\ : Span4Mux_h
    port map (
            O => \N__61553\,
            I => \N__61510\
        );

    \I__14353\ : InMux
    port map (
            O => \N__61552\,
            I => \N__61501\
        );

    \I__14352\ : InMux
    port map (
            O => \N__61551\,
            I => \N__61501\
        );

    \I__14351\ : InMux
    port map (
            O => \N__61550\,
            I => \N__61501\
        );

    \I__14350\ : InMux
    port map (
            O => \N__61549\,
            I => \N__61501\
        );

    \I__14349\ : InMux
    port map (
            O => \N__61546\,
            I => \N__61498\
        );

    \I__14348\ : LocalMux
    port map (
            O => \N__61543\,
            I => \N__61485\
        );

    \I__14347\ : LocalMux
    port map (
            O => \N__61538\,
            I => \N__61485\
        );

    \I__14346\ : LocalMux
    port map (
            O => \N__61531\,
            I => \N__61485\
        );

    \I__14345\ : Sp12to4
    port map (
            O => \N__61522\,
            I => \N__61485\
        );

    \I__14344\ : Span12Mux_s7_h
    port map (
            O => \N__61519\,
            I => \N__61485\
        );

    \I__14343\ : Sp12to4
    port map (
            O => \N__61516\,
            I => \N__61485\
        );

    \I__14342\ : LocalMux
    port map (
            O => \N__61513\,
            I => \N__61478\
        );

    \I__14341\ : Span4Mux_h
    port map (
            O => \N__61510\,
            I => \N__61478\
        );

    \I__14340\ : LocalMux
    port map (
            O => \N__61501\,
            I => \N__61478\
        );

    \I__14339\ : LocalMux
    port map (
            O => \N__61498\,
            I => \N__61475\
        );

    \I__14338\ : Span12Mux_h
    port map (
            O => \N__61485\,
            I => \N__61472\
        );

    \I__14337\ : Sp12to4
    port map (
            O => \N__61478\,
            I => \N__61469\
        );

    \I__14336\ : Span12Mux_h
    port map (
            O => \N__61475\,
            I => \N__61466\
        );

    \I__14335\ : Span12Mux_v
    port map (
            O => \N__61472\,
            I => \N__61461\
        );

    \I__14334\ : Span12Mux_v
    port map (
            O => \N__61469\,
            I => \N__61461\
        );

    \I__14333\ : Odrv12
    port map (
            O => \N__61466\,
            I => \c0.n19098\
        );

    \I__14332\ : Odrv12
    port map (
            O => \N__61461\,
            I => \c0.n19098\
        );

    \I__14331\ : InMux
    port map (
            O => \N__61456\,
            I => \N__61450\
        );

    \I__14330\ : InMux
    port map (
            O => \N__61455\,
            I => \N__61443\
        );

    \I__14329\ : InMux
    port map (
            O => \N__61454\,
            I => \N__61443\
        );

    \I__14328\ : InMux
    port map (
            O => \N__61453\,
            I => \N__61440\
        );

    \I__14327\ : LocalMux
    port map (
            O => \N__61450\,
            I => \N__61437\
        );

    \I__14326\ : CascadeMux
    port map (
            O => \N__61449\,
            I => \N__61434\
        );

    \I__14325\ : InMux
    port map (
            O => \N__61448\,
            I => \N__61431\
        );

    \I__14324\ : LocalMux
    port map (
            O => \N__61443\,
            I => \N__61425\
        );

    \I__14323\ : LocalMux
    port map (
            O => \N__61440\,
            I => \N__61425\
        );

    \I__14322\ : Span4Mux_h
    port map (
            O => \N__61437\,
            I => \N__61421\
        );

    \I__14321\ : InMux
    port map (
            O => \N__61434\,
            I => \N__61418\
        );

    \I__14320\ : LocalMux
    port map (
            O => \N__61431\,
            I => \N__61415\
        );

    \I__14319\ : InMux
    port map (
            O => \N__61430\,
            I => \N__61412\
        );

    \I__14318\ : Span4Mux_v
    port map (
            O => \N__61425\,
            I => \N__61409\
        );

    \I__14317\ : CascadeMux
    port map (
            O => \N__61424\,
            I => \N__61404\
        );

    \I__14316\ : Span4Mux_v
    port map (
            O => \N__61421\,
            I => \N__61401\
        );

    \I__14315\ : LocalMux
    port map (
            O => \N__61418\,
            I => \N__61398\
        );

    \I__14314\ : Span4Mux_v
    port map (
            O => \N__61415\,
            I => \N__61395\
        );

    \I__14313\ : LocalMux
    port map (
            O => \N__61412\,
            I => \N__61392\
        );

    \I__14312\ : Span4Mux_v
    port map (
            O => \N__61409\,
            I => \N__61389\
        );

    \I__14311\ : InMux
    port map (
            O => \N__61408\,
            I => \N__61384\
        );

    \I__14310\ : InMux
    port map (
            O => \N__61407\,
            I => \N__61384\
        );

    \I__14309\ : InMux
    port map (
            O => \N__61404\,
            I => \N__61381\
        );

    \I__14308\ : Sp12to4
    port map (
            O => \N__61401\,
            I => \N__61378\
        );

    \I__14307\ : Span4Mux_v
    port map (
            O => \N__61398\,
            I => \N__61373\
        );

    \I__14306\ : Span4Mux_v
    port map (
            O => \N__61395\,
            I => \N__61373\
        );

    \I__14305\ : Span4Mux_v
    port map (
            O => \N__61392\,
            I => \N__61368\
        );

    \I__14304\ : Span4Mux_h
    port map (
            O => \N__61389\,
            I => \N__61368\
        );

    \I__14303\ : LocalMux
    port map (
            O => \N__61384\,
            I => \N__61361\
        );

    \I__14302\ : LocalMux
    port map (
            O => \N__61381\,
            I => \N__61361\
        );

    \I__14301\ : Span12Mux_v
    port map (
            O => \N__61378\,
            I => \N__61361\
        );

    \I__14300\ : Sp12to4
    port map (
            O => \N__61373\,
            I => \N__61354\
        );

    \I__14299\ : Sp12to4
    port map (
            O => \N__61368\,
            I => \N__61354\
        );

    \I__14298\ : Span12Mux_v
    port map (
            O => \N__61361\,
            I => \N__61354\
        );

    \I__14297\ : Odrv12
    port map (
            O => \N__61354\,
            I => \c0.n9_adj_3251\
        );

    \I__14296\ : InMux
    port map (
            O => \N__61351\,
            I => \N__61348\
        );

    \I__14295\ : LocalMux
    port map (
            O => \N__61348\,
            I => \N__61342\
        );

    \I__14294\ : InMux
    port map (
            O => \N__61347\,
            I => \N__61337\
        );

    \I__14293\ : InMux
    port map (
            O => \N__61346\,
            I => \N__61337\
        );

    \I__14292\ : CascadeMux
    port map (
            O => \N__61345\,
            I => \N__61334\
        );

    \I__14291\ : Span4Mux_h
    port map (
            O => \N__61342\,
            I => \N__61331\
        );

    \I__14290\ : LocalMux
    port map (
            O => \N__61337\,
            I => \N__61328\
        );

    \I__14289\ : InMux
    port map (
            O => \N__61334\,
            I => \N__61323\
        );

    \I__14288\ : Span4Mux_h
    port map (
            O => \N__61331\,
            I => \N__61318\
        );

    \I__14287\ : Span4Mux_v
    port map (
            O => \N__61328\,
            I => \N__61318\
        );

    \I__14286\ : InMux
    port map (
            O => \N__61327\,
            I => \N__61313\
        );

    \I__14285\ : InMux
    port map (
            O => \N__61326\,
            I => \N__61313\
        );

    \I__14284\ : LocalMux
    port map (
            O => \N__61323\,
            I => \c0.data_in_frame_3_4\
        );

    \I__14283\ : Odrv4
    port map (
            O => \N__61318\,
            I => \c0.data_in_frame_3_4\
        );

    \I__14282\ : LocalMux
    port map (
            O => \N__61313\,
            I => \c0.data_in_frame_3_4\
        );

    \I__14281\ : InMux
    port map (
            O => \N__61306\,
            I => \N__61303\
        );

    \I__14280\ : LocalMux
    port map (
            O => \N__61303\,
            I => \c0.n12_adj_2998\
        );

    \I__14279\ : InMux
    port map (
            O => \N__61300\,
            I => \N__61297\
        );

    \I__14278\ : LocalMux
    port map (
            O => \N__61297\,
            I => \N__61294\
        );

    \I__14277\ : Span4Mux_h
    port map (
            O => \N__61294\,
            I => \N__61291\
        );

    \I__14276\ : Span4Mux_h
    port map (
            O => \N__61291\,
            I => \N__61288\
        );

    \I__14275\ : Odrv4
    port map (
            O => \N__61288\,
            I => \c0.n19176\
        );

    \I__14274\ : InMux
    port map (
            O => \N__61285\,
            I => \N__61281\
        );

    \I__14273\ : InMux
    port map (
            O => \N__61284\,
            I => \N__61278\
        );

    \I__14272\ : LocalMux
    port map (
            O => \N__61281\,
            I => \N__61275\
        );

    \I__14271\ : LocalMux
    port map (
            O => \N__61278\,
            I => \N__61272\
        );

    \I__14270\ : Span4Mux_h
    port map (
            O => \N__61275\,
            I => \N__61269\
        );

    \I__14269\ : Span12Mux_v
    port map (
            O => \N__61272\,
            I => \N__61266\
        );

    \I__14268\ : Odrv4
    port map (
            O => \N__61269\,
            I => \c0.n11953\
        );

    \I__14267\ : Odrv12
    port map (
            O => \N__61266\,
            I => \c0.n11953\
        );

    \I__14266\ : InMux
    port map (
            O => \N__61261\,
            I => \N__61258\
        );

    \I__14265\ : LocalMux
    port map (
            O => \N__61258\,
            I => \N__61255\
        );

    \I__14264\ : Span4Mux_v
    port map (
            O => \N__61255\,
            I => \N__61251\
        );

    \I__14263\ : InMux
    port map (
            O => \N__61254\,
            I => \N__61248\
        );

    \I__14262\ : Sp12to4
    port map (
            O => \N__61251\,
            I => \N__61241\
        );

    \I__14261\ : LocalMux
    port map (
            O => \N__61248\,
            I => \N__61241\
        );

    \I__14260\ : InMux
    port map (
            O => \N__61247\,
            I => \N__61236\
        );

    \I__14259\ : InMux
    port map (
            O => \N__61246\,
            I => \N__61236\
        );

    \I__14258\ : Odrv12
    port map (
            O => \N__61241\,
            I => \c0.data_in_frame_5_2\
        );

    \I__14257\ : LocalMux
    port map (
            O => \N__61236\,
            I => \c0.data_in_frame_5_2\
        );

    \I__14256\ : InMux
    port map (
            O => \N__61231\,
            I => \N__61228\
        );

    \I__14255\ : LocalMux
    port map (
            O => \N__61228\,
            I => \N__61222\
        );

    \I__14254\ : InMux
    port map (
            O => \N__61227\,
            I => \N__61219\
        );

    \I__14253\ : InMux
    port map (
            O => \N__61226\,
            I => \N__61216\
        );

    \I__14252\ : InMux
    port map (
            O => \N__61225\,
            I => \N__61213\
        );

    \I__14251\ : Span4Mux_v
    port map (
            O => \N__61222\,
            I => \N__61209\
        );

    \I__14250\ : LocalMux
    port map (
            O => \N__61219\,
            I => \N__61206\
        );

    \I__14249\ : LocalMux
    port map (
            O => \N__61216\,
            I => \N__61202\
        );

    \I__14248\ : LocalMux
    port map (
            O => \N__61213\,
            I => \N__61199\
        );

    \I__14247\ : InMux
    port map (
            O => \N__61212\,
            I => \N__61190\
        );

    \I__14246\ : Span4Mux_h
    port map (
            O => \N__61209\,
            I => \N__61187\
        );

    \I__14245\ : Span4Mux_h
    port map (
            O => \N__61206\,
            I => \N__61184\
        );

    \I__14244\ : InMux
    port map (
            O => \N__61205\,
            I => \N__61181\
        );

    \I__14243\ : Span4Mux_h
    port map (
            O => \N__61202\,
            I => \N__61176\
        );

    \I__14242\ : Span4Mux_h
    port map (
            O => \N__61199\,
            I => \N__61176\
        );

    \I__14241\ : InMux
    port map (
            O => \N__61198\,
            I => \N__61173\
        );

    \I__14240\ : InMux
    port map (
            O => \N__61197\,
            I => \N__61170\
        );

    \I__14239\ : InMux
    port map (
            O => \N__61196\,
            I => \N__61163\
        );

    \I__14238\ : InMux
    port map (
            O => \N__61195\,
            I => \N__61163\
        );

    \I__14237\ : InMux
    port map (
            O => \N__61194\,
            I => \N__61163\
        );

    \I__14236\ : InMux
    port map (
            O => \N__61193\,
            I => \N__61160\
        );

    \I__14235\ : LocalMux
    port map (
            O => \N__61190\,
            I => data_in_frame_1_3
        );

    \I__14234\ : Odrv4
    port map (
            O => \N__61187\,
            I => data_in_frame_1_3
        );

    \I__14233\ : Odrv4
    port map (
            O => \N__61184\,
            I => data_in_frame_1_3
        );

    \I__14232\ : LocalMux
    port map (
            O => \N__61181\,
            I => data_in_frame_1_3
        );

    \I__14231\ : Odrv4
    port map (
            O => \N__61176\,
            I => data_in_frame_1_3
        );

    \I__14230\ : LocalMux
    port map (
            O => \N__61173\,
            I => data_in_frame_1_3
        );

    \I__14229\ : LocalMux
    port map (
            O => \N__61170\,
            I => data_in_frame_1_3
        );

    \I__14228\ : LocalMux
    port map (
            O => \N__61163\,
            I => data_in_frame_1_3
        );

    \I__14227\ : LocalMux
    port map (
            O => \N__61160\,
            I => data_in_frame_1_3
        );

    \I__14226\ : CascadeMux
    port map (
            O => \N__61141\,
            I => \N__61138\
        );

    \I__14225\ : InMux
    port map (
            O => \N__61138\,
            I => \N__61135\
        );

    \I__14224\ : LocalMux
    port map (
            O => \N__61135\,
            I => \c0.n55_adj_3500\
        );

    \I__14223\ : CascadeMux
    port map (
            O => \N__61132\,
            I => \N__61128\
        );

    \I__14222\ : InMux
    port map (
            O => \N__61131\,
            I => \N__61123\
        );

    \I__14221\ : InMux
    port map (
            O => \N__61128\,
            I => \N__61119\
        );

    \I__14220\ : InMux
    port map (
            O => \N__61127\,
            I => \N__61112\
        );

    \I__14219\ : InMux
    port map (
            O => \N__61126\,
            I => \N__61112\
        );

    \I__14218\ : LocalMux
    port map (
            O => \N__61123\,
            I => \N__61109\
        );

    \I__14217\ : InMux
    port map (
            O => \N__61122\,
            I => \N__61106\
        );

    \I__14216\ : LocalMux
    port map (
            O => \N__61119\,
            I => \N__61103\
        );

    \I__14215\ : InMux
    port map (
            O => \N__61118\,
            I => \N__61100\
        );

    \I__14214\ : InMux
    port map (
            O => \N__61117\,
            I => \N__61096\
        );

    \I__14213\ : LocalMux
    port map (
            O => \N__61112\,
            I => \N__61093\
        );

    \I__14212\ : Span4Mux_h
    port map (
            O => \N__61109\,
            I => \N__61087\
        );

    \I__14211\ : LocalMux
    port map (
            O => \N__61106\,
            I => \N__61087\
        );

    \I__14210\ : Span4Mux_h
    port map (
            O => \N__61103\,
            I => \N__61082\
        );

    \I__14209\ : LocalMux
    port map (
            O => \N__61100\,
            I => \N__61082\
        );

    \I__14208\ : CascadeMux
    port map (
            O => \N__61099\,
            I => \N__61074\
        );

    \I__14207\ : LocalMux
    port map (
            O => \N__61096\,
            I => \N__61070\
        );

    \I__14206\ : Span4Mux_v
    port map (
            O => \N__61093\,
            I => \N__61067\
        );

    \I__14205\ : InMux
    port map (
            O => \N__61092\,
            I => \N__61064\
        );

    \I__14204\ : Span4Mux_v
    port map (
            O => \N__61087\,
            I => \N__61061\
        );

    \I__14203\ : Span4Mux_h
    port map (
            O => \N__61082\,
            I => \N__61058\
        );

    \I__14202\ : InMux
    port map (
            O => \N__61081\,
            I => \N__61055\
        );

    \I__14201\ : InMux
    port map (
            O => \N__61080\,
            I => \N__61048\
        );

    \I__14200\ : InMux
    port map (
            O => \N__61079\,
            I => \N__61048\
        );

    \I__14199\ : InMux
    port map (
            O => \N__61078\,
            I => \N__61048\
        );

    \I__14198\ : InMux
    port map (
            O => \N__61077\,
            I => \N__61045\
        );

    \I__14197\ : InMux
    port map (
            O => \N__61074\,
            I => \N__61040\
        );

    \I__14196\ : InMux
    port map (
            O => \N__61073\,
            I => \N__61040\
        );

    \I__14195\ : Span4Mux_h
    port map (
            O => \N__61070\,
            I => \N__61033\
        );

    \I__14194\ : Span4Mux_h
    port map (
            O => \N__61067\,
            I => \N__61033\
        );

    \I__14193\ : LocalMux
    port map (
            O => \N__61064\,
            I => \N__61033\
        );

    \I__14192\ : Odrv4
    port map (
            O => \N__61061\,
            I => data_in_frame_0_2
        );

    \I__14191\ : Odrv4
    port map (
            O => \N__61058\,
            I => data_in_frame_0_2
        );

    \I__14190\ : LocalMux
    port map (
            O => \N__61055\,
            I => data_in_frame_0_2
        );

    \I__14189\ : LocalMux
    port map (
            O => \N__61048\,
            I => data_in_frame_0_2
        );

    \I__14188\ : LocalMux
    port map (
            O => \N__61045\,
            I => data_in_frame_0_2
        );

    \I__14187\ : LocalMux
    port map (
            O => \N__61040\,
            I => data_in_frame_0_2
        );

    \I__14186\ : Odrv4
    port map (
            O => \N__61033\,
            I => data_in_frame_0_2
        );

    \I__14185\ : InMux
    port map (
            O => \N__61018\,
            I => \N__61015\
        );

    \I__14184\ : LocalMux
    port map (
            O => \N__61015\,
            I => \c0.n7\
        );

    \I__14183\ : CascadeMux
    port map (
            O => \N__61012\,
            I => \N__61008\
        );

    \I__14182\ : CascadeMux
    port map (
            O => \N__61011\,
            I => \N__61005\
        );

    \I__14181\ : InMux
    port map (
            O => \N__61008\,
            I => \N__61002\
        );

    \I__14180\ : InMux
    port map (
            O => \N__61005\,
            I => \N__60999\
        );

    \I__14179\ : LocalMux
    port map (
            O => \N__61002\,
            I => \N__60994\
        );

    \I__14178\ : LocalMux
    port map (
            O => \N__60999\,
            I => \N__60994\
        );

    \I__14177\ : Span4Mux_h
    port map (
            O => \N__60994\,
            I => \N__60991\
        );

    \I__14176\ : Odrv4
    port map (
            O => \N__60991\,
            I => \c0.n19241\
        );

    \I__14175\ : CascadeMux
    port map (
            O => \N__60988\,
            I => \N__60984\
        );

    \I__14174\ : InMux
    port map (
            O => \N__60987\,
            I => \N__60980\
        );

    \I__14173\ : InMux
    port map (
            O => \N__60984\,
            I => \N__60977\
        );

    \I__14172\ : CascadeMux
    port map (
            O => \N__60983\,
            I => \N__60973\
        );

    \I__14171\ : LocalMux
    port map (
            O => \N__60980\,
            I => \N__60970\
        );

    \I__14170\ : LocalMux
    port map (
            O => \N__60977\,
            I => \N__60967\
        );

    \I__14169\ : InMux
    port map (
            O => \N__60976\,
            I => \N__60964\
        );

    \I__14168\ : InMux
    port map (
            O => \N__60973\,
            I => \N__60961\
        );

    \I__14167\ : Span4Mux_h
    port map (
            O => \N__60970\,
            I => \N__60958\
        );

    \I__14166\ : Span4Mux_h
    port map (
            O => \N__60967\,
            I => \N__60953\
        );

    \I__14165\ : LocalMux
    port map (
            O => \N__60964\,
            I => \N__60950\
        );

    \I__14164\ : LocalMux
    port map (
            O => \N__60961\,
            I => \N__60945\
        );

    \I__14163\ : Span4Mux_h
    port map (
            O => \N__60958\,
            I => \N__60945\
        );

    \I__14162\ : InMux
    port map (
            O => \N__60957\,
            I => \N__60940\
        );

    \I__14161\ : InMux
    port map (
            O => \N__60956\,
            I => \N__60940\
        );

    \I__14160\ : Odrv4
    port map (
            O => \N__60953\,
            I => \c0.data_in_frame_2_4\
        );

    \I__14159\ : Odrv12
    port map (
            O => \N__60950\,
            I => \c0.data_in_frame_2_4\
        );

    \I__14158\ : Odrv4
    port map (
            O => \N__60945\,
            I => \c0.data_in_frame_2_4\
        );

    \I__14157\ : LocalMux
    port map (
            O => \N__60940\,
            I => \c0.data_in_frame_2_4\
        );

    \I__14156\ : InMux
    port map (
            O => \N__60931\,
            I => \N__60928\
        );

    \I__14155\ : LocalMux
    port map (
            O => \N__60928\,
            I => \N__60923\
        );

    \I__14154\ : InMux
    port map (
            O => \N__60927\,
            I => \N__60917\
        );

    \I__14153\ : InMux
    port map (
            O => \N__60926\,
            I => \N__60917\
        );

    \I__14152\ : Span4Mux_v
    port map (
            O => \N__60923\,
            I => \N__60913\
        );

    \I__14151\ : InMux
    port map (
            O => \N__60922\,
            I => \N__60910\
        );

    \I__14150\ : LocalMux
    port map (
            O => \N__60917\,
            I => \N__60902\
        );

    \I__14149\ : InMux
    port map (
            O => \N__60916\,
            I => \N__60896\
        );

    \I__14148\ : Span4Mux_h
    port map (
            O => \N__60913\,
            I => \N__60893\
        );

    \I__14147\ : LocalMux
    port map (
            O => \N__60910\,
            I => \N__60890\
        );

    \I__14146\ : InMux
    port map (
            O => \N__60909\,
            I => \N__60887\
        );

    \I__14145\ : InMux
    port map (
            O => \N__60908\,
            I => \N__60884\
        );

    \I__14144\ : InMux
    port map (
            O => \N__60907\,
            I => \N__60881\
        );

    \I__14143\ : InMux
    port map (
            O => \N__60906\,
            I => \N__60876\
        );

    \I__14142\ : InMux
    port map (
            O => \N__60905\,
            I => \N__60876\
        );

    \I__14141\ : Span4Mux_h
    port map (
            O => \N__60902\,
            I => \N__60873\
        );

    \I__14140\ : InMux
    port map (
            O => \N__60901\,
            I => \N__60868\
        );

    \I__14139\ : InMux
    port map (
            O => \N__60900\,
            I => \N__60868\
        );

    \I__14138\ : InMux
    port map (
            O => \N__60899\,
            I => \N__60865\
        );

    \I__14137\ : LocalMux
    port map (
            O => \N__60896\,
            I => data_in_frame_1_4
        );

    \I__14136\ : Odrv4
    port map (
            O => \N__60893\,
            I => data_in_frame_1_4
        );

    \I__14135\ : Odrv4
    port map (
            O => \N__60890\,
            I => data_in_frame_1_4
        );

    \I__14134\ : LocalMux
    port map (
            O => \N__60887\,
            I => data_in_frame_1_4
        );

    \I__14133\ : LocalMux
    port map (
            O => \N__60884\,
            I => data_in_frame_1_4
        );

    \I__14132\ : LocalMux
    port map (
            O => \N__60881\,
            I => data_in_frame_1_4
        );

    \I__14131\ : LocalMux
    port map (
            O => \N__60876\,
            I => data_in_frame_1_4
        );

    \I__14130\ : Odrv4
    port map (
            O => \N__60873\,
            I => data_in_frame_1_4
        );

    \I__14129\ : LocalMux
    port map (
            O => \N__60868\,
            I => data_in_frame_1_4
        );

    \I__14128\ : LocalMux
    port map (
            O => \N__60865\,
            I => data_in_frame_1_4
        );

    \I__14127\ : InMux
    port map (
            O => \N__60844\,
            I => \N__60839\
        );

    \I__14126\ : InMux
    port map (
            O => \N__60843\,
            I => \N__60836\
        );

    \I__14125\ : InMux
    port map (
            O => \N__60842\,
            I => \N__60833\
        );

    \I__14124\ : LocalMux
    port map (
            O => \N__60839\,
            I => \N__60830\
        );

    \I__14123\ : LocalMux
    port map (
            O => \N__60836\,
            I => \N__60826\
        );

    \I__14122\ : LocalMux
    port map (
            O => \N__60833\,
            I => \N__60823\
        );

    \I__14121\ : Span12Mux_h
    port map (
            O => \N__60830\,
            I => \N__60820\
        );

    \I__14120\ : InMux
    port map (
            O => \N__60829\,
            I => \N__60817\
        );

    \I__14119\ : Span4Mux_v
    port map (
            O => \N__60826\,
            I => \N__60814\
        );

    \I__14118\ : Span4Mux_h
    port map (
            O => \N__60823\,
            I => \N__60811\
        );

    \I__14117\ : Span12Mux_v
    port map (
            O => \N__60820\,
            I => \N__60808\
        );

    \I__14116\ : LocalMux
    port map (
            O => \N__60817\,
            I => \N__60805\
        );

    \I__14115\ : Span4Mux_v
    port map (
            O => \N__60814\,
            I => \N__60802\
        );

    \I__14114\ : Odrv4
    port map (
            O => \N__60811\,
            I => \c0.n11833\
        );

    \I__14113\ : Odrv12
    port map (
            O => \N__60808\,
            I => \c0.n11833\
        );

    \I__14112\ : Odrv4
    port map (
            O => \N__60805\,
            I => \c0.n11833\
        );

    \I__14111\ : Odrv4
    port map (
            O => \N__60802\,
            I => \c0.n11833\
        );

    \I__14110\ : InMux
    port map (
            O => \N__60793\,
            I => \N__60788\
        );

    \I__14109\ : InMux
    port map (
            O => \N__60792\,
            I => \N__60785\
        );

    \I__14108\ : InMux
    port map (
            O => \N__60791\,
            I => \N__60782\
        );

    \I__14107\ : LocalMux
    port map (
            O => \N__60788\,
            I => \N__60779\
        );

    \I__14106\ : LocalMux
    port map (
            O => \N__60785\,
            I => \N__60775\
        );

    \I__14105\ : LocalMux
    port map (
            O => \N__60782\,
            I => \N__60772\
        );

    \I__14104\ : Span4Mux_v
    port map (
            O => \N__60779\,
            I => \N__60768\
        );

    \I__14103\ : InMux
    port map (
            O => \N__60778\,
            I => \N__60765\
        );

    \I__14102\ : Span4Mux_h
    port map (
            O => \N__60775\,
            I => \N__60762\
        );

    \I__14101\ : Span4Mux_v
    port map (
            O => \N__60772\,
            I => \N__60759\
        );

    \I__14100\ : InMux
    port map (
            O => \N__60771\,
            I => \N__60756\
        );

    \I__14099\ : Odrv4
    port map (
            O => \N__60768\,
            I => \c0.n19456\
        );

    \I__14098\ : LocalMux
    port map (
            O => \N__60765\,
            I => \c0.n19456\
        );

    \I__14097\ : Odrv4
    port map (
            O => \N__60762\,
            I => \c0.n19456\
        );

    \I__14096\ : Odrv4
    port map (
            O => \N__60759\,
            I => \c0.n19456\
        );

    \I__14095\ : LocalMux
    port map (
            O => \N__60756\,
            I => \c0.n19456\
        );

    \I__14094\ : InMux
    port map (
            O => \N__60745\,
            I => \N__60742\
        );

    \I__14093\ : LocalMux
    port map (
            O => \N__60742\,
            I => \N__60739\
        );

    \I__14092\ : Span4Mux_v
    port map (
            O => \N__60739\,
            I => \N__60736\
        );

    \I__14091\ : Odrv4
    port map (
            O => \N__60736\,
            I => \c0.n5595\
        );

    \I__14090\ : InMux
    port map (
            O => \N__60733\,
            I => \N__60730\
        );

    \I__14089\ : LocalMux
    port map (
            O => \N__60730\,
            I => \N__60726\
        );

    \I__14088\ : InMux
    port map (
            O => \N__60729\,
            I => \N__60723\
        );

    \I__14087\ : Span4Mux_v
    port map (
            O => \N__60726\,
            I => \N__60718\
        );

    \I__14086\ : LocalMux
    port map (
            O => \N__60723\,
            I => \N__60718\
        );

    \I__14085\ : Span4Mux_h
    port map (
            O => \N__60718\,
            I => \N__60714\
        );

    \I__14084\ : InMux
    port map (
            O => \N__60717\,
            I => \N__60711\
        );

    \I__14083\ : Span4Mux_v
    port map (
            O => \N__60714\,
            I => \N__60704\
        );

    \I__14082\ : LocalMux
    port map (
            O => \N__60711\,
            I => \N__60704\
        );

    \I__14081\ : InMux
    port map (
            O => \N__60710\,
            I => \N__60699\
        );

    \I__14080\ : InMux
    port map (
            O => \N__60709\,
            I => \N__60699\
        );

    \I__14079\ : Span4Mux_h
    port map (
            O => \N__60704\,
            I => \N__60696\
        );

    \I__14078\ : LocalMux
    port map (
            O => \N__60699\,
            I => \N__60683\
        );

    \I__14077\ : Span4Mux_v
    port map (
            O => \N__60696\,
            I => \N__60680\
        );

    \I__14076\ : InMux
    port map (
            O => \N__60695\,
            I => \N__60677\
        );

    \I__14075\ : InMux
    port map (
            O => \N__60694\,
            I => \N__60668\
        );

    \I__14074\ : InMux
    port map (
            O => \N__60693\,
            I => \N__60668\
        );

    \I__14073\ : InMux
    port map (
            O => \N__60692\,
            I => \N__60668\
        );

    \I__14072\ : InMux
    port map (
            O => \N__60691\,
            I => \N__60668\
        );

    \I__14071\ : InMux
    port map (
            O => \N__60690\,
            I => \N__60663\
        );

    \I__14070\ : InMux
    port map (
            O => \N__60689\,
            I => \N__60663\
        );

    \I__14069\ : InMux
    port map (
            O => \N__60688\,
            I => \N__60660\
        );

    \I__14068\ : InMux
    port map (
            O => \N__60687\,
            I => \N__60655\
        );

    \I__14067\ : InMux
    port map (
            O => \N__60686\,
            I => \N__60655\
        );

    \I__14066\ : Span4Mux_v
    port map (
            O => \N__60683\,
            I => \N__60647\
        );

    \I__14065\ : Span4Mux_v
    port map (
            O => \N__60680\,
            I => \N__60644\
        );

    \I__14064\ : LocalMux
    port map (
            O => \N__60677\,
            I => \N__60641\
        );

    \I__14063\ : LocalMux
    port map (
            O => \N__60668\,
            I => \N__60636\
        );

    \I__14062\ : LocalMux
    port map (
            O => \N__60663\,
            I => \N__60636\
        );

    \I__14061\ : LocalMux
    port map (
            O => \N__60660\,
            I => \N__60629\
        );

    \I__14060\ : LocalMux
    port map (
            O => \N__60655\,
            I => \N__60626\
        );

    \I__14059\ : InMux
    port map (
            O => \N__60654\,
            I => \N__60621\
        );

    \I__14058\ : InMux
    port map (
            O => \N__60653\,
            I => \N__60621\
        );

    \I__14057\ : InMux
    port map (
            O => \N__60652\,
            I => \N__60612\
        );

    \I__14056\ : InMux
    port map (
            O => \N__60651\,
            I => \N__60612\
        );

    \I__14055\ : InMux
    port map (
            O => \N__60650\,
            I => \N__60609\
        );

    \I__14054\ : Sp12to4
    port map (
            O => \N__60647\,
            I => \N__60606\
        );

    \I__14053\ : Span4Mux_v
    port map (
            O => \N__60644\,
            I => \N__60603\
        );

    \I__14052\ : Span4Mux_v
    port map (
            O => \N__60641\,
            I => \N__60600\
        );

    \I__14051\ : Span4Mux_v
    port map (
            O => \N__60636\,
            I => \N__60597\
        );

    \I__14050\ : InMux
    port map (
            O => \N__60635\,
            I => \N__60592\
        );

    \I__14049\ : InMux
    port map (
            O => \N__60634\,
            I => \N__60592\
        );

    \I__14048\ : InMux
    port map (
            O => \N__60633\,
            I => \N__60589\
        );

    \I__14047\ : InMux
    port map (
            O => \N__60632\,
            I => \N__60586\
        );

    \I__14046\ : Span4Mux_v
    port map (
            O => \N__60629\,
            I => \N__60576\
        );

    \I__14045\ : Span4Mux_h
    port map (
            O => \N__60626\,
            I => \N__60576\
        );

    \I__14044\ : LocalMux
    port map (
            O => \N__60621\,
            I => \N__60576\
        );

    \I__14043\ : InMux
    port map (
            O => \N__60620\,
            I => \N__60567\
        );

    \I__14042\ : InMux
    port map (
            O => \N__60619\,
            I => \N__60567\
        );

    \I__14041\ : InMux
    port map (
            O => \N__60618\,
            I => \N__60567\
        );

    \I__14040\ : InMux
    port map (
            O => \N__60617\,
            I => \N__60567\
        );

    \I__14039\ : LocalMux
    port map (
            O => \N__60612\,
            I => \N__60560\
        );

    \I__14038\ : LocalMux
    port map (
            O => \N__60609\,
            I => \N__60560\
        );

    \I__14037\ : Span12Mux_h
    port map (
            O => \N__60606\,
            I => \N__60560\
        );

    \I__14036\ : Span4Mux_v
    port map (
            O => \N__60603\,
            I => \N__60555\
        );

    \I__14035\ : Span4Mux_h
    port map (
            O => \N__60600\,
            I => \N__60555\
        );

    \I__14034\ : Span4Mux_v
    port map (
            O => \N__60597\,
            I => \N__60552\
        );

    \I__14033\ : LocalMux
    port map (
            O => \N__60592\,
            I => \N__60549\
        );

    \I__14032\ : LocalMux
    port map (
            O => \N__60589\,
            I => \N__60546\
        );

    \I__14031\ : LocalMux
    port map (
            O => \N__60586\,
            I => \N__60543\
        );

    \I__14030\ : InMux
    port map (
            O => \N__60585\,
            I => \N__60538\
        );

    \I__14029\ : InMux
    port map (
            O => \N__60584\,
            I => \N__60538\
        );

    \I__14028\ : InMux
    port map (
            O => \N__60583\,
            I => \N__60535\
        );

    \I__14027\ : Sp12to4
    port map (
            O => \N__60576\,
            I => \N__60528\
        );

    \I__14026\ : LocalMux
    port map (
            O => \N__60567\,
            I => \N__60528\
        );

    \I__14025\ : Span12Mux_v
    port map (
            O => \N__60560\,
            I => \N__60528\
        );

    \I__14024\ : Odrv4
    port map (
            O => \N__60555\,
            I => n2108
        );

    \I__14023\ : Odrv4
    port map (
            O => \N__60552\,
            I => n2108
        );

    \I__14022\ : Odrv12
    port map (
            O => \N__60549\,
            I => n2108
        );

    \I__14021\ : Odrv4
    port map (
            O => \N__60546\,
            I => n2108
        );

    \I__14020\ : Odrv4
    port map (
            O => \N__60543\,
            I => n2108
        );

    \I__14019\ : LocalMux
    port map (
            O => \N__60538\,
            I => n2108
        );

    \I__14018\ : LocalMux
    port map (
            O => \N__60535\,
            I => n2108
        );

    \I__14017\ : Odrv12
    port map (
            O => \N__60528\,
            I => n2108
        );

    \I__14016\ : SRMux
    port map (
            O => \N__60511\,
            I => \N__60508\
        );

    \I__14015\ : LocalMux
    port map (
            O => \N__60508\,
            I => \N__60505\
        );

    \I__14014\ : Span4Mux_h
    port map (
            O => \N__60505\,
            I => \N__60502\
        );

    \I__14013\ : Span4Mux_h
    port map (
            O => \N__60502\,
            I => \N__60499\
        );

    \I__14012\ : Span4Mux_h
    port map (
            O => \N__60499\,
            I => \N__60496\
        );

    \I__14011\ : Odrv4
    port map (
            O => \N__60496\,
            I => \c0.n6_adj_3140\
        );

    \I__14010\ : CascadeMux
    port map (
            O => \N__60493\,
            I => \N__60489\
        );

    \I__14009\ : InMux
    port map (
            O => \N__60492\,
            I => \N__60482\
        );

    \I__14008\ : InMux
    port map (
            O => \N__60489\,
            I => \N__60482\
        );

    \I__14007\ : InMux
    port map (
            O => \N__60488\,
            I => \N__60479\
        );

    \I__14006\ : InMux
    port map (
            O => \N__60487\,
            I => \N__60475\
        );

    \I__14005\ : LocalMux
    port map (
            O => \N__60482\,
            I => \N__60472\
        );

    \I__14004\ : LocalMux
    port map (
            O => \N__60479\,
            I => \N__60469\
        );

    \I__14003\ : InMux
    port map (
            O => \N__60478\,
            I => \N__60466\
        );

    \I__14002\ : LocalMux
    port map (
            O => \N__60475\,
            I => \N__60461\
        );

    \I__14001\ : Span4Mux_h
    port map (
            O => \N__60472\,
            I => \N__60461\
        );

    \I__14000\ : Span4Mux_h
    port map (
            O => \N__60469\,
            I => \N__60458\
        );

    \I__13999\ : LocalMux
    port map (
            O => \N__60466\,
            I => \c0.data_in_frame_6_0\
        );

    \I__13998\ : Odrv4
    port map (
            O => \N__60461\,
            I => \c0.data_in_frame_6_0\
        );

    \I__13997\ : Odrv4
    port map (
            O => \N__60458\,
            I => \c0.data_in_frame_6_0\
        );

    \I__13996\ : InMux
    port map (
            O => \N__60451\,
            I => \N__60445\
        );

    \I__13995\ : InMux
    port map (
            O => \N__60450\,
            I => \N__60442\
        );

    \I__13994\ : CascadeMux
    port map (
            O => \N__60449\,
            I => \N__60439\
        );

    \I__13993\ : InMux
    port map (
            O => \N__60448\,
            I => \N__60436\
        );

    \I__13992\ : LocalMux
    port map (
            O => \N__60445\,
            I => \N__60433\
        );

    \I__13991\ : LocalMux
    port map (
            O => \N__60442\,
            I => \N__60430\
        );

    \I__13990\ : InMux
    port map (
            O => \N__60439\,
            I => \N__60427\
        );

    \I__13989\ : LocalMux
    port map (
            O => \N__60436\,
            I => \N__60422\
        );

    \I__13988\ : Span4Mux_h
    port map (
            O => \N__60433\,
            I => \N__60422\
        );

    \I__13987\ : Span4Mux_h
    port map (
            O => \N__60430\,
            I => \N__60419\
        );

    \I__13986\ : LocalMux
    port map (
            O => \N__60427\,
            I => \c0.data_in_frame_6_2\
        );

    \I__13985\ : Odrv4
    port map (
            O => \N__60422\,
            I => \c0.data_in_frame_6_2\
        );

    \I__13984\ : Odrv4
    port map (
            O => \N__60419\,
            I => \c0.data_in_frame_6_2\
        );

    \I__13983\ : InMux
    port map (
            O => \N__60412\,
            I => \N__60408\
        );

    \I__13982\ : InMux
    port map (
            O => \N__60411\,
            I => \N__60405\
        );

    \I__13981\ : LocalMux
    port map (
            O => \N__60408\,
            I => \N__60402\
        );

    \I__13980\ : LocalMux
    port map (
            O => \N__60405\,
            I => \N__60399\
        );

    \I__13979\ : Span4Mux_v
    port map (
            O => \N__60402\,
            I => \N__60395\
        );

    \I__13978\ : Span4Mux_h
    port map (
            O => \N__60399\,
            I => \N__60392\
        );

    \I__13977\ : InMux
    port map (
            O => \N__60398\,
            I => \N__60385\
        );

    \I__13976\ : Span4Mux_h
    port map (
            O => \N__60395\,
            I => \N__60382\
        );

    \I__13975\ : Span4Mux_h
    port map (
            O => \N__60392\,
            I => \N__60379\
        );

    \I__13974\ : InMux
    port map (
            O => \N__60391\,
            I => \N__60372\
        );

    \I__13973\ : InMux
    port map (
            O => \N__60390\,
            I => \N__60372\
        );

    \I__13972\ : InMux
    port map (
            O => \N__60389\,
            I => \N__60372\
        );

    \I__13971\ : InMux
    port map (
            O => \N__60388\,
            I => \N__60369\
        );

    \I__13970\ : LocalMux
    port map (
            O => \N__60385\,
            I => data_in_frame_1_2
        );

    \I__13969\ : Odrv4
    port map (
            O => \N__60382\,
            I => data_in_frame_1_2
        );

    \I__13968\ : Odrv4
    port map (
            O => \N__60379\,
            I => data_in_frame_1_2
        );

    \I__13967\ : LocalMux
    port map (
            O => \N__60372\,
            I => data_in_frame_1_2
        );

    \I__13966\ : LocalMux
    port map (
            O => \N__60369\,
            I => data_in_frame_1_2
        );

    \I__13965\ : CascadeMux
    port map (
            O => \N__60358\,
            I => \N__60355\
        );

    \I__13964\ : InMux
    port map (
            O => \N__60355\,
            I => \N__60347\
        );

    \I__13963\ : InMux
    port map (
            O => \N__60354\,
            I => \N__60347\
        );

    \I__13962\ : InMux
    port map (
            O => \N__60353\,
            I => \N__60343\
        );

    \I__13961\ : InMux
    port map (
            O => \N__60352\,
            I => \N__60340\
        );

    \I__13960\ : LocalMux
    port map (
            O => \N__60347\,
            I => \N__60337\
        );

    \I__13959\ : InMux
    port map (
            O => \N__60346\,
            I => \N__60333\
        );

    \I__13958\ : LocalMux
    port map (
            O => \N__60343\,
            I => \N__60330\
        );

    \I__13957\ : LocalMux
    port map (
            O => \N__60340\,
            I => \N__60326\
        );

    \I__13956\ : Span4Mux_v
    port map (
            O => \N__60337\,
            I => \N__60323\
        );

    \I__13955\ : InMux
    port map (
            O => \N__60336\,
            I => \N__60320\
        );

    \I__13954\ : LocalMux
    port map (
            O => \N__60333\,
            I => \N__60316\
        );

    \I__13953\ : Sp12to4
    port map (
            O => \N__60330\,
            I => \N__60313\
        );

    \I__13952\ : CascadeMux
    port map (
            O => \N__60329\,
            I => \N__60310\
        );

    \I__13951\ : Span4Mux_v
    port map (
            O => \N__60326\,
            I => \N__60302\
        );

    \I__13950\ : Span4Mux_h
    port map (
            O => \N__60323\,
            I => \N__60302\
        );

    \I__13949\ : LocalMux
    port map (
            O => \N__60320\,
            I => \N__60302\
        );

    \I__13948\ : InMux
    port map (
            O => \N__60319\,
            I => \N__60299\
        );

    \I__13947\ : Span4Mux_v
    port map (
            O => \N__60316\,
            I => \N__60296\
        );

    \I__13946\ : Span12Mux_s10_v
    port map (
            O => \N__60313\,
            I => \N__60293\
        );

    \I__13945\ : InMux
    port map (
            O => \N__60310\,
            I => \N__60288\
        );

    \I__13944\ : InMux
    port map (
            O => \N__60309\,
            I => \N__60288\
        );

    \I__13943\ : Span4Mux_h
    port map (
            O => \N__60302\,
            I => \N__60281\
        );

    \I__13942\ : LocalMux
    port map (
            O => \N__60299\,
            I => \N__60281\
        );

    \I__13941\ : Span4Mux_v
    port map (
            O => \N__60296\,
            I => \N__60281\
        );

    \I__13940\ : Odrv12
    port map (
            O => \N__60293\,
            I => \c0.n9_adj_3101\
        );

    \I__13939\ : LocalMux
    port map (
            O => \N__60288\,
            I => \c0.n9_adj_3101\
        );

    \I__13938\ : Odrv4
    port map (
            O => \N__60281\,
            I => \c0.n9_adj_3101\
        );

    \I__13937\ : InMux
    port map (
            O => \N__60274\,
            I => \N__60269\
        );

    \I__13936\ : InMux
    port map (
            O => \N__60273\,
            I => \N__60265\
        );

    \I__13935\ : InMux
    port map (
            O => \N__60272\,
            I => \N__60260\
        );

    \I__13934\ : LocalMux
    port map (
            O => \N__60269\,
            I => \N__60257\
        );

    \I__13933\ : InMux
    port map (
            O => \N__60268\,
            I => \N__60253\
        );

    \I__13932\ : LocalMux
    port map (
            O => \N__60265\,
            I => \N__60249\
        );

    \I__13931\ : CascadeMux
    port map (
            O => \N__60264\,
            I => \N__60246\
        );

    \I__13930\ : CascadeMux
    port map (
            O => \N__60263\,
            I => \N__60243\
        );

    \I__13929\ : LocalMux
    port map (
            O => \N__60260\,
            I => \N__60239\
        );

    \I__13928\ : Span4Mux_v
    port map (
            O => \N__60257\,
            I => \N__60236\
        );

    \I__13927\ : InMux
    port map (
            O => \N__60256\,
            I => \N__60232\
        );

    \I__13926\ : LocalMux
    port map (
            O => \N__60253\,
            I => \N__60229\
        );

    \I__13925\ : InMux
    port map (
            O => \N__60252\,
            I => \N__60226\
        );

    \I__13924\ : Span4Mux_v
    port map (
            O => \N__60249\,
            I => \N__60223\
        );

    \I__13923\ : InMux
    port map (
            O => \N__60246\,
            I => \N__60220\
        );

    \I__13922\ : InMux
    port map (
            O => \N__60243\,
            I => \N__60215\
        );

    \I__13921\ : InMux
    port map (
            O => \N__60242\,
            I => \N__60215\
        );

    \I__13920\ : Span4Mux_v
    port map (
            O => \N__60239\,
            I => \N__60212\
        );

    \I__13919\ : Span4Mux_v
    port map (
            O => \N__60236\,
            I => \N__60209\
        );

    \I__13918\ : CascadeMux
    port map (
            O => \N__60235\,
            I => \N__60205\
        );

    \I__13917\ : LocalMux
    port map (
            O => \N__60232\,
            I => \N__60201\
        );

    \I__13916\ : Span4Mux_v
    port map (
            O => \N__60229\,
            I => \N__60198\
        );

    \I__13915\ : LocalMux
    port map (
            O => \N__60226\,
            I => \N__60195\
        );

    \I__13914\ : Span4Mux_h
    port map (
            O => \N__60223\,
            I => \N__60192\
        );

    \I__13913\ : LocalMux
    port map (
            O => \N__60220\,
            I => \N__60189\
        );

    \I__13912\ : LocalMux
    port map (
            O => \N__60215\,
            I => \N__60186\
        );

    \I__13911\ : Span4Mux_v
    port map (
            O => \N__60212\,
            I => \N__60183\
        );

    \I__13910\ : Span4Mux_h
    port map (
            O => \N__60209\,
            I => \N__60180\
        );

    \I__13909\ : InMux
    port map (
            O => \N__60208\,
            I => \N__60177\
        );

    \I__13908\ : InMux
    port map (
            O => \N__60205\,
            I => \N__60174\
        );

    \I__13907\ : InMux
    port map (
            O => \N__60204\,
            I => \N__60171\
        );

    \I__13906\ : Span4Mux_v
    port map (
            O => \N__60201\,
            I => \N__60168\
        );

    \I__13905\ : Span4Mux_h
    port map (
            O => \N__60198\,
            I => \N__60163\
        );

    \I__13904\ : Span4Mux_v
    port map (
            O => \N__60195\,
            I => \N__60163\
        );

    \I__13903\ : Span4Mux_h
    port map (
            O => \N__60192\,
            I => \N__60154\
        );

    \I__13902\ : Span4Mux_v
    port map (
            O => \N__60189\,
            I => \N__60154\
        );

    \I__13901\ : Span4Mux_v
    port map (
            O => \N__60186\,
            I => \N__60154\
        );

    \I__13900\ : Span4Mux_v
    port map (
            O => \N__60183\,
            I => \N__60154\
        );

    \I__13899\ : Span4Mux_v
    port map (
            O => \N__60180\,
            I => \N__60151\
        );

    \I__13898\ : LocalMux
    port map (
            O => \N__60177\,
            I => \N__60148\
        );

    \I__13897\ : LocalMux
    port map (
            O => \N__60174\,
            I => \FRAME_MATCHER_i_0\
        );

    \I__13896\ : LocalMux
    port map (
            O => \N__60171\,
            I => \FRAME_MATCHER_i_0\
        );

    \I__13895\ : Odrv4
    port map (
            O => \N__60168\,
            I => \FRAME_MATCHER_i_0\
        );

    \I__13894\ : Odrv4
    port map (
            O => \N__60163\,
            I => \FRAME_MATCHER_i_0\
        );

    \I__13893\ : Odrv4
    port map (
            O => \N__60154\,
            I => \FRAME_MATCHER_i_0\
        );

    \I__13892\ : Odrv4
    port map (
            O => \N__60151\,
            I => \FRAME_MATCHER_i_0\
        );

    \I__13891\ : Odrv4
    port map (
            O => \N__60148\,
            I => \FRAME_MATCHER_i_0\
        );

    \I__13890\ : CascadeMux
    port map (
            O => \N__60133\,
            I => \N__60129\
        );

    \I__13889\ : InMux
    port map (
            O => \N__60132\,
            I => \N__60125\
        );

    \I__13888\ : InMux
    port map (
            O => \N__60129\,
            I => \N__60122\
        );

    \I__13887\ : InMux
    port map (
            O => \N__60128\,
            I => \N__60118\
        );

    \I__13886\ : LocalMux
    port map (
            O => \N__60125\,
            I => \N__60112\
        );

    \I__13885\ : LocalMux
    port map (
            O => \N__60122\,
            I => \N__60109\
        );

    \I__13884\ : InMux
    port map (
            O => \N__60121\,
            I => \N__60105\
        );

    \I__13883\ : LocalMux
    port map (
            O => \N__60118\,
            I => \N__60101\
        );

    \I__13882\ : InMux
    port map (
            O => \N__60117\,
            I => \N__60098\
        );

    \I__13881\ : InMux
    port map (
            O => \N__60116\,
            I => \N__60095\
        );

    \I__13880\ : InMux
    port map (
            O => \N__60115\,
            I => \N__60092\
        );

    \I__13879\ : Span4Mux_h
    port map (
            O => \N__60112\,
            I => \N__60089\
        );

    \I__13878\ : Span4Mux_v
    port map (
            O => \N__60109\,
            I => \N__60086\
        );

    \I__13877\ : InMux
    port map (
            O => \N__60108\,
            I => \N__60083\
        );

    \I__13876\ : LocalMux
    port map (
            O => \N__60105\,
            I => \N__60080\
        );

    \I__13875\ : InMux
    port map (
            O => \N__60104\,
            I => \N__60077\
        );

    \I__13874\ : Span4Mux_h
    port map (
            O => \N__60101\,
            I => \N__60072\
        );

    \I__13873\ : LocalMux
    port map (
            O => \N__60098\,
            I => \N__60072\
        );

    \I__13872\ : LocalMux
    port map (
            O => \N__60095\,
            I => \N__60069\
        );

    \I__13871\ : LocalMux
    port map (
            O => \N__60092\,
            I => \N__60064\
        );

    \I__13870\ : Span4Mux_h
    port map (
            O => \N__60089\,
            I => \N__60064\
        );

    \I__13869\ : Sp12to4
    port map (
            O => \N__60086\,
            I => \N__60061\
        );

    \I__13868\ : LocalMux
    port map (
            O => \N__60083\,
            I => \N__60058\
        );

    \I__13867\ : Span4Mux_v
    port map (
            O => \N__60080\,
            I => \N__60053\
        );

    \I__13866\ : LocalMux
    port map (
            O => \N__60077\,
            I => \N__60053\
        );

    \I__13865\ : Span4Mux_v
    port map (
            O => \N__60072\,
            I => \N__60050\
        );

    \I__13864\ : Span4Mux_h
    port map (
            O => \N__60069\,
            I => \N__60042\
        );

    \I__13863\ : Span4Mux_v
    port map (
            O => \N__60064\,
            I => \N__60042\
        );

    \I__13862\ : Span12Mux_h
    port map (
            O => \N__60061\,
            I => \N__60038\
        );

    \I__13861\ : Span4Mux_h
    port map (
            O => \N__60058\,
            I => \N__60035\
        );

    \I__13860\ : Span4Mux_v
    port map (
            O => \N__60053\,
            I => \N__60032\
        );

    \I__13859\ : Sp12to4
    port map (
            O => \N__60050\,
            I => \N__60029\
        );

    \I__13858\ : InMux
    port map (
            O => \N__60049\,
            I => \N__60022\
        );

    \I__13857\ : InMux
    port map (
            O => \N__60048\,
            I => \N__60022\
        );

    \I__13856\ : InMux
    port map (
            O => \N__60047\,
            I => \N__60022\
        );

    \I__13855\ : Sp12to4
    port map (
            O => \N__60042\,
            I => \N__60019\
        );

    \I__13854\ : InMux
    port map (
            O => \N__60041\,
            I => \N__60016\
        );

    \I__13853\ : Odrv12
    port map (
            O => \N__60038\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__13852\ : Odrv4
    port map (
            O => \N__60035\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__13851\ : Odrv4
    port map (
            O => \N__60032\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__13850\ : Odrv12
    port map (
            O => \N__60029\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__13849\ : LocalMux
    port map (
            O => \N__60022\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__13848\ : Odrv12
    port map (
            O => \N__60019\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__13847\ : LocalMux
    port map (
            O => \N__60016\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__13846\ : InMux
    port map (
            O => \N__60001\,
            I => \N__59997\
        );

    \I__13845\ : InMux
    port map (
            O => \N__60000\,
            I => \N__59993\
        );

    \I__13844\ : LocalMux
    port map (
            O => \N__59997\,
            I => \N__59989\
        );

    \I__13843\ : InMux
    port map (
            O => \N__59996\,
            I => \N__59986\
        );

    \I__13842\ : LocalMux
    port map (
            O => \N__59993\,
            I => \N__59982\
        );

    \I__13841\ : InMux
    port map (
            O => \N__59992\,
            I => \N__59979\
        );

    \I__13840\ : Span4Mux_v
    port map (
            O => \N__59989\,
            I => \N__59972\
        );

    \I__13839\ : LocalMux
    port map (
            O => \N__59986\,
            I => \N__59972\
        );

    \I__13838\ : InMux
    port map (
            O => \N__59985\,
            I => \N__59969\
        );

    \I__13837\ : Span4Mux_h
    port map (
            O => \N__59982\,
            I => \N__59966\
        );

    \I__13836\ : LocalMux
    port map (
            O => \N__59979\,
            I => \N__59962\
        );

    \I__13835\ : InMux
    port map (
            O => \N__59978\,
            I => \N__59959\
        );

    \I__13834\ : InMux
    port map (
            O => \N__59977\,
            I => \N__59956\
        );

    \I__13833\ : Span4Mux_h
    port map (
            O => \N__59972\,
            I => \N__59951\
        );

    \I__13832\ : LocalMux
    port map (
            O => \N__59969\,
            I => \N__59951\
        );

    \I__13831\ : Span4Mux_h
    port map (
            O => \N__59966\,
            I => \N__59948\
        );

    \I__13830\ : CascadeMux
    port map (
            O => \N__59965\,
            I => \N__59945\
        );

    \I__13829\ : Span4Mux_v
    port map (
            O => \N__59962\,
            I => \N__59939\
        );

    \I__13828\ : LocalMux
    port map (
            O => \N__59959\,
            I => \N__59939\
        );

    \I__13827\ : LocalMux
    port map (
            O => \N__59956\,
            I => \N__59934\
        );

    \I__13826\ : Span4Mux_h
    port map (
            O => \N__59951\,
            I => \N__59934\
        );

    \I__13825\ : Span4Mux_v
    port map (
            O => \N__59948\,
            I => \N__59931\
        );

    \I__13824\ : InMux
    port map (
            O => \N__59945\,
            I => \N__59928\
        );

    \I__13823\ : CascadeMux
    port map (
            O => \N__59944\,
            I => \N__59924\
        );

    \I__13822\ : Span4Mux_h
    port map (
            O => \N__59939\,
            I => \N__59914\
        );

    \I__13821\ : Span4Mux_h
    port map (
            O => \N__59934\,
            I => \N__59914\
        );

    \I__13820\ : Span4Mux_v
    port map (
            O => \N__59931\,
            I => \N__59914\
        );

    \I__13819\ : LocalMux
    port map (
            O => \N__59928\,
            I => \N__59911\
        );

    \I__13818\ : InMux
    port map (
            O => \N__59927\,
            I => \N__59908\
        );

    \I__13817\ : InMux
    port map (
            O => \N__59924\,
            I => \N__59899\
        );

    \I__13816\ : InMux
    port map (
            O => \N__59923\,
            I => \N__59899\
        );

    \I__13815\ : InMux
    port map (
            O => \N__59922\,
            I => \N__59899\
        );

    \I__13814\ : InMux
    port map (
            O => \N__59921\,
            I => \N__59899\
        );

    \I__13813\ : Span4Mux_v
    port map (
            O => \N__59914\,
            I => \N__59896\
        );

    \I__13812\ : Span12Mux_v
    port map (
            O => \N__59911\,
            I => \N__59893\
        );

    \I__13811\ : LocalMux
    port map (
            O => \N__59908\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__13810\ : LocalMux
    port map (
            O => \N__59899\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__13809\ : Odrv4
    port map (
            O => \N__59896\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__13808\ : Odrv12
    port map (
            O => \N__59893\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__13807\ : InMux
    port map (
            O => \N__59884\,
            I => \N__59880\
        );

    \I__13806\ : InMux
    port map (
            O => \N__59883\,
            I => \N__59877\
        );

    \I__13805\ : LocalMux
    port map (
            O => \N__59880\,
            I => \N__59870\
        );

    \I__13804\ : LocalMux
    port map (
            O => \N__59877\,
            I => \N__59870\
        );

    \I__13803\ : InMux
    port map (
            O => \N__59876\,
            I => \N__59861\
        );

    \I__13802\ : InMux
    port map (
            O => \N__59875\,
            I => \N__59861\
        );

    \I__13801\ : Span4Mux_h
    port map (
            O => \N__59870\,
            I => \N__59858\
        );

    \I__13800\ : InMux
    port map (
            O => \N__59869\,
            I => \N__59855\
        );

    \I__13799\ : InMux
    port map (
            O => \N__59868\,
            I => \N__59848\
        );

    \I__13798\ : InMux
    port map (
            O => \N__59867\,
            I => \N__59848\
        );

    \I__13797\ : InMux
    port map (
            O => \N__59866\,
            I => \N__59848\
        );

    \I__13796\ : LocalMux
    port map (
            O => \N__59861\,
            I => \N__59845\
        );

    \I__13795\ : Span4Mux_h
    port map (
            O => \N__59858\,
            I => \N__59842\
        );

    \I__13794\ : LocalMux
    port map (
            O => \N__59855\,
            I => n19100
        );

    \I__13793\ : LocalMux
    port map (
            O => \N__59848\,
            I => n19100
        );

    \I__13792\ : Odrv12
    port map (
            O => \N__59845\,
            I => n19100
        );

    \I__13791\ : Odrv4
    port map (
            O => \N__59842\,
            I => n19100
        );

    \I__13790\ : InMux
    port map (
            O => \N__59833\,
            I => \N__59829\
        );

    \I__13789\ : InMux
    port map (
            O => \N__59832\,
            I => \N__59825\
        );

    \I__13788\ : LocalMux
    port map (
            O => \N__59829\,
            I => \N__59822\
        );

    \I__13787\ : InMux
    port map (
            O => \N__59828\,
            I => \N__59819\
        );

    \I__13786\ : LocalMux
    port map (
            O => \N__59825\,
            I => \c0.n17942\
        );

    \I__13785\ : Odrv12
    port map (
            O => \N__59822\,
            I => \c0.n17942\
        );

    \I__13784\ : LocalMux
    port map (
            O => \N__59819\,
            I => \c0.n17942\
        );

    \I__13783\ : CascadeMux
    port map (
            O => \N__59812\,
            I => \c0.n77_adj_3396_cascade_\
        );

    \I__13782\ : InMux
    port map (
            O => \N__59809\,
            I => \N__59806\
        );

    \I__13781\ : LocalMux
    port map (
            O => \N__59806\,
            I => \N__59803\
        );

    \I__13780\ : Span4Mux_h
    port map (
            O => \N__59803\,
            I => \N__59800\
        );

    \I__13779\ : Span4Mux_v
    port map (
            O => \N__59800\,
            I => \N__59797\
        );

    \I__13778\ : Odrv4
    port map (
            O => \N__59797\,
            I => \c0.n90_adj_3400\
        );

    \I__13777\ : CascadeMux
    port map (
            O => \N__59794\,
            I => \N__59791\
        );

    \I__13776\ : InMux
    port map (
            O => \N__59791\,
            I => \N__59788\
        );

    \I__13775\ : LocalMux
    port map (
            O => \N__59788\,
            I => \N__59785\
        );

    \I__13774\ : Span4Mux_v
    port map (
            O => \N__59785\,
            I => \N__59780\
        );

    \I__13773\ : CascadeMux
    port map (
            O => \N__59784\,
            I => \N__59776\
        );

    \I__13772\ : CascadeMux
    port map (
            O => \N__59783\,
            I => \N__59772\
        );

    \I__13771\ : Span4Mux_h
    port map (
            O => \N__59780\,
            I => \N__59769\
        );

    \I__13770\ : InMux
    port map (
            O => \N__59779\,
            I => \N__59766\
        );

    \I__13769\ : InMux
    port map (
            O => \N__59776\,
            I => \N__59763\
        );

    \I__13768\ : InMux
    port map (
            O => \N__59775\,
            I => \N__59760\
        );

    \I__13767\ : InMux
    port map (
            O => \N__59772\,
            I => \N__59757\
        );

    \I__13766\ : Sp12to4
    port map (
            O => \N__59769\,
            I => \N__59748\
        );

    \I__13765\ : LocalMux
    port map (
            O => \N__59766\,
            I => \N__59748\
        );

    \I__13764\ : LocalMux
    port map (
            O => \N__59763\,
            I => \N__59748\
        );

    \I__13763\ : LocalMux
    port map (
            O => \N__59760\,
            I => \N__59748\
        );

    \I__13762\ : LocalMux
    port map (
            O => \N__59757\,
            I => \c0.data_in_frame_25_7\
        );

    \I__13761\ : Odrv12
    port map (
            O => \N__59748\,
            I => \c0.data_in_frame_25_7\
        );

    \I__13760\ : InMux
    port map (
            O => \N__59743\,
            I => \N__59739\
        );

    \I__13759\ : InMux
    port map (
            O => \N__59742\,
            I => \N__59735\
        );

    \I__13758\ : LocalMux
    port map (
            O => \N__59739\,
            I => \N__59732\
        );

    \I__13757\ : InMux
    port map (
            O => \N__59738\,
            I => \N__59729\
        );

    \I__13756\ : LocalMux
    port map (
            O => \N__59735\,
            I => \N__59726\
        );

    \I__13755\ : Span4Mux_v
    port map (
            O => \N__59732\,
            I => \N__59723\
        );

    \I__13754\ : LocalMux
    port map (
            O => \N__59729\,
            I => \N__59720\
        );

    \I__13753\ : Span4Mux_v
    port map (
            O => \N__59726\,
            I => \N__59712\
        );

    \I__13752\ : Span4Mux_h
    port map (
            O => \N__59723\,
            I => \N__59712\
        );

    \I__13751\ : Span4Mux_v
    port map (
            O => \N__59720\,
            I => \N__59712\
        );

    \I__13750\ : InMux
    port map (
            O => \N__59719\,
            I => \N__59709\
        );

    \I__13749\ : Span4Mux_v
    port map (
            O => \N__59712\,
            I => \N__59706\
        );

    \I__13748\ : LocalMux
    port map (
            O => \N__59709\,
            I => \c0.data_in_frame_25_5\
        );

    \I__13747\ : Odrv4
    port map (
            O => \N__59706\,
            I => \c0.data_in_frame_25_5\
        );

    \I__13746\ : CascadeMux
    port map (
            O => \N__59701\,
            I => \N__59696\
        );

    \I__13745\ : InMux
    port map (
            O => \N__59700\,
            I => \N__59693\
        );

    \I__13744\ : InMux
    port map (
            O => \N__59699\,
            I => \N__59689\
        );

    \I__13743\ : InMux
    port map (
            O => \N__59696\,
            I => \N__59685\
        );

    \I__13742\ : LocalMux
    port map (
            O => \N__59693\,
            I => \N__59682\
        );

    \I__13741\ : CascadeMux
    port map (
            O => \N__59692\,
            I => \N__59679\
        );

    \I__13740\ : LocalMux
    port map (
            O => \N__59689\,
            I => \N__59676\
        );

    \I__13739\ : InMux
    port map (
            O => \N__59688\,
            I => \N__59673\
        );

    \I__13738\ : LocalMux
    port map (
            O => \N__59685\,
            I => \N__59670\
        );

    \I__13737\ : Span4Mux_v
    port map (
            O => \N__59682\,
            I => \N__59666\
        );

    \I__13736\ : InMux
    port map (
            O => \N__59679\,
            I => \N__59663\
        );

    \I__13735\ : Span4Mux_v
    port map (
            O => \N__59676\,
            I => \N__59660\
        );

    \I__13734\ : LocalMux
    port map (
            O => \N__59673\,
            I => \N__59657\
        );

    \I__13733\ : Span4Mux_v
    port map (
            O => \N__59670\,
            I => \N__59654\
        );

    \I__13732\ : CascadeMux
    port map (
            O => \N__59669\,
            I => \N__59651\
        );

    \I__13731\ : Sp12to4
    port map (
            O => \N__59666\,
            I => \N__59644\
        );

    \I__13730\ : LocalMux
    port map (
            O => \N__59663\,
            I => \N__59644\
        );

    \I__13729\ : Sp12to4
    port map (
            O => \N__59660\,
            I => \N__59644\
        );

    \I__13728\ : Span4Mux_v
    port map (
            O => \N__59657\,
            I => \N__59639\
        );

    \I__13727\ : Span4Mux_h
    port map (
            O => \N__59654\,
            I => \N__59639\
        );

    \I__13726\ : InMux
    port map (
            O => \N__59651\,
            I => \N__59636\
        );

    \I__13725\ : Span12Mux_h
    port map (
            O => \N__59644\,
            I => \N__59633\
        );

    \I__13724\ : Span4Mux_v
    port map (
            O => \N__59639\,
            I => \N__59630\
        );

    \I__13723\ : LocalMux
    port map (
            O => \N__59636\,
            I => \c0.data_in_frame_25_4\
        );

    \I__13722\ : Odrv12
    port map (
            O => \N__59633\,
            I => \c0.data_in_frame_25_4\
        );

    \I__13721\ : Odrv4
    port map (
            O => \N__59630\,
            I => \c0.data_in_frame_25_4\
        );

    \I__13720\ : CascadeMux
    port map (
            O => \N__59623\,
            I => \c0.n19214_cascade_\
        );

    \I__13719\ : InMux
    port map (
            O => \N__59620\,
            I => \N__59617\
        );

    \I__13718\ : LocalMux
    port map (
            O => \N__59617\,
            I => \N__59613\
        );

    \I__13717\ : InMux
    port map (
            O => \N__59616\,
            I => \N__59609\
        );

    \I__13716\ : Span4Mux_h
    port map (
            O => \N__59613\,
            I => \N__59606\
        );

    \I__13715\ : InMux
    port map (
            O => \N__59612\,
            I => \N__59603\
        );

    \I__13714\ : LocalMux
    port map (
            O => \N__59609\,
            I => data_in_frame_24_5
        );

    \I__13713\ : Odrv4
    port map (
            O => \N__59606\,
            I => data_in_frame_24_5
        );

    \I__13712\ : LocalMux
    port map (
            O => \N__59603\,
            I => data_in_frame_24_5
        );

    \I__13711\ : InMux
    port map (
            O => \N__59596\,
            I => \N__59592\
        );

    \I__13710\ : InMux
    port map (
            O => \N__59595\,
            I => \N__59589\
        );

    \I__13709\ : LocalMux
    port map (
            O => \N__59592\,
            I => \N__59585\
        );

    \I__13708\ : LocalMux
    port map (
            O => \N__59589\,
            I => \N__59582\
        );

    \I__13707\ : InMux
    port map (
            O => \N__59588\,
            I => \N__59579\
        );

    \I__13706\ : Span4Mux_v
    port map (
            O => \N__59585\,
            I => \N__59576\
        );

    \I__13705\ : Span4Mux_v
    port map (
            O => \N__59582\,
            I => \N__59571\
        );

    \I__13704\ : LocalMux
    port map (
            O => \N__59579\,
            I => \N__59571\
        );

    \I__13703\ : Span4Mux_h
    port map (
            O => \N__59576\,
            I => \N__59568\
        );

    \I__13702\ : Span4Mux_h
    port map (
            O => \N__59571\,
            I => \N__59565\
        );

    \I__13701\ : Odrv4
    port map (
            O => \N__59568\,
            I => \c0.n12_adj_3214\
        );

    \I__13700\ : Odrv4
    port map (
            O => \N__59565\,
            I => \c0.n12_adj_3214\
        );

    \I__13699\ : InMux
    port map (
            O => \N__59560\,
            I => \N__59557\
        );

    \I__13698\ : LocalMux
    port map (
            O => \N__59557\,
            I => \N__59553\
        );

    \I__13697\ : CascadeMux
    port map (
            O => \N__59556\,
            I => \N__59550\
        );

    \I__13696\ : Span4Mux_h
    port map (
            O => \N__59553\,
            I => \N__59545\
        );

    \I__13695\ : InMux
    port map (
            O => \N__59550\,
            I => \N__59540\
        );

    \I__13694\ : InMux
    port map (
            O => \N__59549\,
            I => \N__59540\
        );

    \I__13693\ : InMux
    port map (
            O => \N__59548\,
            I => \N__59537\
        );

    \I__13692\ : Odrv4
    port map (
            O => \N__59545\,
            I => \c0.data_in_frame_25_6\
        );

    \I__13691\ : LocalMux
    port map (
            O => \N__59540\,
            I => \c0.data_in_frame_25_6\
        );

    \I__13690\ : LocalMux
    port map (
            O => \N__59537\,
            I => \c0.data_in_frame_25_6\
        );

    \I__13689\ : InMux
    port map (
            O => \N__59530\,
            I => \N__59527\
        );

    \I__13688\ : LocalMux
    port map (
            O => \N__59527\,
            I => \N__59524\
        );

    \I__13687\ : Span4Mux_h
    port map (
            O => \N__59524\,
            I => \N__59521\
        );

    \I__13686\ : Span4Mux_v
    port map (
            O => \N__59521\,
            I => \N__59518\
        );

    \I__13685\ : Span4Mux_v
    port map (
            O => \N__59518\,
            I => \N__59515\
        );

    \I__13684\ : Odrv4
    port map (
            O => \N__59515\,
            I => \c0.n5784\
        );

    \I__13683\ : InMux
    port map (
            O => \N__59512\,
            I => \N__59508\
        );

    \I__13682\ : InMux
    port map (
            O => \N__59511\,
            I => \N__59505\
        );

    \I__13681\ : LocalMux
    port map (
            O => \N__59508\,
            I => \N__59501\
        );

    \I__13680\ : LocalMux
    port map (
            O => \N__59505\,
            I => \N__59498\
        );

    \I__13679\ : InMux
    port map (
            O => \N__59504\,
            I => \N__59495\
        );

    \I__13678\ : Span4Mux_v
    port map (
            O => \N__59501\,
            I => \N__59488\
        );

    \I__13677\ : Span4Mux_v
    port map (
            O => \N__59498\,
            I => \N__59488\
        );

    \I__13676\ : LocalMux
    port map (
            O => \N__59495\,
            I => \N__59488\
        );

    \I__13675\ : Odrv4
    port map (
            O => \N__59488\,
            I => \c0.n18431\
        );

    \I__13674\ : InMux
    port map (
            O => \N__59485\,
            I => \N__59482\
        );

    \I__13673\ : LocalMux
    port map (
            O => \N__59482\,
            I => \N__59475\
        );

    \I__13672\ : InMux
    port map (
            O => \N__59481\,
            I => \N__59472\
        );

    \I__13671\ : InMux
    port map (
            O => \N__59480\,
            I => \N__59469\
        );

    \I__13670\ : InMux
    port map (
            O => \N__59479\,
            I => \N__59466\
        );

    \I__13669\ : InMux
    port map (
            O => \N__59478\,
            I => \N__59463\
        );

    \I__13668\ : Span4Mux_v
    port map (
            O => \N__59475\,
            I => \N__59460\
        );

    \I__13667\ : LocalMux
    port map (
            O => \N__59472\,
            I => \N__59456\
        );

    \I__13666\ : LocalMux
    port map (
            O => \N__59469\,
            I => \N__59452\
        );

    \I__13665\ : LocalMux
    port map (
            O => \N__59466\,
            I => \N__59449\
        );

    \I__13664\ : LocalMux
    port map (
            O => \N__59463\,
            I => \N__59443\
        );

    \I__13663\ : Span4Mux_v
    port map (
            O => \N__59460\,
            I => \N__59443\
        );

    \I__13662\ : InMux
    port map (
            O => \N__59459\,
            I => \N__59440\
        );

    \I__13661\ : Span4Mux_v
    port map (
            O => \N__59456\,
            I => \N__59436\
        );

    \I__13660\ : InMux
    port map (
            O => \N__59455\,
            I => \N__59433\
        );

    \I__13659\ : Span4Mux_h
    port map (
            O => \N__59452\,
            I => \N__59429\
        );

    \I__13658\ : Span4Mux_v
    port map (
            O => \N__59449\,
            I => \N__59426\
        );

    \I__13657\ : InMux
    port map (
            O => \N__59448\,
            I => \N__59423\
        );

    \I__13656\ : Span4Mux_h
    port map (
            O => \N__59443\,
            I => \N__59418\
        );

    \I__13655\ : LocalMux
    port map (
            O => \N__59440\,
            I => \N__59418\
        );

    \I__13654\ : InMux
    port map (
            O => \N__59439\,
            I => \N__59415\
        );

    \I__13653\ : Span4Mux_v
    port map (
            O => \N__59436\,
            I => \N__59412\
        );

    \I__13652\ : LocalMux
    port map (
            O => \N__59433\,
            I => \N__59409\
        );

    \I__13651\ : InMux
    port map (
            O => \N__59432\,
            I => \N__59406\
        );

    \I__13650\ : Span4Mux_v
    port map (
            O => \N__59429\,
            I => \N__59403\
        );

    \I__13649\ : Span4Mux_h
    port map (
            O => \N__59426\,
            I => \N__59396\
        );

    \I__13648\ : LocalMux
    port map (
            O => \N__59423\,
            I => \N__59396\
        );

    \I__13647\ : Span4Mux_v
    port map (
            O => \N__59418\,
            I => \N__59396\
        );

    \I__13646\ : LocalMux
    port map (
            O => \N__59415\,
            I => \N__59393\
        );

    \I__13645\ : Odrv4
    port map (
            O => \N__59412\,
            I => \c0.n15701\
        );

    \I__13644\ : Odrv4
    port map (
            O => \N__59409\,
            I => \c0.n15701\
        );

    \I__13643\ : LocalMux
    port map (
            O => \N__59406\,
            I => \c0.n15701\
        );

    \I__13642\ : Odrv4
    port map (
            O => \N__59403\,
            I => \c0.n15701\
        );

    \I__13641\ : Odrv4
    port map (
            O => \N__59396\,
            I => \c0.n15701\
        );

    \I__13640\ : Odrv4
    port map (
            O => \N__59393\,
            I => \c0.n15701\
        );

    \I__13639\ : InMux
    port map (
            O => \N__59380\,
            I => \N__59377\
        );

    \I__13638\ : LocalMux
    port map (
            O => \N__59377\,
            I => \N__59374\
        );

    \I__13637\ : Span4Mux_v
    port map (
            O => \N__59374\,
            I => \N__59371\
        );

    \I__13636\ : Span4Mux_h
    port map (
            O => \N__59371\,
            I => \N__59368\
        );

    \I__13635\ : Span4Mux_v
    port map (
            O => \N__59368\,
            I => \N__59365\
        );

    \I__13634\ : Span4Mux_h
    port map (
            O => \N__59365\,
            I => \N__59362\
        );

    \I__13633\ : Odrv4
    port map (
            O => \N__59362\,
            I => \c0.n7_adj_3047\
        );

    \I__13632\ : InMux
    port map (
            O => \N__59359\,
            I => \N__59355\
        );

    \I__13631\ : InMux
    port map (
            O => \N__59358\,
            I => \N__59352\
        );

    \I__13630\ : LocalMux
    port map (
            O => \N__59355\,
            I => \N__59349\
        );

    \I__13629\ : LocalMux
    port map (
            O => \N__59352\,
            I => \N__59346\
        );

    \I__13628\ : Span4Mux_h
    port map (
            O => \N__59349\,
            I => \N__59340\
        );

    \I__13627\ : Span4Mux_v
    port map (
            O => \N__59346\,
            I => \N__59340\
        );

    \I__13626\ : InMux
    port map (
            O => \N__59345\,
            I => \N__59337\
        );

    \I__13625\ : Odrv4
    port map (
            O => \N__59340\,
            I => \c0.n20965\
        );

    \I__13624\ : LocalMux
    port map (
            O => \N__59337\,
            I => \c0.n20965\
        );

    \I__13623\ : InMux
    port map (
            O => \N__59332\,
            I => \N__59329\
        );

    \I__13622\ : LocalMux
    port map (
            O => \N__59329\,
            I => \N__59326\
        );

    \I__13621\ : Span4Mux_h
    port map (
            O => \N__59326\,
            I => \N__59321\
        );

    \I__13620\ : CascadeMux
    port map (
            O => \N__59325\,
            I => \N__59318\
        );

    \I__13619\ : CascadeMux
    port map (
            O => \N__59324\,
            I => \N__59315\
        );

    \I__13618\ : Span4Mux_h
    port map (
            O => \N__59321\,
            I => \N__59312\
        );

    \I__13617\ : InMux
    port map (
            O => \N__59318\,
            I => \N__59307\
        );

    \I__13616\ : InMux
    port map (
            O => \N__59315\,
            I => \N__59307\
        );

    \I__13615\ : Odrv4
    port map (
            O => \N__59312\,
            I => \c0.data_in_frame_26_0\
        );

    \I__13614\ : LocalMux
    port map (
            O => \N__59307\,
            I => \c0.data_in_frame_26_0\
        );

    \I__13613\ : InMux
    port map (
            O => \N__59302\,
            I => \N__59297\
        );

    \I__13612\ : InMux
    port map (
            O => \N__59301\,
            I => \N__59294\
        );

    \I__13611\ : CascadeMux
    port map (
            O => \N__59300\,
            I => \N__59291\
        );

    \I__13610\ : LocalMux
    port map (
            O => \N__59297\,
            I => \N__59288\
        );

    \I__13609\ : LocalMux
    port map (
            O => \N__59294\,
            I => \N__59285\
        );

    \I__13608\ : InMux
    port map (
            O => \N__59291\,
            I => \N__59282\
        );

    \I__13607\ : Span4Mux_h
    port map (
            O => \N__59288\,
            I => \N__59279\
        );

    \I__13606\ : Span4Mux_h
    port map (
            O => \N__59285\,
            I => \N__59276\
        );

    \I__13605\ : LocalMux
    port map (
            O => \N__59282\,
            I => \N__59269\
        );

    \I__13604\ : Span4Mux_h
    port map (
            O => \N__59279\,
            I => \N__59269\
        );

    \I__13603\ : Span4Mux_h
    port map (
            O => \N__59276\,
            I => \N__59266\
        );

    \I__13602\ : InMux
    port map (
            O => \N__59275\,
            I => \N__59261\
        );

    \I__13601\ : InMux
    port map (
            O => \N__59274\,
            I => \N__59261\
        );

    \I__13600\ : Odrv4
    port map (
            O => \N__59269\,
            I => \c0.data_in_frame_27_1\
        );

    \I__13599\ : Odrv4
    port map (
            O => \N__59266\,
            I => \c0.data_in_frame_27_1\
        );

    \I__13598\ : LocalMux
    port map (
            O => \N__59261\,
            I => \c0.data_in_frame_27_1\
        );

    \I__13597\ : CascadeMux
    port map (
            O => \N__59254\,
            I => \N__59251\
        );

    \I__13596\ : InMux
    port map (
            O => \N__59251\,
            I => \N__59247\
        );

    \I__13595\ : InMux
    port map (
            O => \N__59250\,
            I => \N__59244\
        );

    \I__13594\ : LocalMux
    port map (
            O => \N__59247\,
            I => \N__59241\
        );

    \I__13593\ : LocalMux
    port map (
            O => \N__59244\,
            I => \N__59238\
        );

    \I__13592\ : Span4Mux_h
    port map (
            O => \N__59241\,
            I => \N__59232\
        );

    \I__13591\ : Span4Mux_h
    port map (
            O => \N__59238\,
            I => \N__59232\
        );

    \I__13590\ : InMux
    port map (
            O => \N__59237\,
            I => \N__59227\
        );

    \I__13589\ : Span4Mux_h
    port map (
            O => \N__59232\,
            I => \N__59224\
        );

    \I__13588\ : InMux
    port map (
            O => \N__59231\,
            I => \N__59219\
        );

    \I__13587\ : InMux
    port map (
            O => \N__59230\,
            I => \N__59219\
        );

    \I__13586\ : LocalMux
    port map (
            O => \N__59227\,
            I => \c0.data_in_frame_27_2\
        );

    \I__13585\ : Odrv4
    port map (
            O => \N__59224\,
            I => \c0.data_in_frame_27_2\
        );

    \I__13584\ : LocalMux
    port map (
            O => \N__59219\,
            I => \c0.data_in_frame_27_2\
        );

    \I__13583\ : InMux
    port map (
            O => \N__59212\,
            I => \N__59208\
        );

    \I__13582\ : CascadeMux
    port map (
            O => \N__59211\,
            I => \N__59205\
        );

    \I__13581\ : LocalMux
    port map (
            O => \N__59208\,
            I => \N__59202\
        );

    \I__13580\ : InMux
    port map (
            O => \N__59205\,
            I => \N__59199\
        );

    \I__13579\ : Span12Mux_s9_v
    port map (
            O => \N__59202\,
            I => \N__59196\
        );

    \I__13578\ : LocalMux
    port map (
            O => \N__59199\,
            I => \c0.data_in_frame_28_2\
        );

    \I__13577\ : Odrv12
    port map (
            O => \N__59196\,
            I => \c0.data_in_frame_28_2\
        );

    \I__13576\ : InMux
    port map (
            O => \N__59191\,
            I => \N__59187\
        );

    \I__13575\ : InMux
    port map (
            O => \N__59190\,
            I => \N__59184\
        );

    \I__13574\ : LocalMux
    port map (
            O => \N__59187\,
            I => \c0.n20709\
        );

    \I__13573\ : LocalMux
    port map (
            O => \N__59184\,
            I => \c0.n20709\
        );

    \I__13572\ : CascadeMux
    port map (
            O => \N__59179\,
            I => \N__59175\
        );

    \I__13571\ : InMux
    port map (
            O => \N__59178\,
            I => \N__59172\
        );

    \I__13570\ : InMux
    port map (
            O => \N__59175\,
            I => \N__59169\
        );

    \I__13569\ : LocalMux
    port map (
            O => \N__59172\,
            I => \N__59166\
        );

    \I__13568\ : LocalMux
    port map (
            O => \N__59169\,
            I => \N__59162\
        );

    \I__13567\ : Span4Mux_h
    port map (
            O => \N__59166\,
            I => \N__59159\
        );

    \I__13566\ : InMux
    port map (
            O => \N__59165\,
            I => \N__59156\
        );

    \I__13565\ : Odrv4
    port map (
            O => \N__59162\,
            I => \c0.n38_adj_3062\
        );

    \I__13564\ : Odrv4
    port map (
            O => \N__59159\,
            I => \c0.n38_adj_3062\
        );

    \I__13563\ : LocalMux
    port map (
            O => \N__59156\,
            I => \c0.n38_adj_3062\
        );

    \I__13562\ : CascadeMux
    port map (
            O => \N__59149\,
            I => \N__59146\
        );

    \I__13561\ : InMux
    port map (
            O => \N__59146\,
            I => \N__59143\
        );

    \I__13560\ : LocalMux
    port map (
            O => \N__59143\,
            I => \N__59140\
        );

    \I__13559\ : Odrv12
    port map (
            O => \N__59140\,
            I => \c0.n83_adj_3442\
        );

    \I__13558\ : CascadeMux
    port map (
            O => \N__59137\,
            I => \N__59134\
        );

    \I__13557\ : InMux
    port map (
            O => \N__59134\,
            I => \N__59130\
        );

    \I__13556\ : InMux
    port map (
            O => \N__59133\,
            I => \N__59127\
        );

    \I__13555\ : LocalMux
    port map (
            O => \N__59130\,
            I => \N__59123\
        );

    \I__13554\ : LocalMux
    port map (
            O => \N__59127\,
            I => \N__59120\
        );

    \I__13553\ : InMux
    port map (
            O => \N__59126\,
            I => \N__59117\
        );

    \I__13552\ : Span4Mux_v
    port map (
            O => \N__59123\,
            I => \N__59112\
        );

    \I__13551\ : Span4Mux_v
    port map (
            O => \N__59120\,
            I => \N__59107\
        );

    \I__13550\ : LocalMux
    port map (
            O => \N__59117\,
            I => \N__59107\
        );

    \I__13549\ : InMux
    port map (
            O => \N__59116\,
            I => \N__59104\
        );

    \I__13548\ : InMux
    port map (
            O => \N__59115\,
            I => \N__59101\
        );

    \I__13547\ : Span4Mux_h
    port map (
            O => \N__59112\,
            I => \N__59098\
        );

    \I__13546\ : Span4Mux_v
    port map (
            O => \N__59107\,
            I => \N__59095\
        );

    \I__13545\ : LocalMux
    port map (
            O => \N__59104\,
            I => data_in_frame_18_7
        );

    \I__13544\ : LocalMux
    port map (
            O => \N__59101\,
            I => data_in_frame_18_7
        );

    \I__13543\ : Odrv4
    port map (
            O => \N__59098\,
            I => data_in_frame_18_7
        );

    \I__13542\ : Odrv4
    port map (
            O => \N__59095\,
            I => data_in_frame_18_7
        );

    \I__13541\ : InMux
    port map (
            O => \N__59086\,
            I => \N__59082\
        );

    \I__13540\ : InMux
    port map (
            O => \N__59085\,
            I => \N__59079\
        );

    \I__13539\ : LocalMux
    port map (
            O => \N__59082\,
            I => \N__59076\
        );

    \I__13538\ : LocalMux
    port map (
            O => \N__59079\,
            I => \N__59069\
        );

    \I__13537\ : Span4Mux_v
    port map (
            O => \N__59076\,
            I => \N__59066\
        );

    \I__13536\ : InMux
    port map (
            O => \N__59075\,
            I => \N__59061\
        );

    \I__13535\ : InMux
    port map (
            O => \N__59074\,
            I => \N__59061\
        );

    \I__13534\ : InMux
    port map (
            O => \N__59073\,
            I => \N__59056\
        );

    \I__13533\ : InMux
    port map (
            O => \N__59072\,
            I => \N__59056\
        );

    \I__13532\ : Odrv12
    port map (
            O => \N__59069\,
            I => \c0.n12052\
        );

    \I__13531\ : Odrv4
    port map (
            O => \N__59066\,
            I => \c0.n12052\
        );

    \I__13530\ : LocalMux
    port map (
            O => \N__59061\,
            I => \c0.n12052\
        );

    \I__13529\ : LocalMux
    port map (
            O => \N__59056\,
            I => \c0.n12052\
        );

    \I__13528\ : InMux
    port map (
            O => \N__59047\,
            I => \N__59043\
        );

    \I__13527\ : InMux
    port map (
            O => \N__59046\,
            I => \N__59040\
        );

    \I__13526\ : LocalMux
    port map (
            O => \N__59043\,
            I => \N__59036\
        );

    \I__13525\ : LocalMux
    port map (
            O => \N__59040\,
            I => \N__59033\
        );

    \I__13524\ : InMux
    port map (
            O => \N__59039\,
            I => \N__59029\
        );

    \I__13523\ : Span4Mux_v
    port map (
            O => \N__59036\,
            I => \N__59024\
        );

    \I__13522\ : Span4Mux_h
    port map (
            O => \N__59033\,
            I => \N__59024\
        );

    \I__13521\ : InMux
    port map (
            O => \N__59032\,
            I => \N__59021\
        );

    \I__13520\ : LocalMux
    port map (
            O => \N__59029\,
            I => \c0.n19_adj_3056\
        );

    \I__13519\ : Odrv4
    port map (
            O => \N__59024\,
            I => \c0.n19_adj_3056\
        );

    \I__13518\ : LocalMux
    port map (
            O => \N__59021\,
            I => \c0.n19_adj_3056\
        );

    \I__13517\ : CascadeMux
    port map (
            O => \N__59014\,
            I => \c0.n19_adj_3056_cascade_\
        );

    \I__13516\ : InMux
    port map (
            O => \N__59011\,
            I => \N__59006\
        );

    \I__13515\ : InMux
    port map (
            O => \N__59010\,
            I => \N__58999\
        );

    \I__13514\ : InMux
    port map (
            O => \N__59009\,
            I => \N__58995\
        );

    \I__13513\ : LocalMux
    port map (
            O => \N__59006\,
            I => \N__58992\
        );

    \I__13512\ : InMux
    port map (
            O => \N__59005\,
            I => \N__58985\
        );

    \I__13511\ : InMux
    port map (
            O => \N__59004\,
            I => \N__58985\
        );

    \I__13510\ : InMux
    port map (
            O => \N__59003\,
            I => \N__58985\
        );

    \I__13509\ : InMux
    port map (
            O => \N__59002\,
            I => \N__58982\
        );

    \I__13508\ : LocalMux
    port map (
            O => \N__58999\,
            I => \N__58979\
        );

    \I__13507\ : InMux
    port map (
            O => \N__58998\,
            I => \N__58976\
        );

    \I__13506\ : LocalMux
    port map (
            O => \N__58995\,
            I => \N__58967\
        );

    \I__13505\ : Sp12to4
    port map (
            O => \N__58992\,
            I => \N__58967\
        );

    \I__13504\ : LocalMux
    port map (
            O => \N__58985\,
            I => \N__58967\
        );

    \I__13503\ : LocalMux
    port map (
            O => \N__58982\,
            I => \N__58967\
        );

    \I__13502\ : Span4Mux_h
    port map (
            O => \N__58979\,
            I => \N__58962\
        );

    \I__13501\ : LocalMux
    port map (
            O => \N__58976\,
            I => \N__58962\
        );

    \I__13500\ : Span12Mux_v
    port map (
            O => \N__58967\,
            I => \N__58959\
        );

    \I__13499\ : Odrv4
    port map (
            O => \N__58962\,
            I => \c0.n21045\
        );

    \I__13498\ : Odrv12
    port map (
            O => \N__58959\,
            I => \c0.n21045\
        );

    \I__13497\ : InMux
    port map (
            O => \N__58954\,
            I => \N__58951\
        );

    \I__13496\ : LocalMux
    port map (
            O => \N__58951\,
            I => \N__58948\
        );

    \I__13495\ : Span4Mux_h
    port map (
            O => \N__58948\,
            I => \N__58945\
        );

    \I__13494\ : Odrv4
    port map (
            O => \N__58945\,
            I => \c0.n29_adj_3454\
        );

    \I__13493\ : InMux
    port map (
            O => \N__58942\,
            I => \N__58937\
        );

    \I__13492\ : InMux
    port map (
            O => \N__58941\,
            I => \N__58932\
        );

    \I__13491\ : InMux
    port map (
            O => \N__58940\,
            I => \N__58932\
        );

    \I__13490\ : LocalMux
    port map (
            O => \N__58937\,
            I => \N__58926\
        );

    \I__13489\ : LocalMux
    port map (
            O => \N__58932\,
            I => \N__58926\
        );

    \I__13488\ : InMux
    port map (
            O => \N__58931\,
            I => \N__58923\
        );

    \I__13487\ : Span4Mux_v
    port map (
            O => \N__58926\,
            I => \N__58920\
        );

    \I__13486\ : LocalMux
    port map (
            O => \N__58923\,
            I => \N__58917\
        );

    \I__13485\ : Odrv4
    port map (
            O => \N__58920\,
            I => \c0.n18398\
        );

    \I__13484\ : Odrv4
    port map (
            O => \N__58917\,
            I => \c0.n18398\
        );

    \I__13483\ : InMux
    port map (
            O => \N__58912\,
            I => \N__58909\
        );

    \I__13482\ : LocalMux
    port map (
            O => \N__58909\,
            I => \N__58906\
        );

    \I__13481\ : Span4Mux_h
    port map (
            O => \N__58906\,
            I => \N__58903\
        );

    \I__13480\ : Odrv4
    port map (
            O => \N__58903\,
            I => \c0.n6_adj_3239\
        );

    \I__13479\ : InMux
    port map (
            O => \N__58900\,
            I => \N__58896\
        );

    \I__13478\ : CascadeMux
    port map (
            O => \N__58899\,
            I => \N__58892\
        );

    \I__13477\ : LocalMux
    port map (
            O => \N__58896\,
            I => \N__58889\
        );

    \I__13476\ : InMux
    port map (
            O => \N__58895\,
            I => \N__58886\
        );

    \I__13475\ : InMux
    port map (
            O => \N__58892\,
            I => \N__58883\
        );

    \I__13474\ : Span4Mux_v
    port map (
            O => \N__58889\,
            I => \N__58878\
        );

    \I__13473\ : LocalMux
    port map (
            O => \N__58886\,
            I => \N__58878\
        );

    \I__13472\ : LocalMux
    port map (
            O => \N__58883\,
            I => \N__58875\
        );

    \I__13471\ : Span4Mux_h
    port map (
            O => \N__58878\,
            I => \N__58872\
        );

    \I__13470\ : Span4Mux_v
    port map (
            O => \N__58875\,
            I => \N__58868\
        );

    \I__13469\ : Span4Mux_h
    port map (
            O => \N__58872\,
            I => \N__58865\
        );

    \I__13468\ : InMux
    port map (
            O => \N__58871\,
            I => \N__58862\
        );

    \I__13467\ : Span4Mux_h
    port map (
            O => \N__58868\,
            I => \N__58859\
        );

    \I__13466\ : Span4Mux_v
    port map (
            O => \N__58865\,
            I => \N__58856\
        );

    \I__13465\ : LocalMux
    port map (
            O => \N__58862\,
            I => data_in_frame_22_2
        );

    \I__13464\ : Odrv4
    port map (
            O => \N__58859\,
            I => data_in_frame_22_2
        );

    \I__13463\ : Odrv4
    port map (
            O => \N__58856\,
            I => data_in_frame_22_2
        );

    \I__13462\ : CascadeMux
    port map (
            O => \N__58849\,
            I => \N__58846\
        );

    \I__13461\ : InMux
    port map (
            O => \N__58846\,
            I => \N__58843\
        );

    \I__13460\ : LocalMux
    port map (
            O => \N__58843\,
            I => \c0.n19354\
        );

    \I__13459\ : InMux
    port map (
            O => \N__58840\,
            I => \N__58836\
        );

    \I__13458\ : InMux
    port map (
            O => \N__58839\,
            I => \N__58833\
        );

    \I__13457\ : LocalMux
    port map (
            O => \N__58836\,
            I => \N__58829\
        );

    \I__13456\ : LocalMux
    port map (
            O => \N__58833\,
            I => \N__58826\
        );

    \I__13455\ : InMux
    port map (
            O => \N__58832\,
            I => \N__58823\
        );

    \I__13454\ : Span4Mux_v
    port map (
            O => \N__58829\,
            I => \N__58819\
        );

    \I__13453\ : Span4Mux_v
    port map (
            O => \N__58826\,
            I => \N__58814\
        );

    \I__13452\ : LocalMux
    port map (
            O => \N__58823\,
            I => \N__58814\
        );

    \I__13451\ : InMux
    port map (
            O => \N__58822\,
            I => \N__58811\
        );

    \I__13450\ : Sp12to4
    port map (
            O => \N__58819\,
            I => \N__58808\
        );

    \I__13449\ : Span4Mux_h
    port map (
            O => \N__58814\,
            I => \N__58805\
        );

    \I__13448\ : LocalMux
    port map (
            O => \N__58811\,
            I => data_in_frame_22_7
        );

    \I__13447\ : Odrv12
    port map (
            O => \N__58808\,
            I => data_in_frame_22_7
        );

    \I__13446\ : Odrv4
    port map (
            O => \N__58805\,
            I => data_in_frame_22_7
        );

    \I__13445\ : InMux
    port map (
            O => \N__58798\,
            I => \N__58795\
        );

    \I__13444\ : LocalMux
    port map (
            O => \N__58795\,
            I => \N__58791\
        );

    \I__13443\ : InMux
    port map (
            O => \N__58794\,
            I => \N__58787\
        );

    \I__13442\ : Span4Mux_h
    port map (
            O => \N__58791\,
            I => \N__58784\
        );

    \I__13441\ : InMux
    port map (
            O => \N__58790\,
            I => \N__58781\
        );

    \I__13440\ : LocalMux
    port map (
            O => \N__58787\,
            I => \N__58778\
        );

    \I__13439\ : Span4Mux_v
    port map (
            O => \N__58784\,
            I => \N__58775\
        );

    \I__13438\ : LocalMux
    port map (
            O => \N__58781\,
            I => data_in_frame_22_3
        );

    \I__13437\ : Odrv4
    port map (
            O => \N__58778\,
            I => data_in_frame_22_3
        );

    \I__13436\ : Odrv4
    port map (
            O => \N__58775\,
            I => data_in_frame_22_3
        );

    \I__13435\ : InMux
    port map (
            O => \N__58768\,
            I => \N__58765\
        );

    \I__13434\ : LocalMux
    port map (
            O => \N__58765\,
            I => \N__58762\
        );

    \I__13433\ : Span4Mux_v
    port map (
            O => \N__58762\,
            I => \N__58757\
        );

    \I__13432\ : InMux
    port map (
            O => \N__58761\,
            I => \N__58753\
        );

    \I__13431\ : CascadeMux
    port map (
            O => \N__58760\,
            I => \N__58750\
        );

    \I__13430\ : Sp12to4
    port map (
            O => \N__58757\,
            I => \N__58747\
        );

    \I__13429\ : InMux
    port map (
            O => \N__58756\,
            I => \N__58744\
        );

    \I__13428\ : LocalMux
    port map (
            O => \N__58753\,
            I => \N__58741\
        );

    \I__13427\ : InMux
    port map (
            O => \N__58750\,
            I => \N__58738\
        );

    \I__13426\ : Span12Mux_h
    port map (
            O => \N__58747\,
            I => \N__58735\
        );

    \I__13425\ : LocalMux
    port map (
            O => \N__58744\,
            I => data_in_frame_24_0
        );

    \I__13424\ : Odrv4
    port map (
            O => \N__58741\,
            I => data_in_frame_24_0
        );

    \I__13423\ : LocalMux
    port map (
            O => \N__58738\,
            I => data_in_frame_24_0
        );

    \I__13422\ : Odrv12
    port map (
            O => \N__58735\,
            I => data_in_frame_24_0
        );

    \I__13421\ : InMux
    port map (
            O => \N__58726\,
            I => \N__58719\
        );

    \I__13420\ : InMux
    port map (
            O => \N__58725\,
            I => \N__58719\
        );

    \I__13419\ : CascadeMux
    port map (
            O => \N__58724\,
            I => \N__58716\
        );

    \I__13418\ : LocalMux
    port map (
            O => \N__58719\,
            I => \N__58712\
        );

    \I__13417\ : InMux
    port map (
            O => \N__58716\,
            I => \N__58709\
        );

    \I__13416\ : InMux
    port map (
            O => \N__58715\,
            I => \N__58705\
        );

    \I__13415\ : Span4Mux_h
    port map (
            O => \N__58712\,
            I => \N__58700\
        );

    \I__13414\ : LocalMux
    port map (
            O => \N__58709\,
            I => \N__58700\
        );

    \I__13413\ : CascadeMux
    port map (
            O => \N__58708\,
            I => \N__58697\
        );

    \I__13412\ : LocalMux
    port map (
            O => \N__58705\,
            I => \N__58694\
        );

    \I__13411\ : Span4Mux_v
    port map (
            O => \N__58700\,
            I => \N__58691\
        );

    \I__13410\ : InMux
    port map (
            O => \N__58697\,
            I => \N__58688\
        );

    \I__13409\ : Span12Mux_v
    port map (
            O => \N__58694\,
            I => \N__58685\
        );

    \I__13408\ : Sp12to4
    port map (
            O => \N__58691\,
            I => \N__58682\
        );

    \I__13407\ : LocalMux
    port map (
            O => \N__58688\,
            I => \c0.data_in_frame_26_2\
        );

    \I__13406\ : Odrv12
    port map (
            O => \N__58685\,
            I => \c0.data_in_frame_26_2\
        );

    \I__13405\ : Odrv12
    port map (
            O => \N__58682\,
            I => \c0.data_in_frame_26_2\
        );

    \I__13404\ : InMux
    port map (
            O => \N__58675\,
            I => \N__58672\
        );

    \I__13403\ : LocalMux
    port map (
            O => \N__58672\,
            I => \c0.n93_adj_3385\
        );

    \I__13402\ : InMux
    port map (
            O => \N__58669\,
            I => \N__58664\
        );

    \I__13401\ : InMux
    port map (
            O => \N__58668\,
            I => \N__58661\
        );

    \I__13400\ : InMux
    port map (
            O => \N__58667\,
            I => \N__58658\
        );

    \I__13399\ : LocalMux
    port map (
            O => \N__58664\,
            I => \N__58655\
        );

    \I__13398\ : LocalMux
    port map (
            O => \N__58661\,
            I => \N__58650\
        );

    \I__13397\ : LocalMux
    port map (
            O => \N__58658\,
            I => \N__58650\
        );

    \I__13396\ : Span4Mux_h
    port map (
            O => \N__58655\,
            I => \N__58646\
        );

    \I__13395\ : Span4Mux_h
    port map (
            O => \N__58650\,
            I => \N__58643\
        );

    \I__13394\ : InMux
    port map (
            O => \N__58649\,
            I => \N__58640\
        );

    \I__13393\ : Odrv4
    port map (
            O => \N__58646\,
            I => \c0.n32_adj_3057\
        );

    \I__13392\ : Odrv4
    port map (
            O => \N__58643\,
            I => \c0.n32_adj_3057\
        );

    \I__13391\ : LocalMux
    port map (
            O => \N__58640\,
            I => \c0.n32_adj_3057\
        );

    \I__13390\ : InMux
    port map (
            O => \N__58633\,
            I => \N__58630\
        );

    \I__13389\ : LocalMux
    port map (
            O => \N__58630\,
            I => \N__58626\
        );

    \I__13388\ : InMux
    port map (
            O => \N__58629\,
            I => \N__58623\
        );

    \I__13387\ : Span4Mux_h
    port map (
            O => \N__58626\,
            I => \N__58620\
        );

    \I__13386\ : LocalMux
    port map (
            O => \N__58623\,
            I => \N__58617\
        );

    \I__13385\ : Odrv4
    port map (
            O => \N__58620\,
            I => \c0.n62\
        );

    \I__13384\ : Odrv4
    port map (
            O => \N__58617\,
            I => \c0.n62\
        );

    \I__13383\ : InMux
    port map (
            O => \N__58612\,
            I => \N__58609\
        );

    \I__13382\ : LocalMux
    port map (
            O => \N__58609\,
            I => \c0.n68\
        );

    \I__13381\ : InMux
    port map (
            O => \N__58606\,
            I => \N__58603\
        );

    \I__13380\ : LocalMux
    port map (
            O => \N__58603\,
            I => \N__58600\
        );

    \I__13379\ : Span4Mux_v
    port map (
            O => \N__58600\,
            I => \N__58595\
        );

    \I__13378\ : InMux
    port map (
            O => \N__58599\,
            I => \N__58592\
        );

    \I__13377\ : InMux
    port map (
            O => \N__58598\,
            I => \N__58589\
        );

    \I__13376\ : Odrv4
    port map (
            O => \N__58595\,
            I => \c0.n19502\
        );

    \I__13375\ : LocalMux
    port map (
            O => \N__58592\,
            I => \c0.n19502\
        );

    \I__13374\ : LocalMux
    port map (
            O => \N__58589\,
            I => \c0.n19502\
        );

    \I__13373\ : InMux
    port map (
            O => \N__58582\,
            I => \N__58579\
        );

    \I__13372\ : LocalMux
    port map (
            O => \N__58579\,
            I => \N__58576\
        );

    \I__13371\ : Odrv12
    port map (
            O => \N__58576\,
            I => \c0.n20_adj_3536\
        );

    \I__13370\ : CascadeMux
    port map (
            O => \N__58573\,
            I => \N__58570\
        );

    \I__13369\ : InMux
    port map (
            O => \N__58570\,
            I => \N__58567\
        );

    \I__13368\ : LocalMux
    port map (
            O => \N__58567\,
            I => \N__58564\
        );

    \I__13367\ : Span4Mux_v
    port map (
            O => \N__58564\,
            I => \N__58561\
        );

    \I__13366\ : Span4Mux_h
    port map (
            O => \N__58561\,
            I => \N__58558\
        );

    \I__13365\ : Span4Mux_v
    port map (
            O => \N__58558\,
            I => \N__58555\
        );

    \I__13364\ : Odrv4
    port map (
            O => \N__58555\,
            I => \c0.n23_adj_3534\
        );

    \I__13363\ : CascadeMux
    port map (
            O => \N__58552\,
            I => \N__58547\
        );

    \I__13362\ : InMux
    port map (
            O => \N__58551\,
            I => \N__58544\
        );

    \I__13361\ : CascadeMux
    port map (
            O => \N__58550\,
            I => \N__58541\
        );

    \I__13360\ : InMux
    port map (
            O => \N__58547\,
            I => \N__58538\
        );

    \I__13359\ : LocalMux
    port map (
            O => \N__58544\,
            I => \N__58535\
        );

    \I__13358\ : InMux
    port map (
            O => \N__58541\,
            I => \N__58532\
        );

    \I__13357\ : LocalMux
    port map (
            O => \N__58538\,
            I => \N__58529\
        );

    \I__13356\ : Span4Mux_h
    port map (
            O => \N__58535\,
            I => \N__58526\
        );

    \I__13355\ : LocalMux
    port map (
            O => \N__58532\,
            I => \N__58523\
        );

    \I__13354\ : Span4Mux_v
    port map (
            O => \N__58529\,
            I => \N__58518\
        );

    \I__13353\ : Span4Mux_h
    port map (
            O => \N__58526\,
            I => \N__58518\
        );

    \I__13352\ : Span4Mux_h
    port map (
            O => \N__58523\,
            I => \N__58515\
        );

    \I__13351\ : Odrv4
    port map (
            O => \N__58518\,
            I => \c0.n40_adj_3374\
        );

    \I__13350\ : Odrv4
    port map (
            O => \N__58515\,
            I => \c0.n40_adj_3374\
        );

    \I__13349\ : CascadeMux
    port map (
            O => \N__58510\,
            I => \c0.n38_adj_3062_cascade_\
        );

    \I__13348\ : InMux
    port map (
            O => \N__58507\,
            I => \N__58503\
        );

    \I__13347\ : InMux
    port map (
            O => \N__58506\,
            I => \N__58500\
        );

    \I__13346\ : LocalMux
    port map (
            O => \N__58503\,
            I => \c0.n39_adj_3384\
        );

    \I__13345\ : LocalMux
    port map (
            O => \N__58500\,
            I => \c0.n39_adj_3384\
        );

    \I__13344\ : InMux
    port map (
            O => \N__58495\,
            I => \N__58492\
        );

    \I__13343\ : LocalMux
    port map (
            O => \N__58492\,
            I => \N__58488\
        );

    \I__13342\ : InMux
    port map (
            O => \N__58491\,
            I => \N__58485\
        );

    \I__13341\ : Span4Mux_h
    port map (
            O => \N__58488\,
            I => \N__58482\
        );

    \I__13340\ : LocalMux
    port map (
            O => \N__58485\,
            I => \N__58479\
        );

    \I__13339\ : Span4Mux_h
    port map (
            O => \N__58482\,
            I => \N__58476\
        );

    \I__13338\ : Span4Mux_h
    port map (
            O => \N__58479\,
            I => \N__58473\
        );

    \I__13337\ : Odrv4
    port map (
            O => \N__58476\,
            I => \c0.n93_adj_3329\
        );

    \I__13336\ : Odrv4
    port map (
            O => \N__58473\,
            I => \c0.n93_adj_3329\
        );

    \I__13335\ : InMux
    port map (
            O => \N__58468\,
            I => \N__58463\
        );

    \I__13334\ : CascadeMux
    port map (
            O => \N__58467\,
            I => \N__58458\
        );

    \I__13333\ : InMux
    port map (
            O => \N__58466\,
            I => \N__58455\
        );

    \I__13332\ : LocalMux
    port map (
            O => \N__58463\,
            I => \N__58452\
        );

    \I__13331\ : InMux
    port map (
            O => \N__58462\,
            I => \N__58449\
        );

    \I__13330\ : InMux
    port map (
            O => \N__58461\,
            I => \N__58446\
        );

    \I__13329\ : InMux
    port map (
            O => \N__58458\,
            I => \N__58443\
        );

    \I__13328\ : LocalMux
    port map (
            O => \N__58455\,
            I => \N__58440\
        );

    \I__13327\ : Span4Mux_v
    port map (
            O => \N__58452\,
            I => \N__58433\
        );

    \I__13326\ : LocalMux
    port map (
            O => \N__58449\,
            I => \N__58433\
        );

    \I__13325\ : LocalMux
    port map (
            O => \N__58446\,
            I => \N__58433\
        );

    \I__13324\ : LocalMux
    port map (
            O => \N__58443\,
            I => \N__58428\
        );

    \I__13323\ : Span4Mux_v
    port map (
            O => \N__58440\,
            I => \N__58423\
        );

    \I__13322\ : Span4Mux_v
    port map (
            O => \N__58433\,
            I => \N__58423\
        );

    \I__13321\ : InMux
    port map (
            O => \N__58432\,
            I => \N__58420\
        );

    \I__13320\ : InMux
    port map (
            O => \N__58431\,
            I => \N__58417\
        );

    \I__13319\ : Odrv12
    port map (
            O => \N__58428\,
            I => \c0.data_in_frame_8_3\
        );

    \I__13318\ : Odrv4
    port map (
            O => \N__58423\,
            I => \c0.data_in_frame_8_3\
        );

    \I__13317\ : LocalMux
    port map (
            O => \N__58420\,
            I => \c0.data_in_frame_8_3\
        );

    \I__13316\ : LocalMux
    port map (
            O => \N__58417\,
            I => \c0.data_in_frame_8_3\
        );

    \I__13315\ : CascadeMux
    port map (
            O => \N__58408\,
            I => \N__58405\
        );

    \I__13314\ : InMux
    port map (
            O => \N__58405\,
            I => \N__58401\
        );

    \I__13313\ : InMux
    port map (
            O => \N__58404\,
            I => \N__58398\
        );

    \I__13312\ : LocalMux
    port map (
            O => \N__58401\,
            I => \N__58395\
        );

    \I__13311\ : LocalMux
    port map (
            O => \N__58398\,
            I => \N__58392\
        );

    \I__13310\ : Span4Mux_v
    port map (
            O => \N__58395\,
            I => \N__58387\
        );

    \I__13309\ : Span4Mux_v
    port map (
            O => \N__58392\,
            I => \N__58387\
        );

    \I__13308\ : Span4Mux_h
    port map (
            O => \N__58387\,
            I => \N__58384\
        );

    \I__13307\ : Odrv4
    port map (
            O => \N__58384\,
            I => \c0.n19505\
        );

    \I__13306\ : InMux
    port map (
            O => \N__58381\,
            I => \N__58378\
        );

    \I__13305\ : LocalMux
    port map (
            O => \N__58378\,
            I => \c0.n26_adj_3537\
        );

    \I__13304\ : CascadeMux
    port map (
            O => \N__58375\,
            I => \c0.n20917_cascade_\
        );

    \I__13303\ : InMux
    port map (
            O => \N__58372\,
            I => \N__58369\
        );

    \I__13302\ : LocalMux
    port map (
            O => \N__58369\,
            I => \N__58365\
        );

    \I__13301\ : InMux
    port map (
            O => \N__58368\,
            I => \N__58362\
        );

    \I__13300\ : Span4Mux_v
    port map (
            O => \N__58365\,
            I => \N__58359\
        );

    \I__13299\ : LocalMux
    port map (
            O => \N__58362\,
            I => \N__58354\
        );

    \I__13298\ : Span4Mux_h
    port map (
            O => \N__58359\,
            I => \N__58354\
        );

    \I__13297\ : Span4Mux_v
    port map (
            O => \N__58354\,
            I => \N__58350\
        );

    \I__13296\ : InMux
    port map (
            O => \N__58353\,
            I => \N__58347\
        );

    \I__13295\ : Odrv4
    port map (
            O => \N__58350\,
            I => \c0.n19524\
        );

    \I__13294\ : LocalMux
    port map (
            O => \N__58347\,
            I => \c0.n19524\
        );

    \I__13293\ : CascadeMux
    port map (
            O => \N__58342\,
            I => \c0.n6_adj_3433_cascade_\
        );

    \I__13292\ : CascadeMux
    port map (
            O => \N__58339\,
            I => \c0.n18375_cascade_\
        );

    \I__13291\ : InMux
    port map (
            O => \N__58336\,
            I => \N__58330\
        );

    \I__13290\ : InMux
    port map (
            O => \N__58335\,
            I => \N__58330\
        );

    \I__13289\ : LocalMux
    port map (
            O => \N__58330\,
            I => \c0.n58\
        );

    \I__13288\ : CascadeMux
    port map (
            O => \N__58327\,
            I => \N__58324\
        );

    \I__13287\ : InMux
    port map (
            O => \N__58324\,
            I => \N__58321\
        );

    \I__13286\ : LocalMux
    port map (
            O => \N__58321\,
            I => \N__58318\
        );

    \I__13285\ : Span4Mux_h
    port map (
            O => \N__58318\,
            I => \N__58315\
        );

    \I__13284\ : Span4Mux_h
    port map (
            O => \N__58315\,
            I => \N__58312\
        );

    \I__13283\ : Span4Mux_v
    port map (
            O => \N__58312\,
            I => \N__58309\
        );

    \I__13282\ : Odrv4
    port map (
            O => \N__58309\,
            I => \c0.n16_adj_3489\
        );

    \I__13281\ : InMux
    port map (
            O => \N__58306\,
            I => \N__58300\
        );

    \I__13280\ : InMux
    port map (
            O => \N__58305\,
            I => \N__58300\
        );

    \I__13279\ : LocalMux
    port map (
            O => \N__58300\,
            I => \N__58297\
        );

    \I__13278\ : Span4Mux_h
    port map (
            O => \N__58297\,
            I => \N__58294\
        );

    \I__13277\ : Odrv4
    port map (
            O => \N__58294\,
            I => \c0.n31_adj_3126\
        );

    \I__13276\ : CascadeMux
    port map (
            O => \N__58291\,
            I => \c0.n10_adj_3425_cascade_\
        );

    \I__13275\ : InMux
    port map (
            O => \N__58288\,
            I => \N__58284\
        );

    \I__13274\ : InMux
    port map (
            O => \N__58287\,
            I => \N__58281\
        );

    \I__13273\ : LocalMux
    port map (
            O => \N__58284\,
            I => \c0.n42_adj_3130\
        );

    \I__13272\ : LocalMux
    port map (
            O => \N__58281\,
            I => \c0.n42_adj_3130\
        );

    \I__13271\ : InMux
    port map (
            O => \N__58276\,
            I => \N__58273\
        );

    \I__13270\ : LocalMux
    port map (
            O => \N__58273\,
            I => \N__58270\
        );

    \I__13269\ : Span4Mux_h
    port map (
            O => \N__58270\,
            I => \N__58267\
        );

    \I__13268\ : Odrv4
    port map (
            O => \N__58267\,
            I => \c0.n92_adj_3272\
        );

    \I__13267\ : InMux
    port map (
            O => \N__58264\,
            I => \N__58261\
        );

    \I__13266\ : LocalMux
    port map (
            O => \N__58261\,
            I => \c0.n39_adj_3269\
        );

    \I__13265\ : InMux
    port map (
            O => \N__58258\,
            I => \N__58255\
        );

    \I__13264\ : LocalMux
    port map (
            O => \N__58255\,
            I => \N__58252\
        );

    \I__13263\ : Span4Mux_h
    port map (
            O => \N__58252\,
            I => \N__58249\
        );

    \I__13262\ : Span4Mux_v
    port map (
            O => \N__58249\,
            I => \N__58244\
        );

    \I__13261\ : InMux
    port map (
            O => \N__58248\,
            I => \N__58239\
        );

    \I__13260\ : InMux
    port map (
            O => \N__58247\,
            I => \N__58239\
        );

    \I__13259\ : Span4Mux_h
    port map (
            O => \N__58244\,
            I => \N__58236\
        );

    \I__13258\ : LocalMux
    port map (
            O => \N__58239\,
            I => \N__58233\
        );

    \I__13257\ : Odrv4
    port map (
            O => \N__58236\,
            I => \c0.n36_adj_3275\
        );

    \I__13256\ : Odrv12
    port map (
            O => \N__58233\,
            I => \c0.n36_adj_3275\
        );

    \I__13255\ : CascadeMux
    port map (
            O => \N__58228\,
            I => \N__58224\
        );

    \I__13254\ : InMux
    port map (
            O => \N__58227\,
            I => \N__58221\
        );

    \I__13253\ : InMux
    port map (
            O => \N__58224\,
            I => \N__58218\
        );

    \I__13252\ : LocalMux
    port map (
            O => \N__58221\,
            I => \N__58212\
        );

    \I__13251\ : LocalMux
    port map (
            O => \N__58218\,
            I => \N__58212\
        );

    \I__13250\ : InMux
    port map (
            O => \N__58217\,
            I => \N__58209\
        );

    \I__13249\ : Odrv4
    port map (
            O => \N__58212\,
            I => \c0.n38_adj_3270\
        );

    \I__13248\ : LocalMux
    port map (
            O => \N__58209\,
            I => \c0.n38_adj_3270\
        );

    \I__13247\ : CascadeMux
    port map (
            O => \N__58204\,
            I => \c0.n39_adj_3269_cascade_\
        );

    \I__13246\ : InMux
    port map (
            O => \N__58201\,
            I => \N__58194\
        );

    \I__13245\ : InMux
    port map (
            O => \N__58200\,
            I => \N__58194\
        );

    \I__13244\ : InMux
    port map (
            O => \N__58199\,
            I => \N__58191\
        );

    \I__13243\ : LocalMux
    port map (
            O => \N__58194\,
            I => \c0.n37_adj_3268\
        );

    \I__13242\ : LocalMux
    port map (
            O => \N__58191\,
            I => \c0.n37_adj_3268\
        );

    \I__13241\ : InMux
    port map (
            O => \N__58186\,
            I => \N__58183\
        );

    \I__13240\ : LocalMux
    port map (
            O => \N__58183\,
            I => \N__58180\
        );

    \I__13239\ : Span4Mux_v
    port map (
            O => \N__58180\,
            I => \N__58177\
        );

    \I__13238\ : Span4Mux_h
    port map (
            O => \N__58177\,
            I => \N__58174\
        );

    \I__13237\ : Odrv4
    port map (
            O => \N__58174\,
            I => \c0.n94_adj_3375\
        );

    \I__13236\ : CascadeMux
    port map (
            O => \N__58171\,
            I => \c0.n92_adj_3377_cascade_\
        );

    \I__13235\ : InMux
    port map (
            O => \N__58168\,
            I => \N__58165\
        );

    \I__13234\ : LocalMux
    port map (
            O => \N__58165\,
            I => \N__58162\
        );

    \I__13233\ : Odrv4
    port map (
            O => \N__58162\,
            I => \c0.n91_adj_3389\
        );

    \I__13232\ : InMux
    port map (
            O => \N__58159\,
            I => \N__58156\
        );

    \I__13231\ : LocalMux
    port map (
            O => \N__58156\,
            I => \N__58153\
        );

    \I__13230\ : Odrv12
    port map (
            O => \N__58153\,
            I => \c0.n100_adj_3420\
        );

    \I__13229\ : CascadeMux
    port map (
            O => \N__58150\,
            I => \N__58147\
        );

    \I__13228\ : InMux
    port map (
            O => \N__58147\,
            I => \N__58144\
        );

    \I__13227\ : LocalMux
    port map (
            O => \N__58144\,
            I => \N__58141\
        );

    \I__13226\ : Span4Mux_h
    port map (
            O => \N__58141\,
            I => \N__58138\
        );

    \I__13225\ : Span4Mux_v
    port map (
            O => \N__58138\,
            I => \N__58135\
        );

    \I__13224\ : Span4Mux_h
    port map (
            O => \N__58135\,
            I => \N__58132\
        );

    \I__13223\ : Span4Mux_h
    port map (
            O => \N__58132\,
            I => \N__58127\
        );

    \I__13222\ : InMux
    port map (
            O => \N__58131\,
            I => \N__58124\
        );

    \I__13221\ : InMux
    port map (
            O => \N__58130\,
            I => \N__58121\
        );

    \I__13220\ : Odrv4
    port map (
            O => \N__58127\,
            I => \c0.n11942\
        );

    \I__13219\ : LocalMux
    port map (
            O => \N__58124\,
            I => \c0.n11942\
        );

    \I__13218\ : LocalMux
    port map (
            O => \N__58121\,
            I => \c0.n11942\
        );

    \I__13217\ : CascadeMux
    port map (
            O => \N__58114\,
            I => \N__58111\
        );

    \I__13216\ : InMux
    port map (
            O => \N__58111\,
            I => \N__58108\
        );

    \I__13215\ : LocalMux
    port map (
            O => \N__58108\,
            I => \N__58105\
        );

    \I__13214\ : Span4Mux_h
    port map (
            O => \N__58105\,
            I => \N__58102\
        );

    \I__13213\ : Odrv4
    port map (
            O => \N__58102\,
            I => \c0.n12_adj_3208\
        );

    \I__13212\ : InMux
    port map (
            O => \N__58099\,
            I => \N__58094\
        );

    \I__13211\ : InMux
    port map (
            O => \N__58098\,
            I => \N__58089\
        );

    \I__13210\ : InMux
    port map (
            O => \N__58097\,
            I => \N__58089\
        );

    \I__13209\ : LocalMux
    port map (
            O => \N__58094\,
            I => \c0.n10_adj_3425\
        );

    \I__13208\ : LocalMux
    port map (
            O => \N__58089\,
            I => \c0.n10_adj_3425\
        );

    \I__13207\ : InMux
    port map (
            O => \N__58084\,
            I => \N__58081\
        );

    \I__13206\ : LocalMux
    port map (
            O => \N__58081\,
            I => \N__58078\
        );

    \I__13205\ : Span4Mux_v
    port map (
            O => \N__58078\,
            I => \N__58075\
        );

    \I__13204\ : Odrv4
    port map (
            O => \N__58075\,
            I => \c0.n82\
        );

    \I__13203\ : InMux
    port map (
            O => \N__58072\,
            I => \N__58069\
        );

    \I__13202\ : LocalMux
    port map (
            O => \N__58069\,
            I => \N__58064\
        );

    \I__13201\ : InMux
    port map (
            O => \N__58068\,
            I => \N__58059\
        );

    \I__13200\ : InMux
    port map (
            O => \N__58067\,
            I => \N__58059\
        );

    \I__13199\ : Span4Mux_v
    port map (
            O => \N__58064\,
            I => \N__58054\
        );

    \I__13198\ : LocalMux
    port map (
            O => \N__58059\,
            I => \N__58054\
        );

    \I__13197\ : Span4Mux_h
    port map (
            O => \N__58054\,
            I => \N__58050\
        );

    \I__13196\ : InMux
    port map (
            O => \N__58053\,
            I => \N__58047\
        );

    \I__13195\ : Odrv4
    port map (
            O => \N__58050\,
            I => \c0.n20085\
        );

    \I__13194\ : LocalMux
    port map (
            O => \N__58047\,
            I => \c0.n20085\
        );

    \I__13193\ : InMux
    port map (
            O => \N__58042\,
            I => \N__58038\
        );

    \I__13192\ : InMux
    port map (
            O => \N__58041\,
            I => \N__58034\
        );

    \I__13191\ : LocalMux
    port map (
            O => \N__58038\,
            I => \N__58031\
        );

    \I__13190\ : InMux
    port map (
            O => \N__58037\,
            I => \N__58028\
        );

    \I__13189\ : LocalMux
    port map (
            O => \N__58034\,
            I => \N__58025\
        );

    \I__13188\ : Span4Mux_h
    port map (
            O => \N__58031\,
            I => \N__58017\
        );

    \I__13187\ : LocalMux
    port map (
            O => \N__58028\,
            I => \N__58017\
        );

    \I__13186\ : Span4Mux_v
    port map (
            O => \N__58025\,
            I => \N__58017\
        );

    \I__13185\ : InMux
    port map (
            O => \N__58024\,
            I => \N__58014\
        );

    \I__13184\ : Odrv4
    port map (
            O => \N__58017\,
            I => \c0.n19244\
        );

    \I__13183\ : LocalMux
    port map (
            O => \N__58014\,
            I => \c0.n19244\
        );

    \I__13182\ : InMux
    port map (
            O => \N__58009\,
            I => \N__58006\
        );

    \I__13181\ : LocalMux
    port map (
            O => \N__58006\,
            I => \N__58003\
        );

    \I__13180\ : Span4Mux_h
    port map (
            O => \N__58003\,
            I => \N__58000\
        );

    \I__13179\ : Span4Mux_h
    port map (
            O => \N__58000\,
            I => \N__57997\
        );

    \I__13178\ : Odrv4
    port map (
            O => \N__57997\,
            I => \c0.n88_adj_3422\
        );

    \I__13177\ : InMux
    port map (
            O => \N__57994\,
            I => \N__57991\
        );

    \I__13176\ : LocalMux
    port map (
            O => \N__57991\,
            I => \c0.n25_adj_3510\
        );

    \I__13175\ : InMux
    port map (
            O => \N__57988\,
            I => \N__57982\
        );

    \I__13174\ : InMux
    port map (
            O => \N__57987\,
            I => \N__57982\
        );

    \I__13173\ : LocalMux
    port map (
            O => \N__57982\,
            I => \N__57979\
        );

    \I__13172\ : Span4Mux_h
    port map (
            O => \N__57979\,
            I => \N__57976\
        );

    \I__13171\ : Odrv4
    port map (
            O => \N__57976\,
            I => \c0.n56\
        );

    \I__13170\ : InMux
    port map (
            O => \N__57973\,
            I => \N__57970\
        );

    \I__13169\ : LocalMux
    port map (
            O => \N__57970\,
            I => \N__57966\
        );

    \I__13168\ : InMux
    port map (
            O => \N__57969\,
            I => \N__57963\
        );

    \I__13167\ : Span4Mux_v
    port map (
            O => \N__57966\,
            I => \N__57960\
        );

    \I__13166\ : LocalMux
    port map (
            O => \N__57963\,
            I => \N__57957\
        );

    \I__13165\ : Odrv4
    port map (
            O => \N__57960\,
            I => \c0.n44_adj_3125\
        );

    \I__13164\ : Odrv4
    port map (
            O => \N__57957\,
            I => \c0.n44_adj_3125\
        );

    \I__13163\ : InMux
    port map (
            O => \N__57952\,
            I => \N__57948\
        );

    \I__13162\ : InMux
    port map (
            O => \N__57951\,
            I => \N__57945\
        );

    \I__13161\ : LocalMux
    port map (
            O => \N__57948\,
            I => \c0.n11_adj_3124\
        );

    \I__13160\ : LocalMux
    port map (
            O => \N__57945\,
            I => \c0.n11_adj_3124\
        );

    \I__13159\ : CascadeMux
    port map (
            O => \N__57940\,
            I => \N__57937\
        );

    \I__13158\ : InMux
    port map (
            O => \N__57937\,
            I => \N__57934\
        );

    \I__13157\ : LocalMux
    port map (
            O => \N__57934\,
            I => \c0.n48_adj_3313\
        );

    \I__13156\ : CascadeMux
    port map (
            O => \N__57931\,
            I => \c0.n35_cascade_\
        );

    \I__13155\ : InMux
    port map (
            O => \N__57928\,
            I => \N__57925\
        );

    \I__13154\ : LocalMux
    port map (
            O => \N__57925\,
            I => \c0.n67_adj_3092\
        );

    \I__13153\ : InMux
    port map (
            O => \N__57922\,
            I => \N__57916\
        );

    \I__13152\ : InMux
    port map (
            O => \N__57921\,
            I => \N__57916\
        );

    \I__13151\ : LocalMux
    port map (
            O => \N__57916\,
            I => \N__57913\
        );

    \I__13150\ : Odrv4
    port map (
            O => \N__57913\,
            I => \c0.n43_adj_3089\
        );

    \I__13149\ : CascadeMux
    port map (
            O => \N__57910\,
            I => \N__57906\
        );

    \I__13148\ : CascadeMux
    port map (
            O => \N__57909\,
            I => \N__57903\
        );

    \I__13147\ : InMux
    port map (
            O => \N__57906\,
            I => \N__57900\
        );

    \I__13146\ : InMux
    port map (
            O => \N__57903\,
            I => \N__57897\
        );

    \I__13145\ : LocalMux
    port map (
            O => \N__57900\,
            I => \N__57894\
        );

    \I__13144\ : LocalMux
    port map (
            O => \N__57897\,
            I => \N__57889\
        );

    \I__13143\ : Span4Mux_h
    port map (
            O => \N__57894\,
            I => \N__57889\
        );

    \I__13142\ : Span4Mux_v
    port map (
            O => \N__57889\,
            I => \N__57886\
        );

    \I__13141\ : Odrv4
    port map (
            O => \N__57886\,
            I => \c0.n41_adj_3085\
        );

    \I__13140\ : InMux
    port map (
            O => \N__57883\,
            I => \N__57879\
        );

    \I__13139\ : InMux
    port map (
            O => \N__57882\,
            I => \N__57876\
        );

    \I__13138\ : LocalMux
    port map (
            O => \N__57879\,
            I => \c0.n42_adj_3086\
        );

    \I__13137\ : LocalMux
    port map (
            O => \N__57876\,
            I => \c0.n42_adj_3086\
        );

    \I__13136\ : InMux
    port map (
            O => \N__57871\,
            I => \N__57868\
        );

    \I__13135\ : LocalMux
    port map (
            O => \N__57868\,
            I => \c0.n60_adj_3127\
        );

    \I__13134\ : CascadeMux
    port map (
            O => \N__57865\,
            I => \c0.n55_adj_3128_cascade_\
        );

    \I__13133\ : InMux
    port map (
            O => \N__57862\,
            I => \N__57859\
        );

    \I__13132\ : LocalMux
    port map (
            O => \N__57859\,
            I => \N__57854\
        );

    \I__13131\ : InMux
    port map (
            O => \N__57858\,
            I => \N__57849\
        );

    \I__13130\ : InMux
    port map (
            O => \N__57857\,
            I => \N__57849\
        );

    \I__13129\ : Span4Mux_h
    port map (
            O => \N__57854\,
            I => \N__57846\
        );

    \I__13128\ : LocalMux
    port map (
            O => \N__57849\,
            I => \N__57841\
        );

    \I__13127\ : Span4Mux_h
    port map (
            O => \N__57846\,
            I => \N__57841\
        );

    \I__13126\ : Odrv4
    port map (
            O => \N__57841\,
            I => \c0.n19749\
        );

    \I__13125\ : InMux
    port map (
            O => \N__57838\,
            I => \N__57834\
        );

    \I__13124\ : InMux
    port map (
            O => \N__57837\,
            I => \N__57831\
        );

    \I__13123\ : LocalMux
    port map (
            O => \N__57834\,
            I => \N__57828\
        );

    \I__13122\ : LocalMux
    port map (
            O => \N__57831\,
            I => \N__57825\
        );

    \I__13121\ : Odrv4
    port map (
            O => \N__57828\,
            I => \c0.n69\
        );

    \I__13120\ : Odrv4
    port map (
            O => \N__57825\,
            I => \c0.n69\
        );

    \I__13119\ : CascadeMux
    port map (
            O => \N__57820\,
            I => \N__57816\
        );

    \I__13118\ : InMux
    port map (
            O => \N__57819\,
            I => \N__57813\
        );

    \I__13117\ : InMux
    port map (
            O => \N__57816\,
            I => \N__57810\
        );

    \I__13116\ : LocalMux
    port map (
            O => \N__57813\,
            I => \N__57807\
        );

    \I__13115\ : LocalMux
    port map (
            O => \N__57810\,
            I => \c0.n28_adj_3059\
        );

    \I__13114\ : Odrv4
    port map (
            O => \N__57807\,
            I => \c0.n28_adj_3059\
        );

    \I__13113\ : CascadeMux
    port map (
            O => \N__57802\,
            I => \c0.n38_adj_3058_cascade_\
        );

    \I__13112\ : InMux
    port map (
            O => \N__57799\,
            I => \N__57796\
        );

    \I__13111\ : LocalMux
    port map (
            O => \N__57796\,
            I => \c0.n32_adj_3060\
        );

    \I__13110\ : CascadeMux
    port map (
            O => \N__57793\,
            I => \c0.n8_adj_3061_cascade_\
        );

    \I__13109\ : InMux
    port map (
            O => \N__57790\,
            I => \N__57786\
        );

    \I__13108\ : InMux
    port map (
            O => \N__57789\,
            I => \N__57783\
        );

    \I__13107\ : LocalMux
    port map (
            O => \N__57786\,
            I => \N__57778\
        );

    \I__13106\ : LocalMux
    port map (
            O => \N__57783\,
            I => \N__57778\
        );

    \I__13105\ : Span4Mux_v
    port map (
            O => \N__57778\,
            I => \N__57775\
        );

    \I__13104\ : Span4Mux_h
    port map (
            O => \N__57775\,
            I => \N__57772\
        );

    \I__13103\ : Odrv4
    port map (
            O => \N__57772\,
            I => \c0.n52\
        );

    \I__13102\ : InMux
    port map (
            O => \N__57769\,
            I => \N__57766\
        );

    \I__13101\ : LocalMux
    port map (
            O => \N__57766\,
            I => \c0.n8_adj_3061\
        );

    \I__13100\ : CascadeMux
    port map (
            O => \N__57763\,
            I => \c0.n43_adj_3285_cascade_\
        );

    \I__13099\ : InMux
    port map (
            O => \N__57760\,
            I => \N__57757\
        );

    \I__13098\ : LocalMux
    port map (
            O => \N__57757\,
            I => \c0.n53\
        );

    \I__13097\ : InMux
    port map (
            O => \N__57754\,
            I => \N__57751\
        );

    \I__13096\ : LocalMux
    port map (
            O => \N__57751\,
            I => \N__57748\
        );

    \I__13095\ : Span4Mux_h
    port map (
            O => \N__57748\,
            I => \N__57744\
        );

    \I__13094\ : InMux
    port map (
            O => \N__57747\,
            I => \N__57741\
        );

    \I__13093\ : Odrv4
    port map (
            O => \N__57744\,
            I => \c0.n4_adj_3123\
        );

    \I__13092\ : LocalMux
    port map (
            O => \N__57741\,
            I => \c0.n4_adj_3123\
        );

    \I__13091\ : InMux
    port map (
            O => \N__57736\,
            I => \N__57733\
        );

    \I__13090\ : LocalMux
    port map (
            O => \N__57733\,
            I => \N__57729\
        );

    \I__13089\ : CascadeMux
    port map (
            O => \N__57732\,
            I => \N__57726\
        );

    \I__13088\ : Span4Mux_v
    port map (
            O => \N__57729\,
            I => \N__57720\
        );

    \I__13087\ : InMux
    port map (
            O => \N__57726\,
            I => \N__57717\
        );

    \I__13086\ : InMux
    port map (
            O => \N__57725\,
            I => \N__57714\
        );

    \I__13085\ : CascadeMux
    port map (
            O => \N__57724\,
            I => \N__57710\
        );

    \I__13084\ : InMux
    port map (
            O => \N__57723\,
            I => \N__57706\
        );

    \I__13083\ : Span4Mux_h
    port map (
            O => \N__57720\,
            I => \N__57701\
        );

    \I__13082\ : LocalMux
    port map (
            O => \N__57717\,
            I => \N__57701\
        );

    \I__13081\ : LocalMux
    port map (
            O => \N__57714\,
            I => \N__57698\
        );

    \I__13080\ : InMux
    port map (
            O => \N__57713\,
            I => \N__57693\
        );

    \I__13079\ : InMux
    port map (
            O => \N__57710\,
            I => \N__57693\
        );

    \I__13078\ : InMux
    port map (
            O => \N__57709\,
            I => \N__57689\
        );

    \I__13077\ : LocalMux
    port map (
            O => \N__57706\,
            I => \N__57682\
        );

    \I__13076\ : Span4Mux_h
    port map (
            O => \N__57701\,
            I => \N__57682\
        );

    \I__13075\ : Span4Mux_h
    port map (
            O => \N__57698\,
            I => \N__57682\
        );

    \I__13074\ : LocalMux
    port map (
            O => \N__57693\,
            I => \N__57679\
        );

    \I__13073\ : InMux
    port map (
            O => \N__57692\,
            I => \N__57676\
        );

    \I__13072\ : LocalMux
    port map (
            O => \N__57689\,
            I => \N__57673\
        );

    \I__13071\ : Span4Mux_v
    port map (
            O => \N__57682\,
            I => \N__57670\
        );

    \I__13070\ : Span4Mux_v
    port map (
            O => \N__57679\,
            I => \N__57667\
        );

    \I__13069\ : LocalMux
    port map (
            O => \N__57676\,
            I => data_in_frame_16_7
        );

    \I__13068\ : Odrv12
    port map (
            O => \N__57673\,
            I => data_in_frame_16_7
        );

    \I__13067\ : Odrv4
    port map (
            O => \N__57670\,
            I => data_in_frame_16_7
        );

    \I__13066\ : Odrv4
    port map (
            O => \N__57667\,
            I => data_in_frame_16_7
        );

    \I__13065\ : InMux
    port map (
            O => \N__57658\,
            I => \N__57652\
        );

    \I__13064\ : InMux
    port map (
            O => \N__57657\,
            I => \N__57647\
        );

    \I__13063\ : InMux
    port map (
            O => \N__57656\,
            I => \N__57647\
        );

    \I__13062\ : InMux
    port map (
            O => \N__57655\,
            I => \N__57642\
        );

    \I__13061\ : LocalMux
    port map (
            O => \N__57652\,
            I => \N__57637\
        );

    \I__13060\ : LocalMux
    port map (
            O => \N__57647\,
            I => \N__57637\
        );

    \I__13059\ : InMux
    port map (
            O => \N__57646\,
            I => \N__57634\
        );

    \I__13058\ : InMux
    port map (
            O => \N__57645\,
            I => \N__57629\
        );

    \I__13057\ : LocalMux
    port map (
            O => \N__57642\,
            I => \N__57626\
        );

    \I__13056\ : Span4Mux_v
    port map (
            O => \N__57637\,
            I => \N__57623\
        );

    \I__13055\ : LocalMux
    port map (
            O => \N__57634\,
            I => \N__57620\
        );

    \I__13054\ : CascadeMux
    port map (
            O => \N__57633\,
            I => \N__57617\
        );

    \I__13053\ : InMux
    port map (
            O => \N__57632\,
            I => \N__57614\
        );

    \I__13052\ : LocalMux
    port map (
            O => \N__57629\,
            I => \N__57611\
        );

    \I__13051\ : Span4Mux_v
    port map (
            O => \N__57626\,
            I => \N__57606\
        );

    \I__13050\ : Span4Mux_v
    port map (
            O => \N__57623\,
            I => \N__57606\
        );

    \I__13049\ : Span4Mux_h
    port map (
            O => \N__57620\,
            I => \N__57603\
        );

    \I__13048\ : InMux
    port map (
            O => \N__57617\,
            I => \N__57600\
        );

    \I__13047\ : LocalMux
    port map (
            O => \N__57614\,
            I => \c0.data_in_frame_12_5\
        );

    \I__13046\ : Odrv12
    port map (
            O => \N__57611\,
            I => \c0.data_in_frame_12_5\
        );

    \I__13045\ : Odrv4
    port map (
            O => \N__57606\,
            I => \c0.data_in_frame_12_5\
        );

    \I__13044\ : Odrv4
    port map (
            O => \N__57603\,
            I => \c0.data_in_frame_12_5\
        );

    \I__13043\ : LocalMux
    port map (
            O => \N__57600\,
            I => \c0.data_in_frame_12_5\
        );

    \I__13042\ : CascadeMux
    port map (
            O => \N__57589\,
            I => \c0.n12_adj_3554_cascade_\
        );

    \I__13041\ : InMux
    port map (
            O => \N__57586\,
            I => \N__57583\
        );

    \I__13040\ : LocalMux
    port map (
            O => \N__57583\,
            I => \N__57578\
        );

    \I__13039\ : InMux
    port map (
            O => \N__57582\,
            I => \N__57573\
        );

    \I__13038\ : InMux
    port map (
            O => \N__57581\,
            I => \N__57573\
        );

    \I__13037\ : Span4Mux_v
    port map (
            O => \N__57578\,
            I => \N__57568\
        );

    \I__13036\ : LocalMux
    port map (
            O => \N__57573\,
            I => \N__57565\
        );

    \I__13035\ : InMux
    port map (
            O => \N__57572\,
            I => \N__57562\
        );

    \I__13034\ : InMux
    port map (
            O => \N__57571\,
            I => \N__57559\
        );

    \I__13033\ : Span4Mux_h
    port map (
            O => \N__57568\,
            I => \N__57552\
        );

    \I__13032\ : Span4Mux_v
    port map (
            O => \N__57565\,
            I => \N__57552\
        );

    \I__13031\ : LocalMux
    port map (
            O => \N__57562\,
            I => \N__57552\
        );

    \I__13030\ : LocalMux
    port map (
            O => \N__57559\,
            I => \c0.n20151\
        );

    \I__13029\ : Odrv4
    port map (
            O => \N__57552\,
            I => \c0.n20151\
        );

    \I__13028\ : InMux
    port map (
            O => \N__57547\,
            I => \N__57544\
        );

    \I__13027\ : LocalMux
    port map (
            O => \N__57544\,
            I => \N__57541\
        );

    \I__13026\ : Span4Mux_h
    port map (
            O => \N__57541\,
            I => \N__57538\
        );

    \I__13025\ : Odrv4
    port map (
            O => \N__57538\,
            I => \c0.n20542\
        );

    \I__13024\ : CascadeMux
    port map (
            O => \N__57535\,
            I => \c0.n20542_cascade_\
        );

    \I__13023\ : InMux
    port map (
            O => \N__57532\,
            I => \N__57529\
        );

    \I__13022\ : LocalMux
    port map (
            O => \N__57529\,
            I => \N__57526\
        );

    \I__13021\ : Span4Mux_h
    port map (
            O => \N__57526\,
            I => \N__57522\
        );

    \I__13020\ : InMux
    port map (
            O => \N__57525\,
            I => \N__57519\
        );

    \I__13019\ : Odrv4
    port map (
            O => \N__57522\,
            I => \c0.n45_adj_3423\
        );

    \I__13018\ : LocalMux
    port map (
            O => \N__57519\,
            I => \c0.n45_adj_3423\
        );

    \I__13017\ : CascadeMux
    port map (
            O => \N__57514\,
            I => \c0.n25_adj_3510_cascade_\
        );

    \I__13016\ : InMux
    port map (
            O => \N__57511\,
            I => \N__57508\
        );

    \I__13015\ : LocalMux
    port map (
            O => \N__57508\,
            I => \N__57505\
        );

    \I__13014\ : Odrv4
    port map (
            O => \N__57505\,
            I => \c0.n58_adj_3511\
        );

    \I__13013\ : InMux
    port map (
            O => \N__57502\,
            I => \N__57496\
        );

    \I__13012\ : InMux
    port map (
            O => \N__57501\,
            I => \N__57493\
        );

    \I__13011\ : CascadeMux
    port map (
            O => \N__57500\,
            I => \N__57490\
        );

    \I__13010\ : CascadeMux
    port map (
            O => \N__57499\,
            I => \N__57487\
        );

    \I__13009\ : LocalMux
    port map (
            O => \N__57496\,
            I => \N__57484\
        );

    \I__13008\ : LocalMux
    port map (
            O => \N__57493\,
            I => \N__57481\
        );

    \I__13007\ : InMux
    port map (
            O => \N__57490\,
            I => \N__57478\
        );

    \I__13006\ : InMux
    port map (
            O => \N__57487\,
            I => \N__57475\
        );

    \I__13005\ : Span4Mux_h
    port map (
            O => \N__57484\,
            I => \N__57472\
        );

    \I__13004\ : Span4Mux_v
    port map (
            O => \N__57481\,
            I => \N__57467\
        );

    \I__13003\ : LocalMux
    port map (
            O => \N__57478\,
            I => \N__57467\
        );

    \I__13002\ : LocalMux
    port map (
            O => \N__57475\,
            I => \c0.data_in_frame_14_1\
        );

    \I__13001\ : Odrv4
    port map (
            O => \N__57472\,
            I => \c0.data_in_frame_14_1\
        );

    \I__13000\ : Odrv4
    port map (
            O => \N__57467\,
            I => \c0.data_in_frame_14_1\
        );

    \I__12999\ : CascadeMux
    port map (
            O => \N__57460\,
            I => \N__57457\
        );

    \I__12998\ : InMux
    port map (
            O => \N__57457\,
            I => \N__57447\
        );

    \I__12997\ : InMux
    port map (
            O => \N__57456\,
            I => \N__57447\
        );

    \I__12996\ : InMux
    port map (
            O => \N__57455\,
            I => \N__57447\
        );

    \I__12995\ : InMux
    port map (
            O => \N__57454\,
            I => \N__57444\
        );

    \I__12994\ : LocalMux
    port map (
            O => \N__57447\,
            I => \N__57438\
        );

    \I__12993\ : LocalMux
    port map (
            O => \N__57444\,
            I => \N__57438\
        );

    \I__12992\ : InMux
    port map (
            O => \N__57443\,
            I => \N__57435\
        );

    \I__12991\ : Span4Mux_v
    port map (
            O => \N__57438\,
            I => \N__57429\
        );

    \I__12990\ : LocalMux
    port map (
            O => \N__57435\,
            I => \N__57429\
        );

    \I__12989\ : CascadeMux
    port map (
            O => \N__57434\,
            I => \N__57426\
        );

    \I__12988\ : Span4Mux_h
    port map (
            O => \N__57429\,
            I => \N__57423\
        );

    \I__12987\ : InMux
    port map (
            O => \N__57426\,
            I => \N__57420\
        );

    \I__12986\ : Span4Mux_h
    port map (
            O => \N__57423\,
            I => \N__57417\
        );

    \I__12985\ : LocalMux
    port map (
            O => \N__57420\,
            I => \c0.data_in_frame_15_7\
        );

    \I__12984\ : Odrv4
    port map (
            O => \N__57417\,
            I => \c0.data_in_frame_15_7\
        );

    \I__12983\ : InMux
    port map (
            O => \N__57412\,
            I => \N__57409\
        );

    \I__12982\ : LocalMux
    port map (
            O => \N__57409\,
            I => \N__57405\
        );

    \I__12981\ : CascadeMux
    port map (
            O => \N__57408\,
            I => \N__57402\
        );

    \I__12980\ : Span4Mux_h
    port map (
            O => \N__57405\,
            I => \N__57398\
        );

    \I__12979\ : InMux
    port map (
            O => \N__57402\,
            I => \N__57395\
        );

    \I__12978\ : InMux
    port map (
            O => \N__57401\,
            I => \N__57392\
        );

    \I__12977\ : Span4Mux_h
    port map (
            O => \N__57398\,
            I => \N__57389\
        );

    \I__12976\ : LocalMux
    port map (
            O => \N__57395\,
            I => \N__57384\
        );

    \I__12975\ : LocalMux
    port map (
            O => \N__57392\,
            I => \N__57384\
        );

    \I__12974\ : Odrv4
    port map (
            O => \N__57389\,
            I => \c0.data_in_frame_14_2\
        );

    \I__12973\ : Odrv4
    port map (
            O => \N__57384\,
            I => \c0.data_in_frame_14_2\
        );

    \I__12972\ : CascadeMux
    port map (
            O => \N__57379\,
            I => \N__57376\
        );

    \I__12971\ : InMux
    port map (
            O => \N__57376\,
            I => \N__57373\
        );

    \I__12970\ : LocalMux
    port map (
            O => \N__57373\,
            I => \N__57368\
        );

    \I__12969\ : InMux
    port map (
            O => \N__57372\,
            I => \N__57365\
        );

    \I__12968\ : InMux
    port map (
            O => \N__57371\,
            I => \N__57362\
        );

    \I__12967\ : Span4Mux_h
    port map (
            O => \N__57368\,
            I => \N__57358\
        );

    \I__12966\ : LocalMux
    port map (
            O => \N__57365\,
            I => \N__57355\
        );

    \I__12965\ : LocalMux
    port map (
            O => \N__57362\,
            I => \N__57352\
        );

    \I__12964\ : InMux
    port map (
            O => \N__57361\,
            I => \N__57349\
        );

    \I__12963\ : Span4Mux_v
    port map (
            O => \N__57358\,
            I => \N__57346\
        );

    \I__12962\ : Span4Mux_h
    port map (
            O => \N__57355\,
            I => \N__57343\
        );

    \I__12961\ : Span4Mux_h
    port map (
            O => \N__57352\,
            I => \N__57340\
        );

    \I__12960\ : LocalMux
    port map (
            O => \N__57349\,
            I => \c0.data_in_frame_7_2\
        );

    \I__12959\ : Odrv4
    port map (
            O => \N__57346\,
            I => \c0.data_in_frame_7_2\
        );

    \I__12958\ : Odrv4
    port map (
            O => \N__57343\,
            I => \c0.data_in_frame_7_2\
        );

    \I__12957\ : Odrv4
    port map (
            O => \N__57340\,
            I => \c0.data_in_frame_7_2\
        );

    \I__12956\ : InMux
    port map (
            O => \N__57331\,
            I => \N__57325\
        );

    \I__12955\ : InMux
    port map (
            O => \N__57330\,
            I => \N__57322\
        );

    \I__12954\ : InMux
    port map (
            O => \N__57329\,
            I => \N__57317\
        );

    \I__12953\ : InMux
    port map (
            O => \N__57328\,
            I => \N__57317\
        );

    \I__12952\ : LocalMux
    port map (
            O => \N__57325\,
            I => \N__57314\
        );

    \I__12951\ : LocalMux
    port map (
            O => \N__57322\,
            I => \N__57309\
        );

    \I__12950\ : LocalMux
    port map (
            O => \N__57317\,
            I => \N__57309\
        );

    \I__12949\ : Span4Mux_v
    port map (
            O => \N__57314\,
            I => \N__57302\
        );

    \I__12948\ : Span4Mux_v
    port map (
            O => \N__57309\,
            I => \N__57302\
        );

    \I__12947\ : InMux
    port map (
            O => \N__57308\,
            I => \N__57299\
        );

    \I__12946\ : InMux
    port map (
            O => \N__57307\,
            I => \N__57296\
        );

    \I__12945\ : Odrv4
    port map (
            O => \N__57302\,
            I => \c0.n20981\
        );

    \I__12944\ : LocalMux
    port map (
            O => \N__57299\,
            I => \c0.n20981\
        );

    \I__12943\ : LocalMux
    port map (
            O => \N__57296\,
            I => \c0.n20981\
        );

    \I__12942\ : InMux
    port map (
            O => \N__57289\,
            I => \N__57286\
        );

    \I__12941\ : LocalMux
    port map (
            O => \N__57286\,
            I => \N__57283\
        );

    \I__12940\ : Span4Mux_h
    port map (
            O => \N__57283\,
            I => \N__57280\
        );

    \I__12939\ : Span4Mux_v
    port map (
            O => \N__57280\,
            I => \N__57277\
        );

    \I__12938\ : Span4Mux_h
    port map (
            O => \N__57277\,
            I => \N__57274\
        );

    \I__12937\ : Odrv4
    port map (
            O => \N__57274\,
            I => \c0.n25_adj_3157\
        );

    \I__12936\ : InMux
    port map (
            O => \N__57271\,
            I => \N__57268\
        );

    \I__12935\ : LocalMux
    port map (
            O => \N__57268\,
            I => \N__57264\
        );

    \I__12934\ : InMux
    port map (
            O => \N__57267\,
            I => \N__57261\
        );

    \I__12933\ : Odrv4
    port map (
            O => \N__57264\,
            I => \c0.n5753\
        );

    \I__12932\ : LocalMux
    port map (
            O => \N__57261\,
            I => \c0.n5753\
        );

    \I__12931\ : CascadeMux
    port map (
            O => \N__57256\,
            I => \N__57252\
        );

    \I__12930\ : InMux
    port map (
            O => \N__57255\,
            I => \N__57248\
        );

    \I__12929\ : InMux
    port map (
            O => \N__57252\,
            I => \N__57245\
        );

    \I__12928\ : CascadeMux
    port map (
            O => \N__57251\,
            I => \N__57242\
        );

    \I__12927\ : LocalMux
    port map (
            O => \N__57248\,
            I => \N__57239\
        );

    \I__12926\ : LocalMux
    port map (
            O => \N__57245\,
            I => \N__57236\
        );

    \I__12925\ : InMux
    port map (
            O => \N__57242\,
            I => \N__57232\
        );

    \I__12924\ : Sp12to4
    port map (
            O => \N__57239\,
            I => \N__57229\
        );

    \I__12923\ : Span4Mux_h
    port map (
            O => \N__57236\,
            I => \N__57226\
        );

    \I__12922\ : CascadeMux
    port map (
            O => \N__57235\,
            I => \N__57222\
        );

    \I__12921\ : LocalMux
    port map (
            O => \N__57232\,
            I => \N__57219\
        );

    \I__12920\ : Span12Mux_v
    port map (
            O => \N__57229\,
            I => \N__57216\
        );

    \I__12919\ : Span4Mux_v
    port map (
            O => \N__57226\,
            I => \N__57213\
        );

    \I__12918\ : InMux
    port map (
            O => \N__57225\,
            I => \N__57208\
        );

    \I__12917\ : InMux
    port map (
            O => \N__57222\,
            I => \N__57208\
        );

    \I__12916\ : Span4Mux_h
    port map (
            O => \N__57219\,
            I => \N__57205\
        );

    \I__12915\ : Odrv12
    port map (
            O => \N__57216\,
            I => \c0.data_in_frame_14_0\
        );

    \I__12914\ : Odrv4
    port map (
            O => \N__57213\,
            I => \c0.data_in_frame_14_0\
        );

    \I__12913\ : LocalMux
    port map (
            O => \N__57208\,
            I => \c0.data_in_frame_14_0\
        );

    \I__12912\ : Odrv4
    port map (
            O => \N__57205\,
            I => \c0.data_in_frame_14_0\
        );

    \I__12911\ : InMux
    port map (
            O => \N__57196\,
            I => \N__57192\
        );

    \I__12910\ : CascadeMux
    port map (
            O => \N__57195\,
            I => \N__57188\
        );

    \I__12909\ : LocalMux
    port map (
            O => \N__57192\,
            I => \N__57184\
        );

    \I__12908\ : InMux
    port map (
            O => \N__57191\,
            I => \N__57181\
        );

    \I__12907\ : InMux
    port map (
            O => \N__57188\,
            I => \N__57178\
        );

    \I__12906\ : InMux
    port map (
            O => \N__57187\,
            I => \N__57175\
        );

    \I__12905\ : Span4Mux_v
    port map (
            O => \N__57184\,
            I => \N__57170\
        );

    \I__12904\ : LocalMux
    port map (
            O => \N__57181\,
            I => \N__57170\
        );

    \I__12903\ : LocalMux
    port map (
            O => \N__57178\,
            I => \N__57165\
        );

    \I__12902\ : LocalMux
    port map (
            O => \N__57175\,
            I => \N__57165\
        );

    \I__12901\ : Span4Mux_v
    port map (
            O => \N__57170\,
            I => \N__57162\
        );

    \I__12900\ : Odrv4
    port map (
            O => \N__57165\,
            I => \c0.data_in_frame_12_0\
        );

    \I__12899\ : Odrv4
    port map (
            O => \N__57162\,
            I => \c0.data_in_frame_12_0\
        );

    \I__12898\ : InMux
    port map (
            O => \N__57157\,
            I => \N__57154\
        );

    \I__12897\ : LocalMux
    port map (
            O => \N__57154\,
            I => \N__57149\
        );

    \I__12896\ : InMux
    port map (
            O => \N__57153\,
            I => \N__57144\
        );

    \I__12895\ : InMux
    port map (
            O => \N__57152\,
            I => \N__57144\
        );

    \I__12894\ : Span4Mux_v
    port map (
            O => \N__57149\,
            I => \N__57139\
        );

    \I__12893\ : LocalMux
    port map (
            O => \N__57144\,
            I => \N__57136\
        );

    \I__12892\ : InMux
    port map (
            O => \N__57143\,
            I => \N__57133\
        );

    \I__12891\ : InMux
    port map (
            O => \N__57142\,
            I => \N__57130\
        );

    \I__12890\ : Odrv4
    port map (
            O => \N__57139\,
            I => \c0.n20055\
        );

    \I__12889\ : Odrv4
    port map (
            O => \N__57136\,
            I => \c0.n20055\
        );

    \I__12888\ : LocalMux
    port map (
            O => \N__57133\,
            I => \c0.n20055\
        );

    \I__12887\ : LocalMux
    port map (
            O => \N__57130\,
            I => \c0.n20055\
        );

    \I__12886\ : CascadeMux
    port map (
            O => \N__57121\,
            I => \c0.n20_adj_3536_cascade_\
        );

    \I__12885\ : CascadeMux
    port map (
            O => \N__57118\,
            I => \c0.n12_adj_3558_cascade_\
        );

    \I__12884\ : InMux
    port map (
            O => \N__57115\,
            I => \N__57111\
        );

    \I__12883\ : CascadeMux
    port map (
            O => \N__57114\,
            I => \N__57108\
        );

    \I__12882\ : LocalMux
    port map (
            O => \N__57111\,
            I => \N__57104\
        );

    \I__12881\ : InMux
    port map (
            O => \N__57108\,
            I => \N__57098\
        );

    \I__12880\ : InMux
    port map (
            O => \N__57107\,
            I => \N__57098\
        );

    \I__12879\ : Span4Mux_v
    port map (
            O => \N__57104\,
            I => \N__57095\
        );

    \I__12878\ : InMux
    port map (
            O => \N__57103\,
            I => \N__57092\
        );

    \I__12877\ : LocalMux
    port map (
            O => \N__57098\,
            I => \N__57084\
        );

    \I__12876\ : Span4Mux_h
    port map (
            O => \N__57095\,
            I => \N__57084\
        );

    \I__12875\ : LocalMux
    port map (
            O => \N__57092\,
            I => \N__57084\
        );

    \I__12874\ : InMux
    port map (
            O => \N__57091\,
            I => \N__57081\
        );

    \I__12873\ : Odrv4
    port map (
            O => \N__57084\,
            I => \c0.data_in_frame_8_5\
        );

    \I__12872\ : LocalMux
    port map (
            O => \N__57081\,
            I => \c0.data_in_frame_8_5\
        );

    \I__12871\ : CascadeMux
    port map (
            O => \N__57076\,
            I => \N__57072\
        );

    \I__12870\ : InMux
    port map (
            O => \N__57075\,
            I => \N__57068\
        );

    \I__12869\ : InMux
    port map (
            O => \N__57072\,
            I => \N__57065\
        );

    \I__12868\ : InMux
    port map (
            O => \N__57071\,
            I => \N__57062\
        );

    \I__12867\ : LocalMux
    port map (
            O => \N__57068\,
            I => \N__57059\
        );

    \I__12866\ : LocalMux
    port map (
            O => \N__57065\,
            I => \N__57056\
        );

    \I__12865\ : LocalMux
    port map (
            O => \N__57062\,
            I => \N__57051\
        );

    \I__12864\ : Span4Mux_h
    port map (
            O => \N__57059\,
            I => \N__57051\
        );

    \I__12863\ : Odrv12
    port map (
            O => \N__57056\,
            I => \c0.data_in_frame_12_7\
        );

    \I__12862\ : Odrv4
    port map (
            O => \N__57051\,
            I => \c0.data_in_frame_12_7\
        );

    \I__12861\ : InMux
    port map (
            O => \N__57046\,
            I => \N__57040\
        );

    \I__12860\ : InMux
    port map (
            O => \N__57045\,
            I => \N__57037\
        );

    \I__12859\ : InMux
    port map (
            O => \N__57044\,
            I => \N__57034\
        );

    \I__12858\ : InMux
    port map (
            O => \N__57043\,
            I => \N__57031\
        );

    \I__12857\ : LocalMux
    port map (
            O => \N__57040\,
            I => \N__57028\
        );

    \I__12856\ : LocalMux
    port map (
            O => \N__57037\,
            I => \N__57025\
        );

    \I__12855\ : LocalMux
    port map (
            O => \N__57034\,
            I => \N__57021\
        );

    \I__12854\ : LocalMux
    port map (
            O => \N__57031\,
            I => \N__57018\
        );

    \I__12853\ : Span4Mux_h
    port map (
            O => \N__57028\,
            I => \N__57013\
        );

    \I__12852\ : Span4Mux_h
    port map (
            O => \N__57025\,
            I => \N__57013\
        );

    \I__12851\ : InMux
    port map (
            O => \N__57024\,
            I => \N__57010\
        );

    \I__12850\ : Span4Mux_h
    port map (
            O => \N__57021\,
            I => \N__57007\
        );

    \I__12849\ : Span4Mux_h
    port map (
            O => \N__57018\,
            I => \N__57001\
        );

    \I__12848\ : Span4Mux_v
    port map (
            O => \N__57013\,
            I => \N__56998\
        );

    \I__12847\ : LocalMux
    port map (
            O => \N__57010\,
            I => \N__56993\
        );

    \I__12846\ : Sp12to4
    port map (
            O => \N__57007\,
            I => \N__56993\
        );

    \I__12845\ : InMux
    port map (
            O => \N__57006\,
            I => \N__56988\
        );

    \I__12844\ : InMux
    port map (
            O => \N__57005\,
            I => \N__56988\
        );

    \I__12843\ : InMux
    port map (
            O => \N__57004\,
            I => \N__56985\
        );

    \I__12842\ : Odrv4
    port map (
            O => \N__57001\,
            I => \c0.n5_adj_3031\
        );

    \I__12841\ : Odrv4
    port map (
            O => \N__56998\,
            I => \c0.n5_adj_3031\
        );

    \I__12840\ : Odrv12
    port map (
            O => \N__56993\,
            I => \c0.n5_adj_3031\
        );

    \I__12839\ : LocalMux
    port map (
            O => \N__56988\,
            I => \c0.n5_adj_3031\
        );

    \I__12838\ : LocalMux
    port map (
            O => \N__56985\,
            I => \c0.n5_adj_3031\
        );

    \I__12837\ : CascadeMux
    port map (
            O => \N__56974\,
            I => \c0.n19359_cascade_\
        );

    \I__12836\ : CascadeMux
    port map (
            O => \N__56971\,
            I => \N__56967\
        );

    \I__12835\ : InMux
    port map (
            O => \N__56970\,
            I => \N__56964\
        );

    \I__12834\ : InMux
    port map (
            O => \N__56967\,
            I => \N__56961\
        );

    \I__12833\ : LocalMux
    port map (
            O => \N__56964\,
            I => \N__56958\
        );

    \I__12832\ : LocalMux
    port map (
            O => \N__56961\,
            I => \N__56954\
        );

    \I__12831\ : Span4Mux_h
    port map (
            O => \N__56958\,
            I => \N__56951\
        );

    \I__12830\ : InMux
    port map (
            O => \N__56957\,
            I => \N__56948\
        );

    \I__12829\ : Odrv4
    port map (
            O => \N__56954\,
            I => \c0.data_in_frame_8_4\
        );

    \I__12828\ : Odrv4
    port map (
            O => \N__56951\,
            I => \c0.data_in_frame_8_4\
        );

    \I__12827\ : LocalMux
    port map (
            O => \N__56948\,
            I => \c0.data_in_frame_8_4\
        );

    \I__12826\ : InMux
    port map (
            O => \N__56941\,
            I => \N__56933\
        );

    \I__12825\ : InMux
    port map (
            O => \N__56940\,
            I => \N__56933\
        );

    \I__12824\ : InMux
    port map (
            O => \N__56939\,
            I => \N__56930\
        );

    \I__12823\ : InMux
    port map (
            O => \N__56938\,
            I => \N__56927\
        );

    \I__12822\ : LocalMux
    port map (
            O => \N__56933\,
            I => \N__56922\
        );

    \I__12821\ : LocalMux
    port map (
            O => \N__56930\,
            I => \N__56922\
        );

    \I__12820\ : LocalMux
    port map (
            O => \N__56927\,
            I => \c0.n11478\
        );

    \I__12819\ : Odrv12
    port map (
            O => \N__56922\,
            I => \c0.n11478\
        );

    \I__12818\ : InMux
    port map (
            O => \N__56917\,
            I => \N__56914\
        );

    \I__12817\ : LocalMux
    port map (
            O => \N__56914\,
            I => \c0.n19199\
        );

    \I__12816\ : InMux
    port map (
            O => \N__56911\,
            I => \N__56908\
        );

    \I__12815\ : LocalMux
    port map (
            O => \N__56908\,
            I => \N__56905\
        );

    \I__12814\ : Span4Mux_h
    port map (
            O => \N__56905\,
            I => \N__56899\
        );

    \I__12813\ : InMux
    port map (
            O => \N__56904\,
            I => \N__56896\
        );

    \I__12812\ : InMux
    port map (
            O => \N__56903\,
            I => \N__56891\
        );

    \I__12811\ : InMux
    port map (
            O => \N__56902\,
            I => \N__56891\
        );

    \I__12810\ : Span4Mux_h
    port map (
            O => \N__56899\,
            I => \N__56888\
        );

    \I__12809\ : LocalMux
    port map (
            O => \N__56896\,
            I => \c0.data_in_frame_10_5\
        );

    \I__12808\ : LocalMux
    port map (
            O => \N__56891\,
            I => \c0.data_in_frame_10_5\
        );

    \I__12807\ : Odrv4
    port map (
            O => \N__56888\,
            I => \c0.data_in_frame_10_5\
        );

    \I__12806\ : CascadeMux
    port map (
            O => \N__56881\,
            I => \c0.n19199_cascade_\
        );

    \I__12805\ : CascadeMux
    port map (
            O => \N__56878\,
            I => \N__56875\
        );

    \I__12804\ : InMux
    port map (
            O => \N__56875\,
            I => \N__56872\
        );

    \I__12803\ : LocalMux
    port map (
            O => \N__56872\,
            I => \N__56869\
        );

    \I__12802\ : Span4Mux_h
    port map (
            O => \N__56869\,
            I => \N__56866\
        );

    \I__12801\ : Span4Mux_h
    port map (
            O => \N__56866\,
            I => \N__56863\
        );

    \I__12800\ : Odrv4
    port map (
            O => \N__56863\,
            I => \c0.n19_adj_3540\
        );

    \I__12799\ : CascadeMux
    port map (
            O => \N__56860\,
            I => \N__56857\
        );

    \I__12798\ : InMux
    port map (
            O => \N__56857\,
            I => \N__56854\
        );

    \I__12797\ : LocalMux
    port map (
            O => \N__56854\,
            I => \N__56849\
        );

    \I__12796\ : InMux
    port map (
            O => \N__56853\,
            I => \N__56843\
        );

    \I__12795\ : InMux
    port map (
            O => \N__56852\,
            I => \N__56840\
        );

    \I__12794\ : Span4Mux_h
    port map (
            O => \N__56849\,
            I => \N__56837\
        );

    \I__12793\ : InMux
    port map (
            O => \N__56848\,
            I => \N__56834\
        );

    \I__12792\ : InMux
    port map (
            O => \N__56847\,
            I => \N__56831\
        );

    \I__12791\ : InMux
    port map (
            O => \N__56846\,
            I => \N__56826\
        );

    \I__12790\ : LocalMux
    port map (
            O => \N__56843\,
            I => \N__56818\
        );

    \I__12789\ : LocalMux
    port map (
            O => \N__56840\,
            I => \N__56818\
        );

    \I__12788\ : Span4Mux_h
    port map (
            O => \N__56837\,
            I => \N__56811\
        );

    \I__12787\ : LocalMux
    port map (
            O => \N__56834\,
            I => \N__56811\
        );

    \I__12786\ : LocalMux
    port map (
            O => \N__56831\,
            I => \N__56811\
        );

    \I__12785\ : CascadeMux
    port map (
            O => \N__56830\,
            I => \N__56807\
        );

    \I__12784\ : CascadeMux
    port map (
            O => \N__56829\,
            I => \N__56804\
        );

    \I__12783\ : LocalMux
    port map (
            O => \N__56826\,
            I => \N__56797\
        );

    \I__12782\ : InMux
    port map (
            O => \N__56825\,
            I => \N__56794\
        );

    \I__12781\ : InMux
    port map (
            O => \N__56824\,
            I => \N__56791\
        );

    \I__12780\ : InMux
    port map (
            O => \N__56823\,
            I => \N__56788\
        );

    \I__12779\ : Span4Mux_h
    port map (
            O => \N__56818\,
            I => \N__56783\
        );

    \I__12778\ : Span4Mux_h
    port map (
            O => \N__56811\,
            I => \N__56783\
        );

    \I__12777\ : InMux
    port map (
            O => \N__56810\,
            I => \N__56776\
        );

    \I__12776\ : InMux
    port map (
            O => \N__56807\,
            I => \N__56776\
        );

    \I__12775\ : InMux
    port map (
            O => \N__56804\,
            I => \N__56776\
        );

    \I__12774\ : InMux
    port map (
            O => \N__56803\,
            I => \N__56771\
        );

    \I__12773\ : InMux
    port map (
            O => \N__56802\,
            I => \N__56771\
        );

    \I__12772\ : InMux
    port map (
            O => \N__56801\,
            I => \N__56768\
        );

    \I__12771\ : InMux
    port map (
            O => \N__56800\,
            I => \N__56765\
        );

    \I__12770\ : Span4Mux_h
    port map (
            O => \N__56797\,
            I => \N__56758\
        );

    \I__12769\ : LocalMux
    port map (
            O => \N__56794\,
            I => \N__56758\
        );

    \I__12768\ : LocalMux
    port map (
            O => \N__56791\,
            I => \N__56758\
        );

    \I__12767\ : LocalMux
    port map (
            O => \N__56788\,
            I => data_in_frame_0_1
        );

    \I__12766\ : Odrv4
    port map (
            O => \N__56783\,
            I => data_in_frame_0_1
        );

    \I__12765\ : LocalMux
    port map (
            O => \N__56776\,
            I => data_in_frame_0_1
        );

    \I__12764\ : LocalMux
    port map (
            O => \N__56771\,
            I => data_in_frame_0_1
        );

    \I__12763\ : LocalMux
    port map (
            O => \N__56768\,
            I => data_in_frame_0_1
        );

    \I__12762\ : LocalMux
    port map (
            O => \N__56765\,
            I => data_in_frame_0_1
        );

    \I__12761\ : Odrv4
    port map (
            O => \N__56758\,
            I => data_in_frame_0_1
        );

    \I__12760\ : InMux
    port map (
            O => \N__56743\,
            I => \N__56740\
        );

    \I__12759\ : LocalMux
    port map (
            O => \N__56740\,
            I => \N__56737\
        );

    \I__12758\ : Span4Mux_h
    port map (
            O => \N__56737\,
            I => \N__56734\
        );

    \I__12757\ : Odrv4
    port map (
            O => \N__56734\,
            I => \c0.n17_adj_3544\
        );

    \I__12756\ : CascadeMux
    port map (
            O => \N__56731\,
            I => \N__56728\
        );

    \I__12755\ : InMux
    port map (
            O => \N__56728\,
            I => \N__56723\
        );

    \I__12754\ : InMux
    port map (
            O => \N__56727\,
            I => \N__56720\
        );

    \I__12753\ : InMux
    port map (
            O => \N__56726\,
            I => \N__56716\
        );

    \I__12752\ : LocalMux
    port map (
            O => \N__56723\,
            I => \N__56711\
        );

    \I__12751\ : LocalMux
    port map (
            O => \N__56720\,
            I => \N__56711\
        );

    \I__12750\ : InMux
    port map (
            O => \N__56719\,
            I => \N__56708\
        );

    \I__12749\ : LocalMux
    port map (
            O => \N__56716\,
            I => \N__56704\
        );

    \I__12748\ : Span4Mux_h
    port map (
            O => \N__56711\,
            I => \N__56700\
        );

    \I__12747\ : LocalMux
    port map (
            O => \N__56708\,
            I => \N__56697\
        );

    \I__12746\ : InMux
    port map (
            O => \N__56707\,
            I => \N__56694\
        );

    \I__12745\ : Span4Mux_h
    port map (
            O => \N__56704\,
            I => \N__56691\
        );

    \I__12744\ : InMux
    port map (
            O => \N__56703\,
            I => \N__56688\
        );

    \I__12743\ : Span4Mux_h
    port map (
            O => \N__56700\,
            I => \N__56685\
        );

    \I__12742\ : Span4Mux_h
    port map (
            O => \N__56697\,
            I => \N__56682\
        );

    \I__12741\ : LocalMux
    port map (
            O => \N__56694\,
            I => \c0.data_in_frame_9_1\
        );

    \I__12740\ : Odrv4
    port map (
            O => \N__56691\,
            I => \c0.data_in_frame_9_1\
        );

    \I__12739\ : LocalMux
    port map (
            O => \N__56688\,
            I => \c0.data_in_frame_9_1\
        );

    \I__12738\ : Odrv4
    port map (
            O => \N__56685\,
            I => \c0.data_in_frame_9_1\
        );

    \I__12737\ : Odrv4
    port map (
            O => \N__56682\,
            I => \c0.data_in_frame_9_1\
        );

    \I__12736\ : CascadeMux
    port map (
            O => \N__56671\,
            I => \c0.n11858_cascade_\
        );

    \I__12735\ : InMux
    port map (
            O => \N__56668\,
            I => \N__56665\
        );

    \I__12734\ : LocalMux
    port map (
            O => \N__56665\,
            I => \N__56662\
        );

    \I__12733\ : Span4Mux_v
    port map (
            O => \N__56662\,
            I => \N__56659\
        );

    \I__12732\ : Odrv4
    port map (
            O => \N__56659\,
            I => \c0.n19446\
        );

    \I__12731\ : CascadeMux
    port map (
            O => \N__56656\,
            I => \c0.n19446_cascade_\
        );

    \I__12730\ : InMux
    port map (
            O => \N__56653\,
            I => \N__56647\
        );

    \I__12729\ : InMux
    port map (
            O => \N__56652\,
            I => \N__56643\
        );

    \I__12728\ : InMux
    port map (
            O => \N__56651\,
            I => \N__56637\
        );

    \I__12727\ : InMux
    port map (
            O => \N__56650\,
            I => \N__56637\
        );

    \I__12726\ : LocalMux
    port map (
            O => \N__56647\,
            I => \N__56634\
        );

    \I__12725\ : InMux
    port map (
            O => \N__56646\,
            I => \N__56631\
        );

    \I__12724\ : LocalMux
    port map (
            O => \N__56643\,
            I => \N__56626\
        );

    \I__12723\ : InMux
    port map (
            O => \N__56642\,
            I => \N__56623\
        );

    \I__12722\ : LocalMux
    port map (
            O => \N__56637\,
            I => \N__56620\
        );

    \I__12721\ : Span4Mux_v
    port map (
            O => \N__56634\,
            I => \N__56617\
        );

    \I__12720\ : LocalMux
    port map (
            O => \N__56631\,
            I => \N__56614\
        );

    \I__12719\ : InMux
    port map (
            O => \N__56630\,
            I => \N__56611\
        );

    \I__12718\ : InMux
    port map (
            O => \N__56629\,
            I => \N__56608\
        );

    \I__12717\ : Span4Mux_v
    port map (
            O => \N__56626\,
            I => \N__56605\
        );

    \I__12716\ : LocalMux
    port map (
            O => \N__56623\,
            I => \N__56602\
        );

    \I__12715\ : Span4Mux_v
    port map (
            O => \N__56620\,
            I => \N__56599\
        );

    \I__12714\ : Span4Mux_h
    port map (
            O => \N__56617\,
            I => \N__56594\
        );

    \I__12713\ : Span4Mux_v
    port map (
            O => \N__56614\,
            I => \N__56594\
        );

    \I__12712\ : LocalMux
    port map (
            O => \N__56611\,
            I => \N__56591\
        );

    \I__12711\ : LocalMux
    port map (
            O => \N__56608\,
            I => \c0.data_out_frame_0__7__N_1537\
        );

    \I__12710\ : Odrv4
    port map (
            O => \N__56605\,
            I => \c0.data_out_frame_0__7__N_1537\
        );

    \I__12709\ : Odrv4
    port map (
            O => \N__56602\,
            I => \c0.data_out_frame_0__7__N_1537\
        );

    \I__12708\ : Odrv4
    port map (
            O => \N__56599\,
            I => \c0.data_out_frame_0__7__N_1537\
        );

    \I__12707\ : Odrv4
    port map (
            O => \N__56594\,
            I => \c0.data_out_frame_0__7__N_1537\
        );

    \I__12706\ : Odrv12
    port map (
            O => \N__56591\,
            I => \c0.data_out_frame_0__7__N_1537\
        );

    \I__12705\ : InMux
    port map (
            O => \N__56578\,
            I => \N__56575\
        );

    \I__12704\ : LocalMux
    port map (
            O => \N__56575\,
            I => \N__56572\
        );

    \I__12703\ : Odrv12
    port map (
            O => \N__56572\,
            I => \c0.n11982\
        );

    \I__12702\ : CascadeMux
    port map (
            O => \N__56569\,
            I => \c0.n33_adj_3209_cascade_\
        );

    \I__12701\ : InMux
    port map (
            O => \N__56566\,
            I => \N__56563\
        );

    \I__12700\ : LocalMux
    port map (
            O => \N__56563\,
            I => \N__56557\
        );

    \I__12699\ : InMux
    port map (
            O => \N__56562\,
            I => \N__56552\
        );

    \I__12698\ : InMux
    port map (
            O => \N__56561\,
            I => \N__56552\
        );

    \I__12697\ : InMux
    port map (
            O => \N__56560\,
            I => \N__56549\
        );

    \I__12696\ : Span4Mux_v
    port map (
            O => \N__56557\,
            I => \N__56546\
        );

    \I__12695\ : LocalMux
    port map (
            O => \N__56552\,
            I => \N__56543\
        );

    \I__12694\ : LocalMux
    port map (
            O => \N__56549\,
            I => \N__56540\
        );

    \I__12693\ : Odrv4
    port map (
            O => \N__56546\,
            I => \c0.n5598\
        );

    \I__12692\ : Odrv4
    port map (
            O => \N__56543\,
            I => \c0.n5598\
        );

    \I__12691\ : Odrv4
    port map (
            O => \N__56540\,
            I => \c0.n5598\
        );

    \I__12690\ : CascadeMux
    port map (
            O => \N__56533\,
            I => \N__56530\
        );

    \I__12689\ : InMux
    port map (
            O => \N__56530\,
            I => \N__56525\
        );

    \I__12688\ : InMux
    port map (
            O => \N__56529\,
            I => \N__56521\
        );

    \I__12687\ : InMux
    port map (
            O => \N__56528\,
            I => \N__56518\
        );

    \I__12686\ : LocalMux
    port map (
            O => \N__56525\,
            I => \N__56515\
        );

    \I__12685\ : CascadeMux
    port map (
            O => \N__56524\,
            I => \N__56512\
        );

    \I__12684\ : LocalMux
    port map (
            O => \N__56521\,
            I => \N__56509\
        );

    \I__12683\ : LocalMux
    port map (
            O => \N__56518\,
            I => \N__56504\
        );

    \I__12682\ : Span4Mux_h
    port map (
            O => \N__56515\,
            I => \N__56504\
        );

    \I__12681\ : InMux
    port map (
            O => \N__56512\,
            I => \N__56501\
        );

    \I__12680\ : Span12Mux_h
    port map (
            O => \N__56509\,
            I => \N__56498\
        );

    \I__12679\ : Span4Mux_v
    port map (
            O => \N__56504\,
            I => \N__56495\
        );

    \I__12678\ : LocalMux
    port map (
            O => \N__56501\,
            I => \c0.data_in_frame_17_7\
        );

    \I__12677\ : Odrv12
    port map (
            O => \N__56498\,
            I => \c0.data_in_frame_17_7\
        );

    \I__12676\ : Odrv4
    port map (
            O => \N__56495\,
            I => \c0.data_in_frame_17_7\
        );

    \I__12675\ : InMux
    port map (
            O => \N__56488\,
            I => \N__56485\
        );

    \I__12674\ : LocalMux
    port map (
            O => \N__56485\,
            I => \N__56481\
        );

    \I__12673\ : InMux
    port map (
            O => \N__56484\,
            I => \N__56478\
        );

    \I__12672\ : Span4Mux_v
    port map (
            O => \N__56481\,
            I => \N__56475\
        );

    \I__12671\ : LocalMux
    port map (
            O => \N__56478\,
            I => \c0.n9_adj_3350\
        );

    \I__12670\ : Odrv4
    port map (
            O => \N__56475\,
            I => \c0.n9_adj_3350\
        );

    \I__12669\ : InMux
    port map (
            O => \N__56470\,
            I => \N__56467\
        );

    \I__12668\ : LocalMux
    port map (
            O => \N__56467\,
            I => \N__56464\
        );

    \I__12667\ : Span4Mux_v
    port map (
            O => \N__56464\,
            I => \N__56461\
        );

    \I__12666\ : Odrv4
    port map (
            O => \N__56461\,
            I => \c0.n29_adj_3533\
        );

    \I__12665\ : InMux
    port map (
            O => \N__56458\,
            I => \N__56455\
        );

    \I__12664\ : LocalMux
    port map (
            O => \N__56455\,
            I => \c0.n33_adj_3209\
        );

    \I__12663\ : CascadeMux
    port map (
            O => \N__56452\,
            I => \N__56447\
        );

    \I__12662\ : InMux
    port map (
            O => \N__56451\,
            I => \N__56442\
        );

    \I__12661\ : InMux
    port map (
            O => \N__56450\,
            I => \N__56442\
        );

    \I__12660\ : InMux
    port map (
            O => \N__56447\,
            I => \N__56437\
        );

    \I__12659\ : LocalMux
    port map (
            O => \N__56442\,
            I => \N__56434\
        );

    \I__12658\ : InMux
    port map (
            O => \N__56441\,
            I => \N__56429\
        );

    \I__12657\ : InMux
    port map (
            O => \N__56440\,
            I => \N__56429\
        );

    \I__12656\ : LocalMux
    port map (
            O => \N__56437\,
            I => \N__56426\
        );

    \I__12655\ : Span4Mux_h
    port map (
            O => \N__56434\,
            I => \N__56421\
        );

    \I__12654\ : LocalMux
    port map (
            O => \N__56429\,
            I => \N__56421\
        );

    \I__12653\ : Span4Mux_v
    port map (
            O => \N__56426\,
            I => \N__56418\
        );

    \I__12652\ : Span4Mux_v
    port map (
            O => \N__56421\,
            I => \N__56413\
        );

    \I__12651\ : Span4Mux_h
    port map (
            O => \N__56418\,
            I => \N__56413\
        );

    \I__12650\ : Odrv4
    port map (
            O => \N__56413\,
            I => \c0.n12209\
        );

    \I__12649\ : InMux
    port map (
            O => \N__56410\,
            I => \N__56406\
        );

    \I__12648\ : InMux
    port map (
            O => \N__56409\,
            I => \N__56403\
        );

    \I__12647\ : LocalMux
    port map (
            O => \N__56406\,
            I => \N__56400\
        );

    \I__12646\ : LocalMux
    port map (
            O => \N__56403\,
            I => \N__56393\
        );

    \I__12645\ : Span4Mux_h
    port map (
            O => \N__56400\,
            I => \N__56393\
        );

    \I__12644\ : InMux
    port map (
            O => \N__56399\,
            I => \N__56390\
        );

    \I__12643\ : InMux
    port map (
            O => \N__56398\,
            I => \N__56387\
        );

    \I__12642\ : Span4Mux_v
    port map (
            O => \N__56393\,
            I => \N__56384\
        );

    \I__12641\ : LocalMux
    port map (
            O => \N__56390\,
            I => \N__56379\
        );

    \I__12640\ : LocalMux
    port map (
            O => \N__56387\,
            I => \N__56379\
        );

    \I__12639\ : Span4Mux_v
    port map (
            O => \N__56384\,
            I => \N__56373\
        );

    \I__12638\ : Span4Mux_v
    port map (
            O => \N__56379\,
            I => \N__56373\
        );

    \I__12637\ : InMux
    port map (
            O => \N__56378\,
            I => \N__56370\
        );

    \I__12636\ : Odrv4
    port map (
            O => \N__56373\,
            I => \c0.n9_adj_3027\
        );

    \I__12635\ : LocalMux
    port map (
            O => \N__56370\,
            I => \c0.n9_adj_3027\
        );

    \I__12634\ : InMux
    port map (
            O => \N__56365\,
            I => \N__56362\
        );

    \I__12633\ : LocalMux
    port map (
            O => \N__56362\,
            I => \c0.n45_adj_3224\
        );

    \I__12632\ : CascadeMux
    port map (
            O => \N__56359\,
            I => \N__56356\
        );

    \I__12631\ : InMux
    port map (
            O => \N__56356\,
            I => \N__56353\
        );

    \I__12630\ : LocalMux
    port map (
            O => \N__56353\,
            I => \N__56348\
        );

    \I__12629\ : InMux
    port map (
            O => \N__56352\,
            I => \N__56345\
        );

    \I__12628\ : CascadeMux
    port map (
            O => \N__56351\,
            I => \N__56342\
        );

    \I__12627\ : Span4Mux_h
    port map (
            O => \N__56348\,
            I => \N__56338\
        );

    \I__12626\ : LocalMux
    port map (
            O => \N__56345\,
            I => \N__56335\
        );

    \I__12625\ : InMux
    port map (
            O => \N__56342\,
            I => \N__56332\
        );

    \I__12624\ : InMux
    port map (
            O => \N__56341\,
            I => \N__56329\
        );

    \I__12623\ : Span4Mux_h
    port map (
            O => \N__56338\,
            I => \N__56326\
        );

    \I__12622\ : Span4Mux_h
    port map (
            O => \N__56335\,
            I => \N__56323\
        );

    \I__12621\ : LocalMux
    port map (
            O => \N__56332\,
            I => \c0.data_in_frame_7_6\
        );

    \I__12620\ : LocalMux
    port map (
            O => \N__56329\,
            I => \c0.data_in_frame_7_6\
        );

    \I__12619\ : Odrv4
    port map (
            O => \N__56326\,
            I => \c0.data_in_frame_7_6\
        );

    \I__12618\ : Odrv4
    port map (
            O => \N__56323\,
            I => \c0.data_in_frame_7_6\
        );

    \I__12617\ : InMux
    port map (
            O => \N__56314\,
            I => \N__56308\
        );

    \I__12616\ : InMux
    port map (
            O => \N__56313\,
            I => \N__56308\
        );

    \I__12615\ : LocalMux
    port map (
            O => \N__56308\,
            I => \N__56305\
        );

    \I__12614\ : Sp12to4
    port map (
            O => \N__56305\,
            I => \N__56302\
        );

    \I__12613\ : Odrv12
    port map (
            O => \N__56302\,
            I => \c0.n15\
        );

    \I__12612\ : InMux
    port map (
            O => \N__56299\,
            I => \N__56296\
        );

    \I__12611\ : LocalMux
    port map (
            O => \N__56296\,
            I => \N__56292\
        );

    \I__12610\ : InMux
    port map (
            O => \N__56295\,
            I => \N__56287\
        );

    \I__12609\ : Span4Mux_h
    port map (
            O => \N__56292\,
            I => \N__56284\
        );

    \I__12608\ : InMux
    port map (
            O => \N__56291\,
            I => \N__56279\
        );

    \I__12607\ : InMux
    port map (
            O => \N__56290\,
            I => \N__56279\
        );

    \I__12606\ : LocalMux
    port map (
            O => \N__56287\,
            I => \c0.n23\
        );

    \I__12605\ : Odrv4
    port map (
            O => \N__56284\,
            I => \c0.n23\
        );

    \I__12604\ : LocalMux
    port map (
            O => \N__56279\,
            I => \c0.n23\
        );

    \I__12603\ : InMux
    port map (
            O => \N__56272\,
            I => \N__56269\
        );

    \I__12602\ : LocalMux
    port map (
            O => \N__56269\,
            I => \c0.n51_adj_3426\
        );

    \I__12601\ : InMux
    port map (
            O => \N__56266\,
            I => \N__56263\
        );

    \I__12600\ : LocalMux
    port map (
            O => \N__56263\,
            I => \N__56260\
        );

    \I__12599\ : Span4Mux_v
    port map (
            O => \N__56260\,
            I => \N__56256\
        );

    \I__12598\ : InMux
    port map (
            O => \N__56259\,
            I => \N__56253\
        );

    \I__12597\ : Span4Mux_h
    port map (
            O => \N__56256\,
            I => \N__56248\
        );

    \I__12596\ : LocalMux
    port map (
            O => \N__56253\,
            I => \N__56248\
        );

    \I__12595\ : Span4Mux_h
    port map (
            O => \N__56248\,
            I => \N__56245\
        );

    \I__12594\ : Span4Mux_v
    port map (
            O => \N__56245\,
            I => \N__56242\
        );

    \I__12593\ : Odrv4
    port map (
            O => \N__56242\,
            I => n15645
        );

    \I__12592\ : CascadeMux
    port map (
            O => \N__56239\,
            I => \N__56233\
        );

    \I__12591\ : CascadeMux
    port map (
            O => \N__56238\,
            I => \N__56230\
        );

    \I__12590\ : CascadeMux
    port map (
            O => \N__56237\,
            I => \N__56227\
        );

    \I__12589\ : CascadeMux
    port map (
            O => \N__56236\,
            I => \N__56221\
        );

    \I__12588\ : InMux
    port map (
            O => \N__56233\,
            I => \N__56214\
        );

    \I__12587\ : InMux
    port map (
            O => \N__56230\,
            I => \N__56214\
        );

    \I__12586\ : InMux
    port map (
            O => \N__56227\,
            I => \N__56214\
        );

    \I__12585\ : CascadeMux
    port map (
            O => \N__56226\,
            I => \N__56210\
        );

    \I__12584\ : CascadeMux
    port map (
            O => \N__56225\,
            I => \N__56207\
        );

    \I__12583\ : CascadeMux
    port map (
            O => \N__56224\,
            I => \N__56204\
        );

    \I__12582\ : InMux
    port map (
            O => \N__56221\,
            I => \N__56201\
        );

    \I__12581\ : LocalMux
    port map (
            O => \N__56214\,
            I => \N__56197\
        );

    \I__12580\ : InMux
    port map (
            O => \N__56213\,
            I => \N__56194\
        );

    \I__12579\ : InMux
    port map (
            O => \N__56210\,
            I => \N__56188\
        );

    \I__12578\ : InMux
    port map (
            O => \N__56207\,
            I => \N__56188\
        );

    \I__12577\ : InMux
    port map (
            O => \N__56204\,
            I => \N__56185\
        );

    \I__12576\ : LocalMux
    port map (
            O => \N__56201\,
            I => \N__56182\
        );

    \I__12575\ : InMux
    port map (
            O => \N__56200\,
            I => \N__56179\
        );

    \I__12574\ : Span4Mux_h
    port map (
            O => \N__56197\,
            I => \N__56176\
        );

    \I__12573\ : LocalMux
    port map (
            O => \N__56194\,
            I => \N__56173\
        );

    \I__12572\ : InMux
    port map (
            O => \N__56193\,
            I => \N__56170\
        );

    \I__12571\ : LocalMux
    port map (
            O => \N__56188\,
            I => \N__56167\
        );

    \I__12570\ : LocalMux
    port map (
            O => \N__56185\,
            I => \N__56164\
        );

    \I__12569\ : Sp12to4
    port map (
            O => \N__56182\,
            I => \N__56161\
        );

    \I__12568\ : LocalMux
    port map (
            O => \N__56179\,
            I => \N__56158\
        );

    \I__12567\ : Span4Mux_v
    port map (
            O => \N__56176\,
            I => \N__56155\
        );

    \I__12566\ : Span4Mux_h
    port map (
            O => \N__56173\,
            I => \N__56149\
        );

    \I__12565\ : LocalMux
    port map (
            O => \N__56170\,
            I => \N__56149\
        );

    \I__12564\ : Span4Mux_v
    port map (
            O => \N__56167\,
            I => \N__56146\
        );

    \I__12563\ : Span4Mux_v
    port map (
            O => \N__56164\,
            I => \N__56143\
        );

    \I__12562\ : Span12Mux_s10_v
    port map (
            O => \N__56161\,
            I => \N__56140\
        );

    \I__12561\ : Span4Mux_v
    port map (
            O => \N__56158\,
            I => \N__56135\
        );

    \I__12560\ : Span4Mux_v
    port map (
            O => \N__56155\,
            I => \N__56135\
        );

    \I__12559\ : InMux
    port map (
            O => \N__56154\,
            I => \N__56132\
        );

    \I__12558\ : Span4Mux_v
    port map (
            O => \N__56149\,
            I => \N__56127\
        );

    \I__12557\ : Span4Mux_h
    port map (
            O => \N__56146\,
            I => \N__56127\
        );

    \I__12556\ : Sp12to4
    port map (
            O => \N__56143\,
            I => \N__56123\
        );

    \I__12555\ : Span12Mux_h
    port map (
            O => \N__56140\,
            I => \N__56120\
        );

    \I__12554\ : Span4Mux_h
    port map (
            O => \N__56135\,
            I => \N__56117\
        );

    \I__12553\ : LocalMux
    port map (
            O => \N__56132\,
            I => \N__56114\
        );

    \I__12552\ : Sp12to4
    port map (
            O => \N__56127\,
            I => \N__56111\
        );

    \I__12551\ : InMux
    port map (
            O => \N__56126\,
            I => \N__56108\
        );

    \I__12550\ : Span12Mux_s9_v
    port map (
            O => \N__56123\,
            I => \N__56103\
        );

    \I__12549\ : Span12Mux_v
    port map (
            O => \N__56120\,
            I => \N__56103\
        );

    \I__12548\ : Span4Mux_v
    port map (
            O => \N__56117\,
            I => \N__56098\
        );

    \I__12547\ : Span4Mux_h
    port map (
            O => \N__56114\,
            I => \N__56098\
        );

    \I__12546\ : Span12Mux_h
    port map (
            O => \N__56111\,
            I => \N__56093\
        );

    \I__12545\ : LocalMux
    port map (
            O => \N__56108\,
            I => \N__56093\
        );

    \I__12544\ : Odrv12
    port map (
            O => \N__56103\,
            I => \r_Rx_Data\
        );

    \I__12543\ : Odrv4
    port map (
            O => \N__56098\,
            I => \r_Rx_Data\
        );

    \I__12542\ : Odrv12
    port map (
            O => \N__56093\,
            I => \r_Rx_Data\
        );

    \I__12541\ : InMux
    port map (
            O => \N__56086\,
            I => \N__56081\
        );

    \I__12540\ : InMux
    port map (
            O => \N__56085\,
            I => \N__56077\
        );

    \I__12539\ : InMux
    port map (
            O => \N__56084\,
            I => \N__56074\
        );

    \I__12538\ : LocalMux
    port map (
            O => \N__56081\,
            I => \N__56071\
        );

    \I__12537\ : CascadeMux
    port map (
            O => \N__56080\,
            I => \N__56068\
        );

    \I__12536\ : LocalMux
    port map (
            O => \N__56077\,
            I => \N__56065\
        );

    \I__12535\ : LocalMux
    port map (
            O => \N__56074\,
            I => \N__56062\
        );

    \I__12534\ : Span4Mux_h
    port map (
            O => \N__56071\,
            I => \N__56059\
        );

    \I__12533\ : InMux
    port map (
            O => \N__56068\,
            I => \N__56056\
        );

    \I__12532\ : Span4Mux_v
    port map (
            O => \N__56065\,
            I => \N__56053\
        );

    \I__12531\ : Span4Mux_h
    port map (
            O => \N__56062\,
            I => \N__56048\
        );

    \I__12530\ : Span4Mux_h
    port map (
            O => \N__56059\,
            I => \N__56048\
        );

    \I__12529\ : LocalMux
    port map (
            O => \N__56056\,
            I => \N__56043\
        );

    \I__12528\ : Span4Mux_h
    port map (
            O => \N__56053\,
            I => \N__56043\
        );

    \I__12527\ : Span4Mux_v
    port map (
            O => \N__56048\,
            I => \N__56040\
        );

    \I__12526\ : Span4Mux_h
    port map (
            O => \N__56043\,
            I => \N__56035\
        );

    \I__12525\ : Span4Mux_v
    port map (
            O => \N__56040\,
            I => \N__56035\
        );

    \I__12524\ : Odrv4
    port map (
            O => \N__56035\,
            I => n11466
        );

    \I__12523\ : InMux
    port map (
            O => \N__56032\,
            I => \N__56029\
        );

    \I__12522\ : LocalMux
    port map (
            O => \N__56029\,
            I => \N__56024\
        );

    \I__12521\ : InMux
    port map (
            O => \N__56028\,
            I => \N__56021\
        );

    \I__12520\ : InMux
    port map (
            O => \N__56027\,
            I => \N__56018\
        );

    \I__12519\ : Span4Mux_v
    port map (
            O => \N__56024\,
            I => \N__56014\
        );

    \I__12518\ : LocalMux
    port map (
            O => \N__56021\,
            I => \N__56011\
        );

    \I__12517\ : LocalMux
    port map (
            O => \N__56018\,
            I => \N__56008\
        );

    \I__12516\ : CascadeMux
    port map (
            O => \N__56017\,
            I => \N__56005\
        );

    \I__12515\ : Span4Mux_v
    port map (
            O => \N__56014\,
            I => \N__56002\
        );

    \I__12514\ : Span4Mux_h
    port map (
            O => \N__56011\,
            I => \N__55999\
        );

    \I__12513\ : Span4Mux_h
    port map (
            O => \N__56008\,
            I => \N__55996\
        );

    \I__12512\ : InMux
    port map (
            O => \N__56005\,
            I => \N__55993\
        );

    \I__12511\ : Span4Mux_h
    port map (
            O => \N__56002\,
            I => \N__55988\
        );

    \I__12510\ : Span4Mux_v
    port map (
            O => \N__55999\,
            I => \N__55988\
        );

    \I__12509\ : Span4Mux_h
    port map (
            O => \N__55996\,
            I => \N__55985\
        );

    \I__12508\ : LocalMux
    port map (
            O => \N__55993\,
            I => \c0.data_in_frame_13_7\
        );

    \I__12507\ : Odrv4
    port map (
            O => \N__55988\,
            I => \c0.data_in_frame_13_7\
        );

    \I__12506\ : Odrv4
    port map (
            O => \N__55985\,
            I => \c0.data_in_frame_13_7\
        );

    \I__12505\ : CascadeMux
    port map (
            O => \N__55978\,
            I => \N__55975\
        );

    \I__12504\ : InMux
    port map (
            O => \N__55975\,
            I => \N__55972\
        );

    \I__12503\ : LocalMux
    port map (
            O => \N__55972\,
            I => \N__55969\
        );

    \I__12502\ : Span4Mux_v
    port map (
            O => \N__55969\,
            I => \N__55966\
        );

    \I__12501\ : Span4Mux_v
    port map (
            O => \N__55966\,
            I => \N__55963\
        );

    \I__12500\ : Odrv4
    port map (
            O => \N__55963\,
            I => \c0.n13_adj_3541\
        );

    \I__12499\ : InMux
    port map (
            O => \N__55960\,
            I => \N__55956\
        );

    \I__12498\ : CascadeMux
    port map (
            O => \N__55959\,
            I => \N__55953\
        );

    \I__12497\ : LocalMux
    port map (
            O => \N__55956\,
            I => \N__55948\
        );

    \I__12496\ : InMux
    port map (
            O => \N__55953\,
            I => \N__55945\
        );

    \I__12495\ : InMux
    port map (
            O => \N__55952\,
            I => \N__55942\
        );

    \I__12494\ : CascadeMux
    port map (
            O => \N__55951\,
            I => \N__55939\
        );

    \I__12493\ : Span4Mux_v
    port map (
            O => \N__55948\,
            I => \N__55932\
        );

    \I__12492\ : LocalMux
    port map (
            O => \N__55945\,
            I => \N__55932\
        );

    \I__12491\ : LocalMux
    port map (
            O => \N__55942\,
            I => \N__55932\
        );

    \I__12490\ : InMux
    port map (
            O => \N__55939\,
            I => \N__55929\
        );

    \I__12489\ : Span4Mux_v
    port map (
            O => \N__55932\,
            I => \N__55926\
        );

    \I__12488\ : LocalMux
    port map (
            O => \N__55929\,
            I => \c0.data_in_frame_13_2\
        );

    \I__12487\ : Odrv4
    port map (
            O => \N__55926\,
            I => \c0.data_in_frame_13_2\
        );

    \I__12486\ : InMux
    port map (
            O => \N__55921\,
            I => \N__55916\
        );

    \I__12485\ : CascadeMux
    port map (
            O => \N__55920\,
            I => \N__55913\
        );

    \I__12484\ : InMux
    port map (
            O => \N__55919\,
            I => \N__55910\
        );

    \I__12483\ : LocalMux
    port map (
            O => \N__55916\,
            I => \N__55907\
        );

    \I__12482\ : InMux
    port map (
            O => \N__55913\,
            I => \N__55904\
        );

    \I__12481\ : LocalMux
    port map (
            O => \N__55910\,
            I => \N__55901\
        );

    \I__12480\ : Span4Mux_h
    port map (
            O => \N__55907\,
            I => \N__55898\
        );

    \I__12479\ : LocalMux
    port map (
            O => \N__55904\,
            I => \N__55893\
        );

    \I__12478\ : Span4Mux_v
    port map (
            O => \N__55901\,
            I => \N__55893\
        );

    \I__12477\ : Odrv4
    port map (
            O => \N__55898\,
            I => \c0.data_in_frame_9_5\
        );

    \I__12476\ : Odrv4
    port map (
            O => \N__55893\,
            I => \c0.data_in_frame_9_5\
        );

    \I__12475\ : InMux
    port map (
            O => \N__55888\,
            I => \N__55880\
        );

    \I__12474\ : InMux
    port map (
            O => \N__55887\,
            I => \N__55877\
        );

    \I__12473\ : CascadeMux
    port map (
            O => \N__55886\,
            I => \N__55869\
        );

    \I__12472\ : InMux
    port map (
            O => \N__55885\,
            I => \N__55862\
        );

    \I__12471\ : InMux
    port map (
            O => \N__55884\,
            I => \N__55862\
        );

    \I__12470\ : InMux
    port map (
            O => \N__55883\,
            I => \N__55859\
        );

    \I__12469\ : LocalMux
    port map (
            O => \N__55880\,
            I => \N__55854\
        );

    \I__12468\ : LocalMux
    port map (
            O => \N__55877\,
            I => \N__55854\
        );

    \I__12467\ : InMux
    port map (
            O => \N__55876\,
            I => \N__55849\
        );

    \I__12466\ : InMux
    port map (
            O => \N__55875\,
            I => \N__55849\
        );

    \I__12465\ : InMux
    port map (
            O => \N__55874\,
            I => \N__55842\
        );

    \I__12464\ : InMux
    port map (
            O => \N__55873\,
            I => \N__55842\
        );

    \I__12463\ : InMux
    port map (
            O => \N__55872\,
            I => \N__55842\
        );

    \I__12462\ : InMux
    port map (
            O => \N__55869\,
            I => \N__55839\
        );

    \I__12461\ : CascadeMux
    port map (
            O => \N__55868\,
            I => \N__55836\
        );

    \I__12460\ : InMux
    port map (
            O => \N__55867\,
            I => \N__55833\
        );

    \I__12459\ : LocalMux
    port map (
            O => \N__55862\,
            I => \N__55828\
        );

    \I__12458\ : LocalMux
    port map (
            O => \N__55859\,
            I => \N__55828\
        );

    \I__12457\ : Span4Mux_h
    port map (
            O => \N__55854\,
            I => \N__55825\
        );

    \I__12456\ : LocalMux
    port map (
            O => \N__55849\,
            I => \N__55820\
        );

    \I__12455\ : LocalMux
    port map (
            O => \N__55842\,
            I => \N__55820\
        );

    \I__12454\ : LocalMux
    port map (
            O => \N__55839\,
            I => \N__55816\
        );

    \I__12453\ : InMux
    port map (
            O => \N__55836\,
            I => \N__55813\
        );

    \I__12452\ : LocalMux
    port map (
            O => \N__55833\,
            I => \N__55809\
        );

    \I__12451\ : Span4Mux_v
    port map (
            O => \N__55828\,
            I => \N__55806\
        );

    \I__12450\ : Span4Mux_h
    port map (
            O => \N__55825\,
            I => \N__55801\
        );

    \I__12449\ : Span4Mux_v
    port map (
            O => \N__55820\,
            I => \N__55801\
        );

    \I__12448\ : CascadeMux
    port map (
            O => \N__55819\,
            I => \N__55797\
        );

    \I__12447\ : Span4Mux_v
    port map (
            O => \N__55816\,
            I => \N__55792\
        );

    \I__12446\ : LocalMux
    port map (
            O => \N__55813\,
            I => \N__55789\
        );

    \I__12445\ : InMux
    port map (
            O => \N__55812\,
            I => \N__55786\
        );

    \I__12444\ : Span4Mux_h
    port map (
            O => \N__55809\,
            I => \N__55783\
        );

    \I__12443\ : Span4Mux_h
    port map (
            O => \N__55806\,
            I => \N__55778\
        );

    \I__12442\ : Span4Mux_v
    port map (
            O => \N__55801\,
            I => \N__55778\
        );

    \I__12441\ : InMux
    port map (
            O => \N__55800\,
            I => \N__55775\
        );

    \I__12440\ : InMux
    port map (
            O => \N__55797\,
            I => \N__55768\
        );

    \I__12439\ : InMux
    port map (
            O => \N__55796\,
            I => \N__55768\
        );

    \I__12438\ : InMux
    port map (
            O => \N__55795\,
            I => \N__55768\
        );

    \I__12437\ : Span4Mux_v
    port map (
            O => \N__55792\,
            I => \N__55765\
        );

    \I__12436\ : Span4Mux_v
    port map (
            O => \N__55789\,
            I => \N__55762\
        );

    \I__12435\ : LocalMux
    port map (
            O => \N__55786\,
            I => \N__55757\
        );

    \I__12434\ : Span4Mux_v
    port map (
            O => \N__55783\,
            I => \N__55757\
        );

    \I__12433\ : Span4Mux_h
    port map (
            O => \N__55778\,
            I => \N__55754\
        );

    \I__12432\ : LocalMux
    port map (
            O => \N__55775\,
            I => \N__55747\
        );

    \I__12431\ : LocalMux
    port map (
            O => \N__55768\,
            I => \N__55747\
        );

    \I__12430\ : Sp12to4
    port map (
            O => \N__55765\,
            I => \N__55747\
        );

    \I__12429\ : Span4Mux_h
    port map (
            O => \N__55762\,
            I => \N__55742\
        );

    \I__12428\ : Span4Mux_v
    port map (
            O => \N__55757\,
            I => \N__55742\
        );

    \I__12427\ : Sp12to4
    port map (
            O => \N__55754\,
            I => \N__55737\
        );

    \I__12426\ : Span12Mux_v
    port map (
            O => \N__55747\,
            I => \N__55737\
        );

    \I__12425\ : Odrv4
    port map (
            O => \N__55742\,
            I => \c0.n9_adj_3211\
        );

    \I__12424\ : Odrv12
    port map (
            O => \N__55737\,
            I => \c0.n9_adj_3211\
        );

    \I__12423\ : InMux
    port map (
            O => \N__55732\,
            I => \N__55729\
        );

    \I__12422\ : LocalMux
    port map (
            O => \N__55729\,
            I => \N__55726\
        );

    \I__12421\ : Span4Mux_h
    port map (
            O => \N__55726\,
            I => \N__55721\
        );

    \I__12420\ : InMux
    port map (
            O => \N__55725\,
            I => \N__55718\
        );

    \I__12419\ : InMux
    port map (
            O => \N__55724\,
            I => \N__55715\
        );

    \I__12418\ : Odrv4
    port map (
            O => \N__55721\,
            I => \c0.n6_adj_3019\
        );

    \I__12417\ : LocalMux
    port map (
            O => \N__55718\,
            I => \c0.n6_adj_3019\
        );

    \I__12416\ : LocalMux
    port map (
            O => \N__55715\,
            I => \c0.n6_adj_3019\
        );

    \I__12415\ : CascadeMux
    port map (
            O => \N__55708\,
            I => \N__55705\
        );

    \I__12414\ : InMux
    port map (
            O => \N__55705\,
            I => \N__55701\
        );

    \I__12413\ : InMux
    port map (
            O => \N__55704\,
            I => \N__55698\
        );

    \I__12412\ : LocalMux
    port map (
            O => \N__55701\,
            I => \N__55693\
        );

    \I__12411\ : LocalMux
    port map (
            O => \N__55698\,
            I => \N__55690\
        );

    \I__12410\ : InMux
    port map (
            O => \N__55697\,
            I => \N__55685\
        );

    \I__12409\ : InMux
    port map (
            O => \N__55696\,
            I => \N__55685\
        );

    \I__12408\ : Odrv4
    port map (
            O => \N__55693\,
            I => \c0.data_in_frame_7_5\
        );

    \I__12407\ : Odrv4
    port map (
            O => \N__55690\,
            I => \c0.data_in_frame_7_5\
        );

    \I__12406\ : LocalMux
    port map (
            O => \N__55685\,
            I => \c0.data_in_frame_7_5\
        );

    \I__12405\ : CascadeMux
    port map (
            O => \N__55678\,
            I => \c0.n6_adj_3019_cascade_\
        );

    \I__12404\ : CascadeMux
    port map (
            O => \N__55675\,
            I => \N__55672\
        );

    \I__12403\ : InMux
    port map (
            O => \N__55672\,
            I => \N__55665\
        );

    \I__12402\ : CascadeMux
    port map (
            O => \N__55671\,
            I => \N__55662\
        );

    \I__12401\ : InMux
    port map (
            O => \N__55670\,
            I => \N__55659\
        );

    \I__12400\ : InMux
    port map (
            O => \N__55669\,
            I => \N__55656\
        );

    \I__12399\ : InMux
    port map (
            O => \N__55668\,
            I => \N__55653\
        );

    \I__12398\ : LocalMux
    port map (
            O => \N__55665\,
            I => \N__55650\
        );

    \I__12397\ : InMux
    port map (
            O => \N__55662\,
            I => \N__55647\
        );

    \I__12396\ : LocalMux
    port map (
            O => \N__55659\,
            I => \N__55642\
        );

    \I__12395\ : LocalMux
    port map (
            O => \N__55656\,
            I => \N__55642\
        );

    \I__12394\ : LocalMux
    port map (
            O => \N__55653\,
            I => \N__55639\
        );

    \I__12393\ : Span4Mux_v
    port map (
            O => \N__55650\,
            I => \N__55636\
        );

    \I__12392\ : LocalMux
    port map (
            O => \N__55647\,
            I => \N__55631\
        );

    \I__12391\ : Span4Mux_v
    port map (
            O => \N__55642\,
            I => \N__55631\
        );

    \I__12390\ : Span12Mux_h
    port map (
            O => \N__55639\,
            I => \N__55628\
        );

    \I__12389\ : Span4Mux_v
    port map (
            O => \N__55636\,
            I => \N__55623\
        );

    \I__12388\ : Span4Mux_h
    port map (
            O => \N__55631\,
            I => \N__55623\
        );

    \I__12387\ : Odrv12
    port map (
            O => \N__55628\,
            I => \c0.n20386\
        );

    \I__12386\ : Odrv4
    port map (
            O => \N__55623\,
            I => \c0.n20386\
        );

    \I__12385\ : InMux
    port map (
            O => \N__55618\,
            I => \N__55615\
        );

    \I__12384\ : LocalMux
    port map (
            O => \N__55615\,
            I => \N__55611\
        );

    \I__12383\ : CascadeMux
    port map (
            O => \N__55614\,
            I => \N__55607\
        );

    \I__12382\ : Span4Mux_h
    port map (
            O => \N__55611\,
            I => \N__55604\
        );

    \I__12381\ : InMux
    port map (
            O => \N__55610\,
            I => \N__55601\
        );

    \I__12380\ : InMux
    port map (
            O => \N__55607\,
            I => \N__55598\
        );

    \I__12379\ : Span4Mux_v
    port map (
            O => \N__55604\,
            I => \N__55593\
        );

    \I__12378\ : LocalMux
    port map (
            O => \N__55601\,
            I => \N__55593\
        );

    \I__12377\ : LocalMux
    port map (
            O => \N__55598\,
            I => \c0.data_in_frame_9_6\
        );

    \I__12376\ : Odrv4
    port map (
            O => \N__55593\,
            I => \c0.data_in_frame_9_6\
        );

    \I__12375\ : InMux
    port map (
            O => \N__55588\,
            I => \N__55580\
        );

    \I__12374\ : InMux
    port map (
            O => \N__55587\,
            I => \N__55575\
        );

    \I__12373\ : InMux
    port map (
            O => \N__55586\,
            I => \N__55575\
        );

    \I__12372\ : InMux
    port map (
            O => \N__55585\,
            I => \N__55572\
        );

    \I__12371\ : InMux
    port map (
            O => \N__55584\,
            I => \N__55569\
        );

    \I__12370\ : InMux
    port map (
            O => \N__55583\,
            I => \N__55566\
        );

    \I__12369\ : LocalMux
    port map (
            O => \N__55580\,
            I => \N__55559\
        );

    \I__12368\ : LocalMux
    port map (
            O => \N__55575\,
            I => \N__55559\
        );

    \I__12367\ : LocalMux
    port map (
            O => \N__55572\,
            I => \N__55559\
        );

    \I__12366\ : LocalMux
    port map (
            O => \N__55569\,
            I => \N__55556\
        );

    \I__12365\ : LocalMux
    port map (
            O => \N__55566\,
            I => \c0.data_in_frame_3_7\
        );

    \I__12364\ : Odrv12
    port map (
            O => \N__55559\,
            I => \c0.data_in_frame_3_7\
        );

    \I__12363\ : Odrv4
    port map (
            O => \N__55556\,
            I => \c0.data_in_frame_3_7\
        );

    \I__12362\ : InMux
    port map (
            O => \N__55549\,
            I => \N__55545\
        );

    \I__12361\ : CascadeMux
    port map (
            O => \N__55548\,
            I => \N__55541\
        );

    \I__12360\ : LocalMux
    port map (
            O => \N__55545\,
            I => \N__55537\
        );

    \I__12359\ : InMux
    port map (
            O => \N__55544\,
            I => \N__55532\
        );

    \I__12358\ : InMux
    port map (
            O => \N__55541\,
            I => \N__55532\
        );

    \I__12357\ : InMux
    port map (
            O => \N__55540\,
            I => \N__55529\
        );

    \I__12356\ : Span12Mux_h
    port map (
            O => \N__55537\,
            I => \N__55526\
        );

    \I__12355\ : LocalMux
    port map (
            O => \N__55532\,
            I => \N__55523\
        );

    \I__12354\ : LocalMux
    port map (
            O => \N__55529\,
            I => \c0.data_in_frame_5_5\
        );

    \I__12353\ : Odrv12
    port map (
            O => \N__55526\,
            I => \c0.data_in_frame_5_5\
        );

    \I__12352\ : Odrv4
    port map (
            O => \N__55523\,
            I => \c0.data_in_frame_5_5\
        );

    \I__12351\ : InMux
    port map (
            O => \N__55516\,
            I => \N__55512\
        );

    \I__12350\ : CascadeMux
    port map (
            O => \N__55515\,
            I => \N__55506\
        );

    \I__12349\ : LocalMux
    port map (
            O => \N__55512\,
            I => \N__55502\
        );

    \I__12348\ : InMux
    port map (
            O => \N__55511\,
            I => \N__55499\
        );

    \I__12347\ : InMux
    port map (
            O => \N__55510\,
            I => \N__55496\
        );

    \I__12346\ : InMux
    port map (
            O => \N__55509\,
            I => \N__55493\
        );

    \I__12345\ : InMux
    port map (
            O => \N__55506\,
            I => \N__55490\
        );

    \I__12344\ : InMux
    port map (
            O => \N__55505\,
            I => \N__55487\
        );

    \I__12343\ : Span4Mux_h
    port map (
            O => \N__55502\,
            I => \N__55484\
        );

    \I__12342\ : LocalMux
    port map (
            O => \N__55499\,
            I => \N__55477\
        );

    \I__12341\ : LocalMux
    port map (
            O => \N__55496\,
            I => \N__55477\
        );

    \I__12340\ : LocalMux
    port map (
            O => \N__55493\,
            I => \N__55477\
        );

    \I__12339\ : LocalMux
    port map (
            O => \N__55490\,
            I => \c0.data_in_frame_5_3\
        );

    \I__12338\ : LocalMux
    port map (
            O => \N__55487\,
            I => \c0.data_in_frame_5_3\
        );

    \I__12337\ : Odrv4
    port map (
            O => \N__55484\,
            I => \c0.data_in_frame_5_3\
        );

    \I__12336\ : Odrv12
    port map (
            O => \N__55477\,
            I => \c0.data_in_frame_5_3\
        );

    \I__12335\ : InMux
    port map (
            O => \N__55468\,
            I => \N__55462\
        );

    \I__12334\ : InMux
    port map (
            O => \N__55467\,
            I => \N__55459\
        );

    \I__12333\ : InMux
    port map (
            O => \N__55466\,
            I => \N__55454\
        );

    \I__12332\ : InMux
    port map (
            O => \N__55465\,
            I => \N__55454\
        );

    \I__12331\ : LocalMux
    port map (
            O => \N__55462\,
            I => \N__55451\
        );

    \I__12330\ : LocalMux
    port map (
            O => \N__55459\,
            I => \N__55448\
        );

    \I__12329\ : LocalMux
    port map (
            O => \N__55454\,
            I => \N__55445\
        );

    \I__12328\ : Span4Mux_h
    port map (
            O => \N__55451\,
            I => \N__55442\
        );

    \I__12327\ : Span4Mux_v
    port map (
            O => \N__55448\,
            I => \N__55439\
        );

    \I__12326\ : Span4Mux_v
    port map (
            O => \N__55445\,
            I => \N__55436\
        );

    \I__12325\ : Sp12to4
    port map (
            O => \N__55442\,
            I => \N__55433\
        );

    \I__12324\ : Span4Mux_v
    port map (
            O => \N__55439\,
            I => \N__55430\
        );

    \I__12323\ : Sp12to4
    port map (
            O => \N__55436\,
            I => \N__55425\
        );

    \I__12322\ : Span12Mux_v
    port map (
            O => \N__55433\,
            I => \N__55425\
        );

    \I__12321\ : Odrv4
    port map (
            O => \N__55430\,
            I => n11461
        );

    \I__12320\ : Odrv12
    port map (
            O => \N__55425\,
            I => n11461
        );

    \I__12319\ : InMux
    port map (
            O => \N__55420\,
            I => \N__55417\
        );

    \I__12318\ : LocalMux
    port map (
            O => \N__55417\,
            I => \N__55414\
        );

    \I__12317\ : Odrv4
    port map (
            O => \N__55414\,
            I => \c0.n11626\
        );

    \I__12316\ : InMux
    port map (
            O => \N__55411\,
            I => \N__55408\
        );

    \I__12315\ : LocalMux
    port map (
            O => \N__55408\,
            I => \N__55405\
        );

    \I__12314\ : Odrv12
    port map (
            O => \N__55405\,
            I => \c0.n21_adj_3205\
        );

    \I__12313\ : CascadeMux
    port map (
            O => \N__55402\,
            I => \N__55399\
        );

    \I__12312\ : InMux
    port map (
            O => \N__55399\,
            I => \N__55396\
        );

    \I__12311\ : LocalMux
    port map (
            O => \N__55396\,
            I => \N__55393\
        );

    \I__12310\ : Span4Mux_v
    port map (
            O => \N__55393\,
            I => \N__55390\
        );

    \I__12309\ : Span4Mux_h
    port map (
            O => \N__55390\,
            I => \N__55387\
        );

    \I__12308\ : Odrv4
    port map (
            O => \N__55387\,
            I => \c0.n28_adj_3428\
        );

    \I__12307\ : InMux
    port map (
            O => \N__55384\,
            I => \N__55379\
        );

    \I__12306\ : InMux
    port map (
            O => \N__55383\,
            I => \N__55374\
        );

    \I__12305\ : InMux
    port map (
            O => \N__55382\,
            I => \N__55371\
        );

    \I__12304\ : LocalMux
    port map (
            O => \N__55379\,
            I => \N__55368\
        );

    \I__12303\ : InMux
    port map (
            O => \N__55378\,
            I => \N__55365\
        );

    \I__12302\ : InMux
    port map (
            O => \N__55377\,
            I => \N__55361\
        );

    \I__12301\ : LocalMux
    port map (
            O => \N__55374\,
            I => \N__55358\
        );

    \I__12300\ : LocalMux
    port map (
            O => \N__55371\,
            I => \N__55355\
        );

    \I__12299\ : Span4Mux_h
    port map (
            O => \N__55368\,
            I => \N__55350\
        );

    \I__12298\ : LocalMux
    port map (
            O => \N__55365\,
            I => \N__55350\
        );

    \I__12297\ : InMux
    port map (
            O => \N__55364\,
            I => \N__55346\
        );

    \I__12296\ : LocalMux
    port map (
            O => \N__55361\,
            I => \N__55341\
        );

    \I__12295\ : Span4Mux_v
    port map (
            O => \N__55358\,
            I => \N__55338\
        );

    \I__12294\ : Span4Mux_v
    port map (
            O => \N__55355\,
            I => \N__55333\
        );

    \I__12293\ : Span4Mux_v
    port map (
            O => \N__55350\,
            I => \N__55333\
        );

    \I__12292\ : InMux
    port map (
            O => \N__55349\,
            I => \N__55330\
        );

    \I__12291\ : LocalMux
    port map (
            O => \N__55346\,
            I => \N__55327\
        );

    \I__12290\ : InMux
    port map (
            O => \N__55345\,
            I => \N__55322\
        );

    \I__12289\ : InMux
    port map (
            O => \N__55344\,
            I => \N__55322\
        );

    \I__12288\ : Odrv4
    port map (
            O => \N__55341\,
            I => data_in_frame_1_5
        );

    \I__12287\ : Odrv4
    port map (
            O => \N__55338\,
            I => data_in_frame_1_5
        );

    \I__12286\ : Odrv4
    port map (
            O => \N__55333\,
            I => data_in_frame_1_5
        );

    \I__12285\ : LocalMux
    port map (
            O => \N__55330\,
            I => data_in_frame_1_5
        );

    \I__12284\ : Odrv12
    port map (
            O => \N__55327\,
            I => data_in_frame_1_5
        );

    \I__12283\ : LocalMux
    port map (
            O => \N__55322\,
            I => data_in_frame_1_5
        );

    \I__12282\ : CascadeMux
    port map (
            O => \N__55309\,
            I => \N__55305\
        );

    \I__12281\ : InMux
    port map (
            O => \N__55308\,
            I => \N__55300\
        );

    \I__12280\ : InMux
    port map (
            O => \N__55305\,
            I => \N__55300\
        );

    \I__12279\ : LocalMux
    port map (
            O => \N__55300\,
            I => \N__55297\
        );

    \I__12278\ : Odrv12
    port map (
            O => \N__55297\,
            I => \c0.n7_adj_3509\
        );

    \I__12277\ : CascadeMux
    port map (
            O => \N__55294\,
            I => \c0.n7_adj_3509_cascade_\
        );

    \I__12276\ : CascadeMux
    port map (
            O => \N__55291\,
            I => \N__55288\
        );

    \I__12275\ : InMux
    port map (
            O => \N__55288\,
            I => \N__55285\
        );

    \I__12274\ : LocalMux
    port map (
            O => \N__55285\,
            I => \N__55281\
        );

    \I__12273\ : InMux
    port map (
            O => \N__55284\,
            I => \N__55278\
        );

    \I__12272\ : Span4Mux_v
    port map (
            O => \N__55281\,
            I => \N__55272\
        );

    \I__12271\ : LocalMux
    port map (
            O => \N__55278\,
            I => \N__55272\
        );

    \I__12270\ : InMux
    port map (
            O => \N__55277\,
            I => \N__55269\
        );

    \I__12269\ : Odrv4
    port map (
            O => \N__55272\,
            I => \c0.n10_adj_3012\
        );

    \I__12268\ : LocalMux
    port map (
            O => \N__55269\,
            I => \c0.n10_adj_3012\
        );

    \I__12267\ : InMux
    port map (
            O => \N__55264\,
            I => \N__55260\
        );

    \I__12266\ : InMux
    port map (
            O => \N__55263\,
            I => \N__55257\
        );

    \I__12265\ : LocalMux
    port map (
            O => \N__55260\,
            I => \N__55254\
        );

    \I__12264\ : LocalMux
    port map (
            O => \N__55257\,
            I => \N__55251\
        );

    \I__12263\ : Span4Mux_h
    port map (
            O => \N__55254\,
            I => \N__55248\
        );

    \I__12262\ : Span4Mux_h
    port map (
            O => \N__55251\,
            I => \N__55245\
        );

    \I__12261\ : Odrv4
    port map (
            O => \N__55248\,
            I => \c0.n45\
        );

    \I__12260\ : Odrv4
    port map (
            O => \N__55245\,
            I => \c0.n45\
        );

    \I__12259\ : InMux
    port map (
            O => \N__55240\,
            I => \N__55236\
        );

    \I__12258\ : InMux
    port map (
            O => \N__55239\,
            I => \N__55231\
        );

    \I__12257\ : LocalMux
    port map (
            O => \N__55236\,
            I => \N__55228\
        );

    \I__12256\ : InMux
    port map (
            O => \N__55235\,
            I => \N__55225\
        );

    \I__12255\ : CascadeMux
    port map (
            O => \N__55234\,
            I => \N__55222\
        );

    \I__12254\ : LocalMux
    port map (
            O => \N__55231\,
            I => \N__55219\
        );

    \I__12253\ : Span4Mux_v
    port map (
            O => \N__55228\,
            I => \N__55214\
        );

    \I__12252\ : LocalMux
    port map (
            O => \N__55225\,
            I => \N__55214\
        );

    \I__12251\ : InMux
    port map (
            O => \N__55222\,
            I => \N__55209\
        );

    \I__12250\ : Span4Mux_v
    port map (
            O => \N__55219\,
            I => \N__55206\
        );

    \I__12249\ : Span4Mux_h
    port map (
            O => \N__55214\,
            I => \N__55203\
        );

    \I__12248\ : InMux
    port map (
            O => \N__55213\,
            I => \N__55200\
        );

    \I__12247\ : InMux
    port map (
            O => \N__55212\,
            I => \N__55197\
        );

    \I__12246\ : LocalMux
    port map (
            O => \N__55209\,
            I => \c0.data_in_frame_4_1\
        );

    \I__12245\ : Odrv4
    port map (
            O => \N__55206\,
            I => \c0.data_in_frame_4_1\
        );

    \I__12244\ : Odrv4
    port map (
            O => \N__55203\,
            I => \c0.data_in_frame_4_1\
        );

    \I__12243\ : LocalMux
    port map (
            O => \N__55200\,
            I => \c0.data_in_frame_4_1\
        );

    \I__12242\ : LocalMux
    port map (
            O => \N__55197\,
            I => \c0.data_in_frame_4_1\
        );

    \I__12241\ : CascadeMux
    port map (
            O => \N__55186\,
            I => \N__55175\
        );

    \I__12240\ : InMux
    port map (
            O => \N__55185\,
            I => \N__55172\
        );

    \I__12239\ : InMux
    port map (
            O => \N__55184\,
            I => \N__55169\
        );

    \I__12238\ : InMux
    port map (
            O => \N__55183\,
            I => \N__55166\
        );

    \I__12237\ : InMux
    port map (
            O => \N__55182\,
            I => \N__55157\
        );

    \I__12236\ : InMux
    port map (
            O => \N__55181\,
            I => \N__55157\
        );

    \I__12235\ : InMux
    port map (
            O => \N__55180\,
            I => \N__55154\
        );

    \I__12234\ : InMux
    port map (
            O => \N__55179\,
            I => \N__55151\
        );

    \I__12233\ : CascadeMux
    port map (
            O => \N__55178\,
            I => \N__55148\
        );

    \I__12232\ : InMux
    port map (
            O => \N__55175\,
            I => \N__55144\
        );

    \I__12231\ : LocalMux
    port map (
            O => \N__55172\,
            I => \N__55137\
        );

    \I__12230\ : LocalMux
    port map (
            O => \N__55169\,
            I => \N__55137\
        );

    \I__12229\ : LocalMux
    port map (
            O => \N__55166\,
            I => \N__55137\
        );

    \I__12228\ : InMux
    port map (
            O => \N__55165\,
            I => \N__55130\
        );

    \I__12227\ : InMux
    port map (
            O => \N__55164\,
            I => \N__55130\
        );

    \I__12226\ : InMux
    port map (
            O => \N__55163\,
            I => \N__55130\
        );

    \I__12225\ : CascadeMux
    port map (
            O => \N__55162\,
            I => \N__55124\
        );

    \I__12224\ : LocalMux
    port map (
            O => \N__55157\,
            I => \N__55121\
        );

    \I__12223\ : LocalMux
    port map (
            O => \N__55154\,
            I => \N__55118\
        );

    \I__12222\ : LocalMux
    port map (
            O => \N__55151\,
            I => \N__55115\
        );

    \I__12221\ : InMux
    port map (
            O => \N__55148\,
            I => \N__55110\
        );

    \I__12220\ : InMux
    port map (
            O => \N__55147\,
            I => \N__55110\
        );

    \I__12219\ : LocalMux
    port map (
            O => \N__55144\,
            I => \N__55105\
        );

    \I__12218\ : Span4Mux_v
    port map (
            O => \N__55137\,
            I => \N__55100\
        );

    \I__12217\ : LocalMux
    port map (
            O => \N__55130\,
            I => \N__55100\
        );

    \I__12216\ : InMux
    port map (
            O => \N__55129\,
            I => \N__55095\
        );

    \I__12215\ : InMux
    port map (
            O => \N__55128\,
            I => \N__55095\
        );

    \I__12214\ : InMux
    port map (
            O => \N__55127\,
            I => \N__55092\
        );

    \I__12213\ : InMux
    port map (
            O => \N__55124\,
            I => \N__55089\
        );

    \I__12212\ : Span4Mux_v
    port map (
            O => \N__55121\,
            I => \N__55080\
        );

    \I__12211\ : Span4Mux_v
    port map (
            O => \N__55118\,
            I => \N__55080\
        );

    \I__12210\ : Span4Mux_h
    port map (
            O => \N__55115\,
            I => \N__55080\
        );

    \I__12209\ : LocalMux
    port map (
            O => \N__55110\,
            I => \N__55080\
        );

    \I__12208\ : InMux
    port map (
            O => \N__55109\,
            I => \N__55077\
        );

    \I__12207\ : InMux
    port map (
            O => \N__55108\,
            I => \N__55074\
        );

    \I__12206\ : Span4Mux_v
    port map (
            O => \N__55105\,
            I => \N__55069\
        );

    \I__12205\ : Span4Mux_h
    port map (
            O => \N__55100\,
            I => \N__55069\
        );

    \I__12204\ : LocalMux
    port map (
            O => \N__55095\,
            I => data_in_frame_0_6
        );

    \I__12203\ : LocalMux
    port map (
            O => \N__55092\,
            I => data_in_frame_0_6
        );

    \I__12202\ : LocalMux
    port map (
            O => \N__55089\,
            I => data_in_frame_0_6
        );

    \I__12201\ : Odrv4
    port map (
            O => \N__55080\,
            I => data_in_frame_0_6
        );

    \I__12200\ : LocalMux
    port map (
            O => \N__55077\,
            I => data_in_frame_0_6
        );

    \I__12199\ : LocalMux
    port map (
            O => \N__55074\,
            I => data_in_frame_0_6
        );

    \I__12198\ : Odrv4
    port map (
            O => \N__55069\,
            I => data_in_frame_0_6
        );

    \I__12197\ : InMux
    port map (
            O => \N__55054\,
            I => \N__55049\
        );

    \I__12196\ : InMux
    port map (
            O => \N__55053\,
            I => \N__55046\
        );

    \I__12195\ : InMux
    port map (
            O => \N__55052\,
            I => \N__55043\
        );

    \I__12194\ : LocalMux
    port map (
            O => \N__55049\,
            I => \N__55040\
        );

    \I__12193\ : LocalMux
    port map (
            O => \N__55046\,
            I => \N__55035\
        );

    \I__12192\ : LocalMux
    port map (
            O => \N__55043\,
            I => \N__55035\
        );

    \I__12191\ : Span4Mux_h
    port map (
            O => \N__55040\,
            I => \N__55028\
        );

    \I__12190\ : Span4Mux_h
    port map (
            O => \N__55035\,
            I => \N__55025\
        );

    \I__12189\ : InMux
    port map (
            O => \N__55034\,
            I => \N__55022\
        );

    \I__12188\ : InMux
    port map (
            O => \N__55033\,
            I => \N__55017\
        );

    \I__12187\ : InMux
    port map (
            O => \N__55032\,
            I => \N__55017\
        );

    \I__12186\ : CascadeMux
    port map (
            O => \N__55031\,
            I => \N__55011\
        );

    \I__12185\ : Span4Mux_h
    port map (
            O => \N__55028\,
            I => \N__55007\
        );

    \I__12184\ : Span4Mux_v
    port map (
            O => \N__55025\,
            I => \N__55000\
        );

    \I__12183\ : LocalMux
    port map (
            O => \N__55022\,
            I => \N__55000\
        );

    \I__12182\ : LocalMux
    port map (
            O => \N__55017\,
            I => \N__55000\
        );

    \I__12181\ : InMux
    port map (
            O => \N__55016\,
            I => \N__54995\
        );

    \I__12180\ : InMux
    port map (
            O => \N__55015\,
            I => \N__54995\
        );

    \I__12179\ : InMux
    port map (
            O => \N__55014\,
            I => \N__54992\
        );

    \I__12178\ : InMux
    port map (
            O => \N__55011\,
            I => \N__54987\
        );

    \I__12177\ : InMux
    port map (
            O => \N__55010\,
            I => \N__54987\
        );

    \I__12176\ : Odrv4
    port map (
            O => \N__55007\,
            I => data_in_frame_1_0
        );

    \I__12175\ : Odrv4
    port map (
            O => \N__55000\,
            I => data_in_frame_1_0
        );

    \I__12174\ : LocalMux
    port map (
            O => \N__54995\,
            I => data_in_frame_1_0
        );

    \I__12173\ : LocalMux
    port map (
            O => \N__54992\,
            I => data_in_frame_1_0
        );

    \I__12172\ : LocalMux
    port map (
            O => \N__54987\,
            I => data_in_frame_1_0
        );

    \I__12171\ : InMux
    port map (
            O => \N__54976\,
            I => \N__54973\
        );

    \I__12170\ : LocalMux
    port map (
            O => \N__54973\,
            I => \N__54970\
        );

    \I__12169\ : Span4Mux_v
    port map (
            O => \N__54970\,
            I => \N__54967\
        );

    \I__12168\ : Span4Mux_h
    port map (
            O => \N__54967\,
            I => \N__54962\
        );

    \I__12167\ : InMux
    port map (
            O => \N__54966\,
            I => \N__54957\
        );

    \I__12166\ : InMux
    port map (
            O => \N__54965\,
            I => \N__54957\
        );

    \I__12165\ : Odrv4
    port map (
            O => \N__54962\,
            I => \c0.n20341\
        );

    \I__12164\ : LocalMux
    port map (
            O => \N__54957\,
            I => \c0.n20341\
        );

    \I__12163\ : InMux
    port map (
            O => \N__54952\,
            I => \N__54949\
        );

    \I__12162\ : LocalMux
    port map (
            O => \N__54949\,
            I => \N__54946\
        );

    \I__12161\ : Odrv4
    port map (
            O => \N__54946\,
            I => \c0.n58_adj_3497\
        );

    \I__12160\ : InMux
    port map (
            O => \N__54943\,
            I => \N__54940\
        );

    \I__12159\ : LocalMux
    port map (
            O => \N__54940\,
            I => \c0.n56_adj_3505\
        );

    \I__12158\ : InMux
    port map (
            O => \N__54937\,
            I => \N__54934\
        );

    \I__12157\ : LocalMux
    port map (
            O => \N__54934\,
            I => \N__54931\
        );

    \I__12156\ : Span4Mux_h
    port map (
            O => \N__54931\,
            I => \N__54928\
        );

    \I__12155\ : Odrv4
    port map (
            O => \N__54928\,
            I => \c0.n64_adj_3506\
        );

    \I__12154\ : InMux
    port map (
            O => \N__54925\,
            I => \N__54922\
        );

    \I__12153\ : LocalMux
    port map (
            O => \N__54922\,
            I => \N__54919\
        );

    \I__12152\ : Span12Mux_s10_h
    port map (
            O => \N__54919\,
            I => \N__54916\
        );

    \I__12151\ : Odrv12
    port map (
            O => \N__54916\,
            I => \c0.n19217\
        );

    \I__12150\ : CascadeMux
    port map (
            O => \N__54913\,
            I => \c0.n4_adj_3036_cascade_\
        );

    \I__12149\ : InMux
    port map (
            O => \N__54910\,
            I => \N__54907\
        );

    \I__12148\ : LocalMux
    port map (
            O => \N__54907\,
            I => \c0.n57_adj_3499\
        );

    \I__12147\ : CascadeMux
    port map (
            O => \N__54904\,
            I => \c0.n11478_cascade_\
        );

    \I__12146\ : InMux
    port map (
            O => \N__54901\,
            I => \N__54898\
        );

    \I__12145\ : LocalMux
    port map (
            O => \N__54898\,
            I => \c0.n81\
        );

    \I__12144\ : InMux
    port map (
            O => \N__54895\,
            I => \N__54889\
        );

    \I__12143\ : CascadeMux
    port map (
            O => \N__54894\,
            I => \N__54884\
        );

    \I__12142\ : InMux
    port map (
            O => \N__54893\,
            I => \N__54881\
        );

    \I__12141\ : InMux
    port map (
            O => \N__54892\,
            I => \N__54877\
        );

    \I__12140\ : LocalMux
    port map (
            O => \N__54889\,
            I => \N__54873\
        );

    \I__12139\ : InMux
    port map (
            O => \N__54888\,
            I => \N__54868\
        );

    \I__12138\ : InMux
    port map (
            O => \N__54887\,
            I => \N__54868\
        );

    \I__12137\ : InMux
    port map (
            O => \N__54884\,
            I => \N__54865\
        );

    \I__12136\ : LocalMux
    port map (
            O => \N__54881\,
            I => \N__54862\
        );

    \I__12135\ : InMux
    port map (
            O => \N__54880\,
            I => \N__54859\
        );

    \I__12134\ : LocalMux
    port map (
            O => \N__54877\,
            I => \N__54855\
        );

    \I__12133\ : InMux
    port map (
            O => \N__54876\,
            I => \N__54852\
        );

    \I__12132\ : Span4Mux_h
    port map (
            O => \N__54873\,
            I => \N__54846\
        );

    \I__12131\ : LocalMux
    port map (
            O => \N__54868\,
            I => \N__54846\
        );

    \I__12130\ : LocalMux
    port map (
            O => \N__54865\,
            I => \N__54843\
        );

    \I__12129\ : Span4Mux_h
    port map (
            O => \N__54862\,
            I => \N__54837\
        );

    \I__12128\ : LocalMux
    port map (
            O => \N__54859\,
            I => \N__54837\
        );

    \I__12127\ : CascadeMux
    port map (
            O => \N__54858\,
            I => \N__54831\
        );

    \I__12126\ : Span12Mux_h
    port map (
            O => \N__54855\,
            I => \N__54828\
        );

    \I__12125\ : LocalMux
    port map (
            O => \N__54852\,
            I => \N__54825\
        );

    \I__12124\ : InMux
    port map (
            O => \N__54851\,
            I => \N__54822\
        );

    \I__12123\ : Span4Mux_v
    port map (
            O => \N__54846\,
            I => \N__54819\
        );

    \I__12122\ : Span4Mux_h
    port map (
            O => \N__54843\,
            I => \N__54816\
        );

    \I__12121\ : InMux
    port map (
            O => \N__54842\,
            I => \N__54813\
        );

    \I__12120\ : Span4Mux_h
    port map (
            O => \N__54837\,
            I => \N__54810\
        );

    \I__12119\ : InMux
    port map (
            O => \N__54836\,
            I => \N__54807\
        );

    \I__12118\ : InMux
    port map (
            O => \N__54835\,
            I => \N__54800\
        );

    \I__12117\ : InMux
    port map (
            O => \N__54834\,
            I => \N__54800\
        );

    \I__12116\ : InMux
    port map (
            O => \N__54831\,
            I => \N__54800\
        );

    \I__12115\ : Odrv12
    port map (
            O => \N__54828\,
            I => data_in_frame_1_6
        );

    \I__12114\ : Odrv12
    port map (
            O => \N__54825\,
            I => data_in_frame_1_6
        );

    \I__12113\ : LocalMux
    port map (
            O => \N__54822\,
            I => data_in_frame_1_6
        );

    \I__12112\ : Odrv4
    port map (
            O => \N__54819\,
            I => data_in_frame_1_6
        );

    \I__12111\ : Odrv4
    port map (
            O => \N__54816\,
            I => data_in_frame_1_6
        );

    \I__12110\ : LocalMux
    port map (
            O => \N__54813\,
            I => data_in_frame_1_6
        );

    \I__12109\ : Odrv4
    port map (
            O => \N__54810\,
            I => data_in_frame_1_6
        );

    \I__12108\ : LocalMux
    port map (
            O => \N__54807\,
            I => data_in_frame_1_6
        );

    \I__12107\ : LocalMux
    port map (
            O => \N__54800\,
            I => data_in_frame_1_6
        );

    \I__12106\ : InMux
    port map (
            O => \N__54781\,
            I => \N__54778\
        );

    \I__12105\ : LocalMux
    port map (
            O => \N__54778\,
            I => \c0.n11526\
        );

    \I__12104\ : CascadeMux
    port map (
            O => \N__54775\,
            I => \N__54772\
        );

    \I__12103\ : InMux
    port map (
            O => \N__54772\,
            I => \N__54767\
        );

    \I__12102\ : InMux
    port map (
            O => \N__54771\,
            I => \N__54762\
        );

    \I__12101\ : InMux
    port map (
            O => \N__54770\,
            I => \N__54762\
        );

    \I__12100\ : LocalMux
    port map (
            O => \N__54767\,
            I => \c0.data_in_frame_6_5\
        );

    \I__12099\ : LocalMux
    port map (
            O => \N__54762\,
            I => \c0.data_in_frame_6_5\
        );

    \I__12098\ : CascadeMux
    port map (
            O => \N__54757\,
            I => \N__54754\
        );

    \I__12097\ : InMux
    port map (
            O => \N__54754\,
            I => \N__54751\
        );

    \I__12096\ : LocalMux
    port map (
            O => \N__54751\,
            I => \N__54747\
        );

    \I__12095\ : InMux
    port map (
            O => \N__54750\,
            I => \N__54744\
        );

    \I__12094\ : Span4Mux_h
    port map (
            O => \N__54747\,
            I => \N__54741\
        );

    \I__12093\ : LocalMux
    port map (
            O => \N__54744\,
            I => \N__54738\
        );

    \I__12092\ : Odrv4
    port map (
            O => \N__54741\,
            I => \c0.n11549\
        );

    \I__12091\ : Odrv4
    port map (
            O => \N__54738\,
            I => \c0.n11549\
        );

    \I__12090\ : InMux
    port map (
            O => \N__54733\,
            I => \N__54728\
        );

    \I__12089\ : InMux
    port map (
            O => \N__54732\,
            I => \N__54722\
        );

    \I__12088\ : InMux
    port map (
            O => \N__54731\,
            I => \N__54722\
        );

    \I__12087\ : LocalMux
    port map (
            O => \N__54728\,
            I => \N__54719\
        );

    \I__12086\ : InMux
    port map (
            O => \N__54727\,
            I => \N__54716\
        );

    \I__12085\ : LocalMux
    port map (
            O => \N__54722\,
            I => \N__54713\
        );

    \I__12084\ : Odrv12
    port map (
            O => \N__54719\,
            I => \c0.n11651\
        );

    \I__12083\ : LocalMux
    port map (
            O => \N__54716\,
            I => \c0.n11651\
        );

    \I__12082\ : Odrv4
    port map (
            O => \N__54713\,
            I => \c0.n11651\
        );

    \I__12081\ : InMux
    port map (
            O => \N__54706\,
            I => \N__54703\
        );

    \I__12080\ : LocalMux
    port map (
            O => \N__54703\,
            I => \N__54700\
        );

    \I__12079\ : Span4Mux_h
    port map (
            O => \N__54700\,
            I => \N__54697\
        );

    \I__12078\ : Span4Mux_h
    port map (
            O => \N__54697\,
            I => \N__54694\
        );

    \I__12077\ : Odrv4
    port map (
            O => \N__54694\,
            I => \c0.n27_adj_3457\
        );

    \I__12076\ : InMux
    port map (
            O => \N__54691\,
            I => \N__54688\
        );

    \I__12075\ : LocalMux
    port map (
            O => \N__54688\,
            I => \N__54685\
        );

    \I__12074\ : Span4Mux_h
    port map (
            O => \N__54685\,
            I => \N__54681\
        );

    \I__12073\ : CascadeMux
    port map (
            O => \N__54684\,
            I => \N__54677\
        );

    \I__12072\ : Span4Mux_v
    port map (
            O => \N__54681\,
            I => \N__54668\
        );

    \I__12071\ : InMux
    port map (
            O => \N__54680\,
            I => \N__54665\
        );

    \I__12070\ : InMux
    port map (
            O => \N__54677\,
            I => \N__54658\
        );

    \I__12069\ : InMux
    port map (
            O => \N__54676\,
            I => \N__54658\
        );

    \I__12068\ : InMux
    port map (
            O => \N__54675\,
            I => \N__54658\
        );

    \I__12067\ : InMux
    port map (
            O => \N__54674\,
            I => \N__54655\
        );

    \I__12066\ : InMux
    port map (
            O => \N__54673\,
            I => \N__54652\
        );

    \I__12065\ : InMux
    port map (
            O => \N__54672\,
            I => \N__54647\
        );

    \I__12064\ : InMux
    port map (
            O => \N__54671\,
            I => \N__54647\
        );

    \I__12063\ : Odrv4
    port map (
            O => \N__54668\,
            I => data_in_frame_1_7
        );

    \I__12062\ : LocalMux
    port map (
            O => \N__54665\,
            I => data_in_frame_1_7
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__54658\,
            I => data_in_frame_1_7
        );

    \I__12060\ : LocalMux
    port map (
            O => \N__54655\,
            I => data_in_frame_1_7
        );

    \I__12059\ : LocalMux
    port map (
            O => \N__54652\,
            I => data_in_frame_1_7
        );

    \I__12058\ : LocalMux
    port map (
            O => \N__54647\,
            I => data_in_frame_1_7
        );

    \I__12057\ : InMux
    port map (
            O => \N__54634\,
            I => \N__54631\
        );

    \I__12056\ : LocalMux
    port map (
            O => \N__54631\,
            I => \c0.n12_adj_3378\
        );

    \I__12055\ : CascadeMux
    port map (
            O => \N__54628\,
            I => \N__54624\
        );

    \I__12054\ : CascadeMux
    port map (
            O => \N__54627\,
            I => \N__54620\
        );

    \I__12053\ : InMux
    port map (
            O => \N__54624\,
            I => \N__54617\
        );

    \I__12052\ : InMux
    port map (
            O => \N__54623\,
            I => \N__54614\
        );

    \I__12051\ : InMux
    port map (
            O => \N__54620\,
            I => \N__54609\
        );

    \I__12050\ : LocalMux
    port map (
            O => \N__54617\,
            I => \N__54606\
        );

    \I__12049\ : LocalMux
    port map (
            O => \N__54614\,
            I => \N__54603\
        );

    \I__12048\ : InMux
    port map (
            O => \N__54613\,
            I => \N__54598\
        );

    \I__12047\ : InMux
    port map (
            O => \N__54612\,
            I => \N__54598\
        );

    \I__12046\ : LocalMux
    port map (
            O => \N__54609\,
            I => \c0.data_in_frame_2_1\
        );

    \I__12045\ : Odrv12
    port map (
            O => \N__54606\,
            I => \c0.data_in_frame_2_1\
        );

    \I__12044\ : Odrv12
    port map (
            O => \N__54603\,
            I => \c0.data_in_frame_2_1\
        );

    \I__12043\ : LocalMux
    port map (
            O => \N__54598\,
            I => \c0.data_in_frame_2_1\
        );

    \I__12042\ : InMux
    port map (
            O => \N__54589\,
            I => \N__54586\
        );

    \I__12041\ : LocalMux
    port map (
            O => \N__54586\,
            I => \N__54583\
        );

    \I__12040\ : Odrv12
    port map (
            O => \N__54583\,
            I => \c0.n34_adj_3326\
        );

    \I__12039\ : CascadeMux
    port map (
            O => \N__54580\,
            I => \N__54576\
        );

    \I__12038\ : InMux
    port map (
            O => \N__54579\,
            I => \N__54571\
        );

    \I__12037\ : InMux
    port map (
            O => \N__54576\,
            I => \N__54571\
        );

    \I__12036\ : LocalMux
    port map (
            O => \N__54571\,
            I => \c0.n13_adj_3344\
        );

    \I__12035\ : InMux
    port map (
            O => \N__54568\,
            I => \N__54564\
        );

    \I__12034\ : CascadeMux
    port map (
            O => \N__54567\,
            I => \N__54561\
        );

    \I__12033\ : LocalMux
    port map (
            O => \N__54564\,
            I => \N__54557\
        );

    \I__12032\ : InMux
    port map (
            O => \N__54561\,
            I => \N__54553\
        );

    \I__12031\ : InMux
    port map (
            O => \N__54560\,
            I => \N__54550\
        );

    \I__12030\ : Span12Mux_h
    port map (
            O => \N__54557\,
            I => \N__54547\
        );

    \I__12029\ : InMux
    port map (
            O => \N__54556\,
            I => \N__54544\
        );

    \I__12028\ : LocalMux
    port map (
            O => \N__54553\,
            I => \N__54541\
        );

    \I__12027\ : LocalMux
    port map (
            O => \N__54550\,
            I => \c0.n23_adj_3076\
        );

    \I__12026\ : Odrv12
    port map (
            O => \N__54547\,
            I => \c0.n23_adj_3076\
        );

    \I__12025\ : LocalMux
    port map (
            O => \N__54544\,
            I => \c0.n23_adj_3076\
        );

    \I__12024\ : Odrv4
    port map (
            O => \N__54541\,
            I => \c0.n23_adj_3076\
        );

    \I__12023\ : InMux
    port map (
            O => \N__54532\,
            I => \N__54525\
        );

    \I__12022\ : InMux
    port map (
            O => \N__54531\,
            I => \N__54525\
        );

    \I__12021\ : InMux
    port map (
            O => \N__54530\,
            I => \N__54522\
        );

    \I__12020\ : LocalMux
    port map (
            O => \N__54525\,
            I => \N__54519\
        );

    \I__12019\ : LocalMux
    port map (
            O => \N__54522\,
            I => \N__54515\
        );

    \I__12018\ : Span4Mux_v
    port map (
            O => \N__54519\,
            I => \N__54512\
        );

    \I__12017\ : InMux
    port map (
            O => \N__54518\,
            I => \N__54509\
        );

    \I__12016\ : Odrv4
    port map (
            O => \N__54515\,
            I => \c0.n19424\
        );

    \I__12015\ : Odrv4
    port map (
            O => \N__54512\,
            I => \c0.n19424\
        );

    \I__12014\ : LocalMux
    port map (
            O => \N__54509\,
            I => \c0.n19424\
        );

    \I__12013\ : CascadeMux
    port map (
            O => \N__54502\,
            I => \N__54499\
        );

    \I__12012\ : InMux
    port map (
            O => \N__54499\,
            I => \N__54496\
        );

    \I__12011\ : LocalMux
    port map (
            O => \N__54496\,
            I => \N__54493\
        );

    \I__12010\ : Span4Mux_v
    port map (
            O => \N__54493\,
            I => \N__54489\
        );

    \I__12009\ : InMux
    port map (
            O => \N__54492\,
            I => \N__54486\
        );

    \I__12008\ : Odrv4
    port map (
            O => \N__54489\,
            I => \c0.n7_adj_3029\
        );

    \I__12007\ : LocalMux
    port map (
            O => \N__54486\,
            I => \c0.n7_adj_3029\
        );

    \I__12006\ : CascadeMux
    port map (
            O => \N__54481\,
            I => \N__54476\
        );

    \I__12005\ : InMux
    port map (
            O => \N__54480\,
            I => \N__54473\
        );

    \I__12004\ : CascadeMux
    port map (
            O => \N__54479\,
            I => \N__54469\
        );

    \I__12003\ : InMux
    port map (
            O => \N__54476\,
            I => \N__54463\
        );

    \I__12002\ : LocalMux
    port map (
            O => \N__54473\,
            I => \N__54456\
        );

    \I__12001\ : CascadeMux
    port map (
            O => \N__54472\,
            I => \N__54453\
        );

    \I__12000\ : InMux
    port map (
            O => \N__54469\,
            I => \N__54449\
        );

    \I__11999\ : InMux
    port map (
            O => \N__54468\,
            I => \N__54446\
        );

    \I__11998\ : InMux
    port map (
            O => \N__54467\,
            I => \N__54443\
        );

    \I__11997\ : InMux
    port map (
            O => \N__54466\,
            I => \N__54439\
        );

    \I__11996\ : LocalMux
    port map (
            O => \N__54463\,
            I => \N__54436\
        );

    \I__11995\ : InMux
    port map (
            O => \N__54462\,
            I => \N__54431\
        );

    \I__11994\ : InMux
    port map (
            O => \N__54461\,
            I => \N__54431\
        );

    \I__11993\ : InMux
    port map (
            O => \N__54460\,
            I => \N__54428\
        );

    \I__11992\ : CascadeMux
    port map (
            O => \N__54459\,
            I => \N__54424\
        );

    \I__11991\ : Span4Mux_v
    port map (
            O => \N__54456\,
            I => \N__54418\
        );

    \I__11990\ : InMux
    port map (
            O => \N__54453\,
            I => \N__54415\
        );

    \I__11989\ : InMux
    port map (
            O => \N__54452\,
            I => \N__54412\
        );

    \I__11988\ : LocalMux
    port map (
            O => \N__54449\,
            I => \N__54405\
        );

    \I__11987\ : LocalMux
    port map (
            O => \N__54446\,
            I => \N__54405\
        );

    \I__11986\ : LocalMux
    port map (
            O => \N__54443\,
            I => \N__54402\
        );

    \I__11985\ : InMux
    port map (
            O => \N__54442\,
            I => \N__54399\
        );

    \I__11984\ : LocalMux
    port map (
            O => \N__54439\,
            I => \N__54396\
        );

    \I__11983\ : Span4Mux_h
    port map (
            O => \N__54436\,
            I => \N__54388\
        );

    \I__11982\ : LocalMux
    port map (
            O => \N__54431\,
            I => \N__54388\
        );

    \I__11981\ : LocalMux
    port map (
            O => \N__54428\,
            I => \N__54388\
        );

    \I__11980\ : InMux
    port map (
            O => \N__54427\,
            I => \N__54385\
        );

    \I__11979\ : InMux
    port map (
            O => \N__54424\,
            I => \N__54378\
        );

    \I__11978\ : InMux
    port map (
            O => \N__54423\,
            I => \N__54378\
        );

    \I__11977\ : InMux
    port map (
            O => \N__54422\,
            I => \N__54373\
        );

    \I__11976\ : InMux
    port map (
            O => \N__54421\,
            I => \N__54373\
        );

    \I__11975\ : Span4Mux_h
    port map (
            O => \N__54418\,
            I => \N__54370\
        );

    \I__11974\ : LocalMux
    port map (
            O => \N__54415\,
            I => \N__54365\
        );

    \I__11973\ : LocalMux
    port map (
            O => \N__54412\,
            I => \N__54365\
        );

    \I__11972\ : InMux
    port map (
            O => \N__54411\,
            I => \N__54360\
        );

    \I__11971\ : InMux
    port map (
            O => \N__54410\,
            I => \N__54360\
        );

    \I__11970\ : Span4Mux_h
    port map (
            O => \N__54405\,
            I => \N__54351\
        );

    \I__11969\ : Span4Mux_v
    port map (
            O => \N__54402\,
            I => \N__54351\
        );

    \I__11968\ : LocalMux
    port map (
            O => \N__54399\,
            I => \N__54351\
        );

    \I__11967\ : Span4Mux_h
    port map (
            O => \N__54396\,
            I => \N__54351\
        );

    \I__11966\ : InMux
    port map (
            O => \N__54395\,
            I => \N__54348\
        );

    \I__11965\ : Span4Mux_h
    port map (
            O => \N__54388\,
            I => \N__54343\
        );

    \I__11964\ : LocalMux
    port map (
            O => \N__54385\,
            I => \N__54343\
        );

    \I__11963\ : InMux
    port map (
            O => \N__54384\,
            I => \N__54340\
        );

    \I__11962\ : InMux
    port map (
            O => \N__54383\,
            I => \N__54337\
        );

    \I__11961\ : LocalMux
    port map (
            O => \N__54378\,
            I => data_in_frame_0_4
        );

    \I__11960\ : LocalMux
    port map (
            O => \N__54373\,
            I => data_in_frame_0_4
        );

    \I__11959\ : Odrv4
    port map (
            O => \N__54370\,
            I => data_in_frame_0_4
        );

    \I__11958\ : Odrv12
    port map (
            O => \N__54365\,
            I => data_in_frame_0_4
        );

    \I__11957\ : LocalMux
    port map (
            O => \N__54360\,
            I => data_in_frame_0_4
        );

    \I__11956\ : Odrv4
    port map (
            O => \N__54351\,
            I => data_in_frame_0_4
        );

    \I__11955\ : LocalMux
    port map (
            O => \N__54348\,
            I => data_in_frame_0_4
        );

    \I__11954\ : Odrv4
    port map (
            O => \N__54343\,
            I => data_in_frame_0_4
        );

    \I__11953\ : LocalMux
    port map (
            O => \N__54340\,
            I => data_in_frame_0_4
        );

    \I__11952\ : LocalMux
    port map (
            O => \N__54337\,
            I => data_in_frame_0_4
        );

    \I__11951\ : CascadeMux
    port map (
            O => \N__54316\,
            I => \N__54312\
        );

    \I__11950\ : InMux
    port map (
            O => \N__54315\,
            I => \N__54309\
        );

    \I__11949\ : InMux
    port map (
            O => \N__54312\,
            I => \N__54305\
        );

    \I__11948\ : LocalMux
    port map (
            O => \N__54309\,
            I => \N__54302\
        );

    \I__11947\ : InMux
    port map (
            O => \N__54308\,
            I => \N__54299\
        );

    \I__11946\ : LocalMux
    port map (
            O => \N__54305\,
            I => \N__54291\
        );

    \I__11945\ : Span4Mux_h
    port map (
            O => \N__54302\,
            I => \N__54291\
        );

    \I__11944\ : LocalMux
    port map (
            O => \N__54299\,
            I => \N__54288\
        );

    \I__11943\ : InMux
    port map (
            O => \N__54298\,
            I => \N__54285\
        );

    \I__11942\ : InMux
    port map (
            O => \N__54297\,
            I => \N__54280\
        );

    \I__11941\ : InMux
    port map (
            O => \N__54296\,
            I => \N__54280\
        );

    \I__11940\ : Odrv4
    port map (
            O => \N__54291\,
            I => \c0.data_in_frame_2_3\
        );

    \I__11939\ : Odrv12
    port map (
            O => \N__54288\,
            I => \c0.data_in_frame_2_3\
        );

    \I__11938\ : LocalMux
    port map (
            O => \N__54285\,
            I => \c0.data_in_frame_2_3\
        );

    \I__11937\ : LocalMux
    port map (
            O => \N__54280\,
            I => \c0.data_in_frame_2_3\
        );

    \I__11936\ : InMux
    port map (
            O => \N__54271\,
            I => \N__54268\
        );

    \I__11935\ : LocalMux
    port map (
            O => \N__54268\,
            I => \N__54263\
        );

    \I__11934\ : InMux
    port map (
            O => \N__54267\,
            I => \N__54258\
        );

    \I__11933\ : CascadeMux
    port map (
            O => \N__54266\,
            I => \N__54255\
        );

    \I__11932\ : Span4Mux_v
    port map (
            O => \N__54263\,
            I => \N__54251\
        );

    \I__11931\ : InMux
    port map (
            O => \N__54262\,
            I => \N__54246\
        );

    \I__11930\ : InMux
    port map (
            O => \N__54261\,
            I => \N__54246\
        );

    \I__11929\ : LocalMux
    port map (
            O => \N__54258\,
            I => \N__54243\
        );

    \I__11928\ : InMux
    port map (
            O => \N__54255\,
            I => \N__54239\
        );

    \I__11927\ : InMux
    port map (
            O => \N__54254\,
            I => \N__54236\
        );

    \I__11926\ : Span4Mux_h
    port map (
            O => \N__54251\,
            I => \N__54233\
        );

    \I__11925\ : LocalMux
    port map (
            O => \N__54246\,
            I => \N__54230\
        );

    \I__11924\ : Span4Mux_h
    port map (
            O => \N__54243\,
            I => \N__54227\
        );

    \I__11923\ : InMux
    port map (
            O => \N__54242\,
            I => \N__54224\
        );

    \I__11922\ : LocalMux
    port map (
            O => \N__54239\,
            I => \c0.data_in_frame_4_4\
        );

    \I__11921\ : LocalMux
    port map (
            O => \N__54236\,
            I => \c0.data_in_frame_4_4\
        );

    \I__11920\ : Odrv4
    port map (
            O => \N__54233\,
            I => \c0.data_in_frame_4_4\
        );

    \I__11919\ : Odrv4
    port map (
            O => \N__54230\,
            I => \c0.data_in_frame_4_4\
        );

    \I__11918\ : Odrv4
    port map (
            O => \N__54227\,
            I => \c0.data_in_frame_4_4\
        );

    \I__11917\ : LocalMux
    port map (
            O => \N__54224\,
            I => \c0.data_in_frame_4_4\
        );

    \I__11916\ : InMux
    port map (
            O => \N__54211\,
            I => \N__54205\
        );

    \I__11915\ : InMux
    port map (
            O => \N__54210\,
            I => \N__54205\
        );

    \I__11914\ : LocalMux
    port map (
            O => \N__54205\,
            I => \N__54202\
        );

    \I__11913\ : Odrv4
    port map (
            O => \N__54202\,
            I => \c0.n8_adj_3345\
        );

    \I__11912\ : InMux
    port map (
            O => \N__54199\,
            I => \N__54195\
        );

    \I__11911\ : InMux
    port map (
            O => \N__54198\,
            I => \N__54192\
        );

    \I__11910\ : LocalMux
    port map (
            O => \N__54195\,
            I => \c0.n7_adj_3520\
        );

    \I__11909\ : LocalMux
    port map (
            O => \N__54192\,
            I => \c0.n7_adj_3520\
        );

    \I__11908\ : InMux
    port map (
            O => \N__54187\,
            I => \N__54178\
        );

    \I__11907\ : InMux
    port map (
            O => \N__54186\,
            I => \N__54178\
        );

    \I__11906\ : InMux
    port map (
            O => \N__54185\,
            I => \N__54178\
        );

    \I__11905\ : LocalMux
    port map (
            O => \N__54178\,
            I => \N__54175\
        );

    \I__11904\ : Odrv4
    port map (
            O => \N__54175\,
            I => \c0.n9_adj_3346\
        );

    \I__11903\ : CascadeMux
    port map (
            O => \N__54172\,
            I => \c0.n8_adj_3345_cascade_\
        );

    \I__11902\ : CascadeMux
    port map (
            O => \N__54169\,
            I => \c0.n11626_cascade_\
        );

    \I__11901\ : InMux
    port map (
            O => \N__54166\,
            I => \N__54163\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__54163\,
            I => \N__54159\
        );

    \I__11899\ : CascadeMux
    port map (
            O => \N__54162\,
            I => \N__54156\
        );

    \I__11898\ : Span4Mux_h
    port map (
            O => \N__54159\,
            I => \N__54152\
        );

    \I__11897\ : InMux
    port map (
            O => \N__54156\,
            I => \N__54149\
        );

    \I__11896\ : InMux
    port map (
            O => \N__54155\,
            I => \N__54146\
        );

    \I__11895\ : Span4Mux_v
    port map (
            O => \N__54152\,
            I => \N__54143\
        );

    \I__11894\ : LocalMux
    port map (
            O => \N__54149\,
            I => \c0.data_in_frame_8_7\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__54146\,
            I => \c0.data_in_frame_8_7\
        );

    \I__11892\ : Odrv4
    port map (
            O => \N__54143\,
            I => \c0.data_in_frame_8_7\
        );

    \I__11891\ : InMux
    port map (
            O => \N__54136\,
            I => \N__54131\
        );

    \I__11890\ : InMux
    port map (
            O => \N__54135\,
            I => \N__54127\
        );

    \I__11889\ : InMux
    port map (
            O => \N__54134\,
            I => \N__54123\
        );

    \I__11888\ : LocalMux
    port map (
            O => \N__54131\,
            I => \N__54119\
        );

    \I__11887\ : InMux
    port map (
            O => \N__54130\,
            I => \N__54116\
        );

    \I__11886\ : LocalMux
    port map (
            O => \N__54127\,
            I => \N__54112\
        );

    \I__11885\ : InMux
    port map (
            O => \N__54126\,
            I => \N__54109\
        );

    \I__11884\ : LocalMux
    port map (
            O => \N__54123\,
            I => \N__54106\
        );

    \I__11883\ : InMux
    port map (
            O => \N__54122\,
            I => \N__54103\
        );

    \I__11882\ : Span4Mux_v
    port map (
            O => \N__54119\,
            I => \N__54098\
        );

    \I__11881\ : LocalMux
    port map (
            O => \N__54116\,
            I => \N__54098\
        );

    \I__11880\ : InMux
    port map (
            O => \N__54115\,
            I => \N__54091\
        );

    \I__11879\ : Span4Mux_h
    port map (
            O => \N__54112\,
            I => \N__54088\
        );

    \I__11878\ : LocalMux
    port map (
            O => \N__54109\,
            I => \N__54079\
        );

    \I__11877\ : Span4Mux_h
    port map (
            O => \N__54106\,
            I => \N__54079\
        );

    \I__11876\ : LocalMux
    port map (
            O => \N__54103\,
            I => \N__54079\
        );

    \I__11875\ : Span4Mux_v
    port map (
            O => \N__54098\,
            I => \N__54079\
        );

    \I__11874\ : InMux
    port map (
            O => \N__54097\,
            I => \N__54070\
        );

    \I__11873\ : InMux
    port map (
            O => \N__54096\,
            I => \N__54070\
        );

    \I__11872\ : InMux
    port map (
            O => \N__54095\,
            I => \N__54070\
        );

    \I__11871\ : InMux
    port map (
            O => \N__54094\,
            I => \N__54070\
        );

    \I__11870\ : LocalMux
    port map (
            O => \N__54091\,
            I => \N__54067\
        );

    \I__11869\ : Odrv4
    port map (
            O => \N__54088\,
            I => data_in_frame_1_1
        );

    \I__11868\ : Odrv4
    port map (
            O => \N__54079\,
            I => data_in_frame_1_1
        );

    \I__11867\ : LocalMux
    port map (
            O => \N__54070\,
            I => data_in_frame_1_1
        );

    \I__11866\ : Odrv4
    port map (
            O => \N__54067\,
            I => data_in_frame_1_1
        );

    \I__11865\ : InMux
    port map (
            O => \N__54058\,
            I => \N__54055\
        );

    \I__11864\ : LocalMux
    port map (
            O => \N__54055\,
            I => \N__54051\
        );

    \I__11863\ : InMux
    port map (
            O => \N__54054\,
            I => \N__54048\
        );

    \I__11862\ : Span4Mux_v
    port map (
            O => \N__54051\,
            I => \N__54045\
        );

    \I__11861\ : LocalMux
    port map (
            O => \N__54048\,
            I => \N__54042\
        );

    \I__11860\ : Span4Mux_h
    port map (
            O => \N__54045\,
            I => \N__54039\
        );

    \I__11859\ : Span4Mux_v
    port map (
            O => \N__54042\,
            I => \N__54036\
        );

    \I__11858\ : Odrv4
    port map (
            O => \N__54039\,
            I => \c0.n19970\
        );

    \I__11857\ : Odrv4
    port map (
            O => \N__54036\,
            I => \c0.n19970\
        );

    \I__11856\ : InMux
    port map (
            O => \N__54031\,
            I => \N__54028\
        );

    \I__11855\ : LocalMux
    port map (
            O => \N__54028\,
            I => \N__54025\
        );

    \I__11854\ : Odrv12
    port map (
            O => \N__54025\,
            I => \c0.n6_adj_3501\
        );

    \I__11853\ : CascadeMux
    port map (
            O => \N__54022\,
            I => \N__54017\
        );

    \I__11852\ : InMux
    port map (
            O => \N__54021\,
            I => \N__54014\
        );

    \I__11851\ : CascadeMux
    port map (
            O => \N__54020\,
            I => \N__54011\
        );

    \I__11850\ : InMux
    port map (
            O => \N__54017\,
            I => \N__54008\
        );

    \I__11849\ : LocalMux
    port map (
            O => \N__54014\,
            I => \N__54005\
        );

    \I__11848\ : InMux
    port map (
            O => \N__54011\,
            I => \N__54002\
        );

    \I__11847\ : LocalMux
    port map (
            O => \N__54008\,
            I => \N__53999\
        );

    \I__11846\ : Span4Mux_v
    port map (
            O => \N__54005\,
            I => \N__53996\
        );

    \I__11845\ : LocalMux
    port map (
            O => \N__54002\,
            I => \N__53993\
        );

    \I__11844\ : Odrv12
    port map (
            O => \N__53999\,
            I => \c0.data_in_frame_6_3\
        );

    \I__11843\ : Odrv4
    port map (
            O => \N__53996\,
            I => \c0.data_in_frame_6_3\
        );

    \I__11842\ : Odrv4
    port map (
            O => \N__53993\,
            I => \c0.data_in_frame_6_3\
        );

    \I__11841\ : InMux
    port map (
            O => \N__53986\,
            I => \N__53983\
        );

    \I__11840\ : LocalMux
    port map (
            O => \N__53983\,
            I => \N__53980\
        );

    \I__11839\ : Span4Mux_v
    port map (
            O => \N__53980\,
            I => \N__53977\
        );

    \I__11838\ : Odrv4
    port map (
            O => \N__53977\,
            I => \c0.n25_adj_3048\
        );

    \I__11837\ : InMux
    port map (
            O => \N__53974\,
            I => \N__53970\
        );

    \I__11836\ : InMux
    port map (
            O => \N__53973\,
            I => \N__53967\
        );

    \I__11835\ : LocalMux
    port map (
            O => \N__53970\,
            I => \N__53964\
        );

    \I__11834\ : LocalMux
    port map (
            O => \N__53967\,
            I => \N__53960\
        );

    \I__11833\ : Span4Mux_v
    port map (
            O => \N__53964\,
            I => \N__53957\
        );

    \I__11832\ : InMux
    port map (
            O => \N__53963\,
            I => \N__53954\
        );

    \I__11831\ : Odrv4
    port map (
            O => \N__53960\,
            I => \c0.n19312\
        );

    \I__11830\ : Odrv4
    port map (
            O => \N__53957\,
            I => \c0.n19312\
        );

    \I__11829\ : LocalMux
    port map (
            O => \N__53954\,
            I => \c0.n19312\
        );

    \I__11828\ : InMux
    port map (
            O => \N__53947\,
            I => \N__53944\
        );

    \I__11827\ : LocalMux
    port map (
            O => \N__53944\,
            I => \N__53939\
        );

    \I__11826\ : InMux
    port map (
            O => \N__53943\,
            I => \N__53936\
        );

    \I__11825\ : InMux
    port map (
            O => \N__53942\,
            I => \N__53933\
        );

    \I__11824\ : Span4Mux_h
    port map (
            O => \N__53939\,
            I => \N__53930\
        );

    \I__11823\ : LocalMux
    port map (
            O => \N__53936\,
            I => \N__53927\
        );

    \I__11822\ : LocalMux
    port map (
            O => \N__53933\,
            I => \N__53924\
        );

    \I__11821\ : Span4Mux_v
    port map (
            O => \N__53930\,
            I => \N__53921\
        );

    \I__11820\ : Span4Mux_h
    port map (
            O => \N__53927\,
            I => \N__53918\
        );

    \I__11819\ : Odrv12
    port map (
            O => \N__53924\,
            I => \c0.n20512\
        );

    \I__11818\ : Odrv4
    port map (
            O => \N__53921\,
            I => \c0.n20512\
        );

    \I__11817\ : Odrv4
    port map (
            O => \N__53918\,
            I => \c0.n20512\
        );

    \I__11816\ : InMux
    port map (
            O => \N__53911\,
            I => \N__53908\
        );

    \I__11815\ : LocalMux
    port map (
            O => \N__53908\,
            I => \N__53904\
        );

    \I__11814\ : InMux
    port map (
            O => \N__53907\,
            I => \N__53901\
        );

    \I__11813\ : Span4Mux_v
    port map (
            O => \N__53904\,
            I => \N__53898\
        );

    \I__11812\ : LocalMux
    port map (
            O => \N__53901\,
            I => \N__53895\
        );

    \I__11811\ : Span4Mux_v
    port map (
            O => \N__53898\,
            I => \N__53892\
        );

    \I__11810\ : Span4Mux_v
    port map (
            O => \N__53895\,
            I => \N__53889\
        );

    \I__11809\ : Odrv4
    port map (
            O => \N__53892\,
            I => \c0.n19202\
        );

    \I__11808\ : Odrv4
    port map (
            O => \N__53889\,
            I => \c0.n19202\
        );

    \I__11807\ : CascadeMux
    port map (
            O => \N__53884\,
            I => \c0.n12_adj_3210_cascade_\
        );

    \I__11806\ : InMux
    port map (
            O => \N__53881\,
            I => \N__53878\
        );

    \I__11805\ : LocalMux
    port map (
            O => \N__53878\,
            I => \N__53875\
        );

    \I__11804\ : Span4Mux_h
    port map (
            O => \N__53875\,
            I => \N__53871\
        );

    \I__11803\ : InMux
    port map (
            O => \N__53874\,
            I => \N__53865\
        );

    \I__11802\ : Span4Mux_v
    port map (
            O => \N__53871\,
            I => \N__53862\
        );

    \I__11801\ : InMux
    port map (
            O => \N__53870\,
            I => \N__53859\
        );

    \I__11800\ : InMux
    port map (
            O => \N__53869\,
            I => \N__53854\
        );

    \I__11799\ : InMux
    port map (
            O => \N__53868\,
            I => \N__53854\
        );

    \I__11798\ : LocalMux
    port map (
            O => \N__53865\,
            I => \N__53851\
        );

    \I__11797\ : Odrv4
    port map (
            O => \N__53862\,
            I => \c0.n18433\
        );

    \I__11796\ : LocalMux
    port map (
            O => \N__53859\,
            I => \c0.n18433\
        );

    \I__11795\ : LocalMux
    port map (
            O => \N__53854\,
            I => \c0.n18433\
        );

    \I__11794\ : Odrv4
    port map (
            O => \N__53851\,
            I => \c0.n18433\
        );

    \I__11793\ : InMux
    port map (
            O => \N__53842\,
            I => \N__53839\
        );

    \I__11792\ : LocalMux
    port map (
            O => \N__53839\,
            I => \N__53834\
        );

    \I__11791\ : InMux
    port map (
            O => \N__53838\,
            I => \N__53829\
        );

    \I__11790\ : InMux
    port map (
            O => \N__53837\,
            I => \N__53829\
        );

    \I__11789\ : Odrv4
    port map (
            O => \N__53834\,
            I => \c0.n17834\
        );

    \I__11788\ : LocalMux
    port map (
            O => \N__53829\,
            I => \c0.n17834\
        );

    \I__11787\ : CascadeMux
    port map (
            O => \N__53824\,
            I => \N__53821\
        );

    \I__11786\ : InMux
    port map (
            O => \N__53821\,
            I => \N__53818\
        );

    \I__11785\ : LocalMux
    port map (
            O => \N__53818\,
            I => \N__53815\
        );

    \I__11784\ : Span4Mux_h
    port map (
            O => \N__53815\,
            I => \N__53812\
        );

    \I__11783\ : Odrv4
    port map (
            O => \N__53812\,
            I => \c0.n21767\
        );

    \I__11782\ : InMux
    port map (
            O => \N__53809\,
            I => \N__53805\
        );

    \I__11781\ : InMux
    port map (
            O => \N__53808\,
            I => \N__53801\
        );

    \I__11780\ : LocalMux
    port map (
            O => \N__53805\,
            I => \N__53798\
        );

    \I__11779\ : InMux
    port map (
            O => \N__53804\,
            I => \N__53795\
        );

    \I__11778\ : LocalMux
    port map (
            O => \N__53801\,
            I => \N__53791\
        );

    \I__11777\ : Span4Mux_v
    port map (
            O => \N__53798\,
            I => \N__53786\
        );

    \I__11776\ : LocalMux
    port map (
            O => \N__53795\,
            I => \N__53786\
        );

    \I__11775\ : InMux
    port map (
            O => \N__53794\,
            I => \N__53783\
        );

    \I__11774\ : Span12Mux_v
    port map (
            O => \N__53791\,
            I => \N__53780\
        );

    \I__11773\ : Span4Mux_v
    port map (
            O => \N__53786\,
            I => \N__53777\
        );

    \I__11772\ : LocalMux
    port map (
            O => \N__53783\,
            I => data_in_frame_22_6
        );

    \I__11771\ : Odrv12
    port map (
            O => \N__53780\,
            I => data_in_frame_22_6
        );

    \I__11770\ : Odrv4
    port map (
            O => \N__53777\,
            I => data_in_frame_22_6
        );

    \I__11769\ : InMux
    port map (
            O => \N__53770\,
            I => \N__53765\
        );

    \I__11768\ : InMux
    port map (
            O => \N__53769\,
            I => \N__53760\
        );

    \I__11767\ : InMux
    port map (
            O => \N__53768\,
            I => \N__53760\
        );

    \I__11766\ : LocalMux
    port map (
            O => \N__53765\,
            I => data_in_frame_23_0
        );

    \I__11765\ : LocalMux
    port map (
            O => \N__53760\,
            I => data_in_frame_23_0
        );

    \I__11764\ : InMux
    port map (
            O => \N__53755\,
            I => \N__53752\
        );

    \I__11763\ : LocalMux
    port map (
            O => \N__53752\,
            I => \N__53748\
        );

    \I__11762\ : InMux
    port map (
            O => \N__53751\,
            I => \N__53745\
        );

    \I__11761\ : Span4Mux_v
    port map (
            O => \N__53748\,
            I => \N__53741\
        );

    \I__11760\ : LocalMux
    port map (
            O => \N__53745\,
            I => \N__53738\
        );

    \I__11759\ : InMux
    port map (
            O => \N__53744\,
            I => \N__53735\
        );

    \I__11758\ : Span4Mux_h
    port map (
            O => \N__53741\,
            I => \N__53732\
        );

    \I__11757\ : Span4Mux_v
    port map (
            O => \N__53738\,
            I => \N__53729\
        );

    \I__11756\ : LocalMux
    port map (
            O => \N__53735\,
            I => data_in_frame_23_4
        );

    \I__11755\ : Odrv4
    port map (
            O => \N__53732\,
            I => data_in_frame_23_4
        );

    \I__11754\ : Odrv4
    port map (
            O => \N__53729\,
            I => data_in_frame_23_4
        );

    \I__11753\ : InMux
    port map (
            O => \N__53722\,
            I => \N__53715\
        );

    \I__11752\ : InMux
    port map (
            O => \N__53721\,
            I => \N__53715\
        );

    \I__11751\ : InMux
    port map (
            O => \N__53720\,
            I => \N__53711\
        );

    \I__11750\ : LocalMux
    port map (
            O => \N__53715\,
            I => \N__53706\
        );

    \I__11749\ : InMux
    port map (
            O => \N__53714\,
            I => \N__53703\
        );

    \I__11748\ : LocalMux
    port map (
            O => \N__53711\,
            I => \N__53699\
        );

    \I__11747\ : InMux
    port map (
            O => \N__53710\,
            I => \N__53694\
        );

    \I__11746\ : InMux
    port map (
            O => \N__53709\,
            I => \N__53694\
        );

    \I__11745\ : Span4Mux_v
    port map (
            O => \N__53706\,
            I => \N__53688\
        );

    \I__11744\ : LocalMux
    port map (
            O => \N__53703\,
            I => \N__53688\
        );

    \I__11743\ : InMux
    port map (
            O => \N__53702\,
            I => \N__53685\
        );

    \I__11742\ : Span12Mux_v
    port map (
            O => \N__53699\,
            I => \N__53682\
        );

    \I__11741\ : LocalMux
    port map (
            O => \N__53694\,
            I => \N__53679\
        );

    \I__11740\ : InMux
    port map (
            O => \N__53693\,
            I => \N__53676\
        );

    \I__11739\ : Span4Mux_h
    port map (
            O => \N__53688\,
            I => \N__53671\
        );

    \I__11738\ : LocalMux
    port map (
            O => \N__53685\,
            I => \N__53671\
        );

    \I__11737\ : Odrv12
    port map (
            O => \N__53682\,
            I => n19126
        );

    \I__11736\ : Odrv12
    port map (
            O => \N__53679\,
            I => n19126
        );

    \I__11735\ : LocalMux
    port map (
            O => \N__53676\,
            I => n19126
        );

    \I__11734\ : Odrv4
    port map (
            O => \N__53671\,
            I => n19126
        );

    \I__11733\ : CascadeMux
    port map (
            O => \N__53662\,
            I => \N__53659\
        );

    \I__11732\ : InMux
    port map (
            O => \N__53659\,
            I => \N__53654\
        );

    \I__11731\ : CascadeMux
    port map (
            O => \N__53658\,
            I => \N__53651\
        );

    \I__11730\ : CascadeMux
    port map (
            O => \N__53657\,
            I => \N__53648\
        );

    \I__11729\ : LocalMux
    port map (
            O => \N__53654\,
            I => \N__53645\
        );

    \I__11728\ : InMux
    port map (
            O => \N__53651\,
            I => \N__53642\
        );

    \I__11727\ : InMux
    port map (
            O => \N__53648\,
            I => \N__53639\
        );

    \I__11726\ : Span4Mux_h
    port map (
            O => \N__53645\,
            I => \N__53636\
        );

    \I__11725\ : LocalMux
    port map (
            O => \N__53642\,
            I => \N__53633\
        );

    \I__11724\ : LocalMux
    port map (
            O => \N__53639\,
            I => \c0.data_in_frame_11_0\
        );

    \I__11723\ : Odrv4
    port map (
            O => \N__53636\,
            I => \c0.data_in_frame_11_0\
        );

    \I__11722\ : Odrv4
    port map (
            O => \N__53633\,
            I => \c0.data_in_frame_11_0\
        );

    \I__11721\ : InMux
    port map (
            O => \N__53626\,
            I => \N__53623\
        );

    \I__11720\ : LocalMux
    port map (
            O => \N__53623\,
            I => \N__53619\
        );

    \I__11719\ : InMux
    port map (
            O => \N__53622\,
            I => \N__53615\
        );

    \I__11718\ : Span4Mux_v
    port map (
            O => \N__53619\,
            I => \N__53612\
        );

    \I__11717\ : InMux
    port map (
            O => \N__53618\,
            I => \N__53609\
        );

    \I__11716\ : LocalMux
    port map (
            O => \N__53615\,
            I => data_in_frame_24_7
        );

    \I__11715\ : Odrv4
    port map (
            O => \N__53612\,
            I => data_in_frame_24_7
        );

    \I__11714\ : LocalMux
    port map (
            O => \N__53609\,
            I => data_in_frame_24_7
        );

    \I__11713\ : InMux
    port map (
            O => \N__53602\,
            I => \N__53598\
        );

    \I__11712\ : InMux
    port map (
            O => \N__53601\,
            I => \N__53595\
        );

    \I__11711\ : LocalMux
    port map (
            O => \N__53598\,
            I => \N__53592\
        );

    \I__11710\ : LocalMux
    port map (
            O => \N__53595\,
            I => \c0.n12206\
        );

    \I__11709\ : Odrv4
    port map (
            O => \N__53592\,
            I => \c0.n12206\
        );

    \I__11708\ : InMux
    port map (
            O => \N__53587\,
            I => \N__53582\
        );

    \I__11707\ : InMux
    port map (
            O => \N__53586\,
            I => \N__53579\
        );

    \I__11706\ : InMux
    port map (
            O => \N__53585\,
            I => \N__53576\
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__53582\,
            I => \N__53573\
        );

    \I__11704\ : LocalMux
    port map (
            O => \N__53579\,
            I => \N__53570\
        );

    \I__11703\ : LocalMux
    port map (
            O => \N__53576\,
            I => \c0.n19268\
        );

    \I__11702\ : Odrv4
    port map (
            O => \N__53573\,
            I => \c0.n19268\
        );

    \I__11701\ : Odrv12
    port map (
            O => \N__53570\,
            I => \c0.n19268\
        );

    \I__11700\ : CascadeMux
    port map (
            O => \N__53563\,
            I => \c0.n19268_cascade_\
        );

    \I__11699\ : InMux
    port map (
            O => \N__53560\,
            I => \N__53557\
        );

    \I__11698\ : LocalMux
    port map (
            O => \N__53557\,
            I => \N__53553\
        );

    \I__11697\ : InMux
    port map (
            O => \N__53556\,
            I => \N__53550\
        );

    \I__11696\ : Span4Mux_v
    port map (
            O => \N__53553\,
            I => \N__53545\
        );

    \I__11695\ : LocalMux
    port map (
            O => \N__53550\,
            I => \N__53545\
        );

    \I__11694\ : Span4Mux_h
    port map (
            O => \N__53545\,
            I => \N__53542\
        );

    \I__11693\ : Odrv4
    port map (
            O => \N__53542\,
            I => \c0.n20_adj_3301\
        );

    \I__11692\ : InMux
    port map (
            O => \N__53539\,
            I => \N__53532\
        );

    \I__11691\ : InMux
    port map (
            O => \N__53538\,
            I => \N__53532\
        );

    \I__11690\ : InMux
    port map (
            O => \N__53537\,
            I => \N__53529\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__53532\,
            I => \N__53526\
        );

    \I__11688\ : LocalMux
    port map (
            O => \N__53529\,
            I => \N__53523\
        );

    \I__11687\ : Span4Mux_v
    port map (
            O => \N__53526\,
            I => \N__53520\
        );

    \I__11686\ : Span4Mux_v
    port map (
            O => \N__53523\,
            I => \N__53517\
        );

    \I__11685\ : Odrv4
    port map (
            O => \N__53520\,
            I => \c0.n7_adj_3054\
        );

    \I__11684\ : Odrv4
    port map (
            O => \N__53517\,
            I => \c0.n7_adj_3054\
        );

    \I__11683\ : InMux
    port map (
            O => \N__53512\,
            I => \N__53507\
        );

    \I__11682\ : InMux
    port map (
            O => \N__53511\,
            I => \N__53501\
        );

    \I__11681\ : InMux
    port map (
            O => \N__53510\,
            I => \N__53501\
        );

    \I__11680\ : LocalMux
    port map (
            O => \N__53507\,
            I => \N__53498\
        );

    \I__11679\ : InMux
    port map (
            O => \N__53506\,
            I => \N__53495\
        );

    \I__11678\ : LocalMux
    port map (
            O => \N__53501\,
            I => \N__53491\
        );

    \I__11677\ : Span4Mux_v
    port map (
            O => \N__53498\,
            I => \N__53488\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__53495\,
            I => \N__53485\
        );

    \I__11675\ : InMux
    port map (
            O => \N__53494\,
            I => \N__53482\
        );

    \I__11674\ : Odrv4
    port map (
            O => \N__53491\,
            I => \c0.n11601\
        );

    \I__11673\ : Odrv4
    port map (
            O => \N__53488\,
            I => \c0.n11601\
        );

    \I__11672\ : Odrv4
    port map (
            O => \N__53485\,
            I => \c0.n11601\
        );

    \I__11671\ : LocalMux
    port map (
            O => \N__53482\,
            I => \c0.n11601\
        );

    \I__11670\ : InMux
    port map (
            O => \N__53473\,
            I => \N__53470\
        );

    \I__11669\ : LocalMux
    port map (
            O => \N__53470\,
            I => \N__53466\
        );

    \I__11668\ : InMux
    port map (
            O => \N__53469\,
            I => \N__53463\
        );

    \I__11667\ : Span4Mux_v
    port map (
            O => \N__53466\,
            I => \N__53460\
        );

    \I__11666\ : LocalMux
    port map (
            O => \N__53463\,
            I => \N__53456\
        );

    \I__11665\ : Span4Mux_h
    port map (
            O => \N__53460\,
            I => \N__53453\
        );

    \I__11664\ : InMux
    port map (
            O => \N__53459\,
            I => \N__53450\
        );

    \I__11663\ : Odrv12
    port map (
            O => \N__53456\,
            I => \c0.n19764\
        );

    \I__11662\ : Odrv4
    port map (
            O => \N__53453\,
            I => \c0.n19764\
        );

    \I__11661\ : LocalMux
    port map (
            O => \N__53450\,
            I => \c0.n19764\
        );

    \I__11660\ : InMux
    port map (
            O => \N__53443\,
            I => \N__53439\
        );

    \I__11659\ : InMux
    port map (
            O => \N__53442\,
            I => \N__53436\
        );

    \I__11658\ : LocalMux
    port map (
            O => \N__53439\,
            I => \N__53433\
        );

    \I__11657\ : LocalMux
    port map (
            O => \N__53436\,
            I => \N__53430\
        );

    \I__11656\ : Odrv4
    port map (
            O => \N__53433\,
            I => \c0.n42_adj_3055\
        );

    \I__11655\ : Odrv12
    port map (
            O => \N__53430\,
            I => \c0.n42_adj_3055\
        );

    \I__11654\ : InMux
    port map (
            O => \N__53425\,
            I => \N__53422\
        );

    \I__11653\ : LocalMux
    port map (
            O => \N__53422\,
            I => \N__53418\
        );

    \I__11652\ : InMux
    port map (
            O => \N__53421\,
            I => \N__53415\
        );

    \I__11651\ : Span4Mux_v
    port map (
            O => \N__53418\,
            I => \N__53409\
        );

    \I__11650\ : LocalMux
    port map (
            O => \N__53415\,
            I => \N__53409\
        );

    \I__11649\ : InMux
    port map (
            O => \N__53414\,
            I => \N__53406\
        );

    \I__11648\ : Span4Mux_v
    port map (
            O => \N__53409\,
            I => \N__53403\
        );

    \I__11647\ : LocalMux
    port map (
            O => \N__53406\,
            I => \N__53400\
        );

    \I__11646\ : Odrv4
    port map (
            O => \N__53403\,
            I => \c0.n11815\
        );

    \I__11645\ : Odrv4
    port map (
            O => \N__53400\,
            I => \c0.n11815\
        );

    \I__11644\ : CascadeMux
    port map (
            O => \N__53395\,
            I => \N__53392\
        );

    \I__11643\ : InMux
    port map (
            O => \N__53392\,
            I => \N__53386\
        );

    \I__11642\ : InMux
    port map (
            O => \N__53391\,
            I => \N__53386\
        );

    \I__11641\ : LocalMux
    port map (
            O => \N__53386\,
            I => \c0.n4_adj_3100\
        );

    \I__11640\ : InMux
    port map (
            O => \N__53383\,
            I => \N__53380\
        );

    \I__11639\ : LocalMux
    port map (
            O => \N__53380\,
            I => \N__53376\
        );

    \I__11638\ : CascadeMux
    port map (
            O => \N__53379\,
            I => \N__53372\
        );

    \I__11637\ : Span4Mux_v
    port map (
            O => \N__53376\,
            I => \N__53369\
        );

    \I__11636\ : InMux
    port map (
            O => \N__53375\,
            I => \N__53366\
        );

    \I__11635\ : InMux
    port map (
            O => \N__53372\,
            I => \N__53363\
        );

    \I__11634\ : Sp12to4
    port map (
            O => \N__53369\,
            I => \N__53358\
        );

    \I__11633\ : LocalMux
    port map (
            O => \N__53366\,
            I => \N__53358\
        );

    \I__11632\ : LocalMux
    port map (
            O => \N__53363\,
            I => \c0.data_in_frame_25_0\
        );

    \I__11631\ : Odrv12
    port map (
            O => \N__53358\,
            I => \c0.data_in_frame_25_0\
        );

    \I__11630\ : InMux
    port map (
            O => \N__53353\,
            I => \N__53350\
        );

    \I__11629\ : LocalMux
    port map (
            O => \N__53350\,
            I => \N__53347\
        );

    \I__11628\ : Odrv4
    port map (
            O => \N__53347\,
            I => \c0.n19436\
        );

    \I__11627\ : InMux
    port map (
            O => \N__53344\,
            I => \N__53339\
        );

    \I__11626\ : InMux
    port map (
            O => \N__53343\,
            I => \N__53334\
        );

    \I__11625\ : InMux
    port map (
            O => \N__53342\,
            I => \N__53334\
        );

    \I__11624\ : LocalMux
    port map (
            O => \N__53339\,
            I => \N__53330\
        );

    \I__11623\ : LocalMux
    port map (
            O => \N__53334\,
            I => \N__53327\
        );

    \I__11622\ : InMux
    port map (
            O => \N__53333\,
            I => \N__53322\
        );

    \I__11621\ : Span4Mux_v
    port map (
            O => \N__53330\,
            I => \N__53319\
        );

    \I__11620\ : Span4Mux_h
    port map (
            O => \N__53327\,
            I => \N__53316\
        );

    \I__11619\ : InMux
    port map (
            O => \N__53326\,
            I => \N__53311\
        );

    \I__11618\ : InMux
    port map (
            O => \N__53325\,
            I => \N__53311\
        );

    \I__11617\ : LocalMux
    port map (
            O => \N__53322\,
            I => data_in_frame_22_4
        );

    \I__11616\ : Odrv4
    port map (
            O => \N__53319\,
            I => data_in_frame_22_4
        );

    \I__11615\ : Odrv4
    port map (
            O => \N__53316\,
            I => data_in_frame_22_4
        );

    \I__11614\ : LocalMux
    port map (
            O => \N__53311\,
            I => data_in_frame_22_4
        );

    \I__11613\ : CascadeMux
    port map (
            O => \N__53302\,
            I => \c0.n19436_cascade_\
        );

    \I__11612\ : InMux
    port map (
            O => \N__53299\,
            I => \N__53294\
        );

    \I__11611\ : InMux
    port map (
            O => \N__53298\,
            I => \N__53289\
        );

    \I__11610\ : InMux
    port map (
            O => \N__53297\,
            I => \N__53289\
        );

    \I__11609\ : LocalMux
    port map (
            O => \N__53294\,
            I => \c0.n11776\
        );

    \I__11608\ : LocalMux
    port map (
            O => \N__53289\,
            I => \c0.n11776\
        );

    \I__11607\ : CascadeMux
    port map (
            O => \N__53284\,
            I => \N__53281\
        );

    \I__11606\ : InMux
    port map (
            O => \N__53281\,
            I => \N__53275\
        );

    \I__11605\ : InMux
    port map (
            O => \N__53280\,
            I => \N__53275\
        );

    \I__11604\ : LocalMux
    port map (
            O => \N__53275\,
            I => \c0.n6_adj_3112\
        );

    \I__11603\ : InMux
    port map (
            O => \N__53272\,
            I => \N__53266\
        );

    \I__11602\ : InMux
    port map (
            O => \N__53271\,
            I => \N__53266\
        );

    \I__11601\ : LocalMux
    port map (
            O => \N__53266\,
            I => \c0.n19151\
        );

    \I__11600\ : InMux
    port map (
            O => \N__53263\,
            I => \N__53260\
        );

    \I__11599\ : LocalMux
    port map (
            O => \N__53260\,
            I => \N__53256\
        );

    \I__11598\ : InMux
    port map (
            O => \N__53259\,
            I => \N__53252\
        );

    \I__11597\ : Span4Mux_h
    port map (
            O => \N__53256\,
            I => \N__53249\
        );

    \I__11596\ : InMux
    port map (
            O => \N__53255\,
            I => \N__53246\
        );

    \I__11595\ : LocalMux
    port map (
            O => \N__53252\,
            I => \N__53243\
        );

    \I__11594\ : Span4Mux_h
    port map (
            O => \N__53249\,
            I => \N__53238\
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__53246\,
            I => \N__53238\
        );

    \I__11592\ : Span12Mux_h
    port map (
            O => \N__53243\,
            I => \N__53235\
        );

    \I__11591\ : Odrv4
    port map (
            O => \N__53238\,
            I => \c0.n20933\
        );

    \I__11590\ : Odrv12
    port map (
            O => \N__53235\,
            I => \c0.n20933\
        );

    \I__11589\ : InMux
    port map (
            O => \N__53230\,
            I => \N__53212\
        );

    \I__11588\ : InMux
    port map (
            O => \N__53229\,
            I => \N__53205\
        );

    \I__11587\ : InMux
    port map (
            O => \N__53228\,
            I => \N__53202\
        );

    \I__11586\ : InMux
    port map (
            O => \N__53227\,
            I => \N__53199\
        );

    \I__11585\ : InMux
    port map (
            O => \N__53226\,
            I => \N__53196\
        );

    \I__11584\ : InMux
    port map (
            O => \N__53225\,
            I => \N__53192\
        );

    \I__11583\ : CascadeMux
    port map (
            O => \N__53224\,
            I => \N__53189\
        );

    \I__11582\ : InMux
    port map (
            O => \N__53223\,
            I => \N__53180\
        );

    \I__11581\ : InMux
    port map (
            O => \N__53222\,
            I => \N__53180\
        );

    \I__11580\ : InMux
    port map (
            O => \N__53221\,
            I => \N__53180\
        );

    \I__11579\ : InMux
    port map (
            O => \N__53220\,
            I => \N__53165\
        );

    \I__11578\ : InMux
    port map (
            O => \N__53219\,
            I => \N__53165\
        );

    \I__11577\ : InMux
    port map (
            O => \N__53218\,
            I => \N__53165\
        );

    \I__11576\ : InMux
    port map (
            O => \N__53217\,
            I => \N__53160\
        );

    \I__11575\ : InMux
    port map (
            O => \N__53216\,
            I => \N__53160\
        );

    \I__11574\ : InMux
    port map (
            O => \N__53215\,
            I => \N__53157\
        );

    \I__11573\ : LocalMux
    port map (
            O => \N__53212\,
            I => \N__53154\
        );

    \I__11572\ : InMux
    port map (
            O => \N__53211\,
            I => \N__53145\
        );

    \I__11571\ : InMux
    port map (
            O => \N__53210\,
            I => \N__53145\
        );

    \I__11570\ : InMux
    port map (
            O => \N__53209\,
            I => \N__53145\
        );

    \I__11569\ : InMux
    port map (
            O => \N__53208\,
            I => \N__53145\
        );

    \I__11568\ : LocalMux
    port map (
            O => \N__53205\,
            I => \N__53136\
        );

    \I__11567\ : LocalMux
    port map (
            O => \N__53202\,
            I => \N__53136\
        );

    \I__11566\ : LocalMux
    port map (
            O => \N__53199\,
            I => \N__53136\
        );

    \I__11565\ : LocalMux
    port map (
            O => \N__53196\,
            I => \N__53136\
        );

    \I__11564\ : InMux
    port map (
            O => \N__53195\,
            I => \N__53132\
        );

    \I__11563\ : LocalMux
    port map (
            O => \N__53192\,
            I => \N__53129\
        );

    \I__11562\ : InMux
    port map (
            O => \N__53189\,
            I => \N__53122\
        );

    \I__11561\ : InMux
    port map (
            O => \N__53188\,
            I => \N__53122\
        );

    \I__11560\ : InMux
    port map (
            O => \N__53187\,
            I => \N__53122\
        );

    \I__11559\ : LocalMux
    port map (
            O => \N__53180\,
            I => \N__53119\
        );

    \I__11558\ : InMux
    port map (
            O => \N__53179\,
            I => \N__53115\
        );

    \I__11557\ : InMux
    port map (
            O => \N__53178\,
            I => \N__53112\
        );

    \I__11556\ : InMux
    port map (
            O => \N__53177\,
            I => \N__53109\
        );

    \I__11555\ : InMux
    port map (
            O => \N__53176\,
            I => \N__53106\
        );

    \I__11554\ : InMux
    port map (
            O => \N__53175\,
            I => \N__53103\
        );

    \I__11553\ : InMux
    port map (
            O => \N__53174\,
            I => \N__53100\
        );

    \I__11552\ : InMux
    port map (
            O => \N__53173\,
            I => \N__53095\
        );

    \I__11551\ : InMux
    port map (
            O => \N__53172\,
            I => \N__53095\
        );

    \I__11550\ : LocalMux
    port map (
            O => \N__53165\,
            I => \N__53092\
        );

    \I__11549\ : LocalMux
    port map (
            O => \N__53160\,
            I => \N__53087\
        );

    \I__11548\ : LocalMux
    port map (
            O => \N__53157\,
            I => \N__53087\
        );

    \I__11547\ : Span4Mux_h
    port map (
            O => \N__53154\,
            I => \N__53080\
        );

    \I__11546\ : LocalMux
    port map (
            O => \N__53145\,
            I => \N__53080\
        );

    \I__11545\ : Span4Mux_v
    port map (
            O => \N__53136\,
            I => \N__53080\
        );

    \I__11544\ : InMux
    port map (
            O => \N__53135\,
            I => \N__53076\
        );

    \I__11543\ : LocalMux
    port map (
            O => \N__53132\,
            I => \N__53071\
        );

    \I__11542\ : Span4Mux_h
    port map (
            O => \N__53129\,
            I => \N__53071\
        );

    \I__11541\ : LocalMux
    port map (
            O => \N__53122\,
            I => \N__53066\
        );

    \I__11540\ : Span4Mux_v
    port map (
            O => \N__53119\,
            I => \N__53066\
        );

    \I__11539\ : CascadeMux
    port map (
            O => \N__53118\,
            I => \N__53063\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__53115\,
            I => \N__53060\
        );

    \I__11537\ : LocalMux
    port map (
            O => \N__53112\,
            I => \N__53055\
        );

    \I__11536\ : LocalMux
    port map (
            O => \N__53109\,
            I => \N__53055\
        );

    \I__11535\ : LocalMux
    port map (
            O => \N__53106\,
            I => \N__53040\
        );

    \I__11534\ : LocalMux
    port map (
            O => \N__53103\,
            I => \N__53040\
        );

    \I__11533\ : LocalMux
    port map (
            O => \N__53100\,
            I => \N__53040\
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__53095\,
            I => \N__53040\
        );

    \I__11531\ : Span4Mux_h
    port map (
            O => \N__53092\,
            I => \N__53040\
        );

    \I__11530\ : Span4Mux_v
    port map (
            O => \N__53087\,
            I => \N__53040\
        );

    \I__11529\ : Span4Mux_h
    port map (
            O => \N__53080\,
            I => \N__53040\
        );

    \I__11528\ : InMux
    port map (
            O => \N__53079\,
            I => \N__53037\
        );

    \I__11527\ : LocalMux
    port map (
            O => \N__53076\,
            I => \N__53033\
        );

    \I__11526\ : Span4Mux_v
    port map (
            O => \N__53071\,
            I => \N__53030\
        );

    \I__11525\ : Span4Mux_v
    port map (
            O => \N__53066\,
            I => \N__53027\
        );

    \I__11524\ : InMux
    port map (
            O => \N__53063\,
            I => \N__53024\
        );

    \I__11523\ : Span4Mux_h
    port map (
            O => \N__53060\,
            I => \N__53015\
        );

    \I__11522\ : Span4Mux_v
    port map (
            O => \N__53055\,
            I => \N__53015\
        );

    \I__11521\ : Span4Mux_v
    port map (
            O => \N__53040\,
            I => \N__53015\
        );

    \I__11520\ : LocalMux
    port map (
            O => \N__53037\,
            I => \N__53015\
        );

    \I__11519\ : CascadeMux
    port map (
            O => \N__53036\,
            I => \N__53012\
        );

    \I__11518\ : Sp12to4
    port map (
            O => \N__53033\,
            I => \N__53008\
        );

    \I__11517\ : Span4Mux_v
    port map (
            O => \N__53030\,
            I => \N__53005\
        );

    \I__11516\ : Span4Mux_v
    port map (
            O => \N__53027\,
            I => \N__53000\
        );

    \I__11515\ : LocalMux
    port map (
            O => \N__53024\,
            I => \N__53000\
        );

    \I__11514\ : Span4Mux_v
    port map (
            O => \N__53015\,
            I => \N__52997\
        );

    \I__11513\ : InMux
    port map (
            O => \N__53012\,
            I => \N__52993\
        );

    \I__11512\ : InMux
    port map (
            O => \N__53011\,
            I => \N__52990\
        );

    \I__11511\ : Span12Mux_v
    port map (
            O => \N__53008\,
            I => \N__52987\
        );

    \I__11510\ : Span4Mux_v
    port map (
            O => \N__53005\,
            I => \N__52984\
        );

    \I__11509\ : Span4Mux_v
    port map (
            O => \N__53000\,
            I => \N__52981\
        );

    \I__11508\ : Span4Mux_v
    port map (
            O => \N__52997\,
            I => \N__52978\
        );

    \I__11507\ : InMux
    port map (
            O => \N__52996\,
            I => \N__52975\
        );

    \I__11506\ : LocalMux
    port map (
            O => \N__52993\,
            I => rx_data_ready
        );

    \I__11505\ : LocalMux
    port map (
            O => \N__52990\,
            I => rx_data_ready
        );

    \I__11504\ : Odrv12
    port map (
            O => \N__52987\,
            I => rx_data_ready
        );

    \I__11503\ : Odrv4
    port map (
            O => \N__52984\,
            I => rx_data_ready
        );

    \I__11502\ : Odrv4
    port map (
            O => \N__52981\,
            I => rx_data_ready
        );

    \I__11501\ : Odrv4
    port map (
            O => \N__52978\,
            I => rx_data_ready
        );

    \I__11500\ : LocalMux
    port map (
            O => \N__52975\,
            I => rx_data_ready
        );

    \I__11499\ : InMux
    port map (
            O => \N__52960\,
            I => \N__52957\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__52957\,
            I => \N__52953\
        );

    \I__11497\ : CascadeMux
    port map (
            O => \N__52956\,
            I => \N__52950\
        );

    \I__11496\ : Span4Mux_h
    port map (
            O => \N__52953\,
            I => \N__52946\
        );

    \I__11495\ : InMux
    port map (
            O => \N__52950\,
            I => \N__52943\
        );

    \I__11494\ : InMux
    port map (
            O => \N__52949\,
            I => \N__52939\
        );

    \I__11493\ : Span4Mux_h
    port map (
            O => \N__52946\,
            I => \N__52936\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__52943\,
            I => \N__52933\
        );

    \I__11491\ : InMux
    port map (
            O => \N__52942\,
            I => \N__52930\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__52939\,
            I => data_in_3_6
        );

    \I__11489\ : Odrv4
    port map (
            O => \N__52936\,
            I => data_in_3_6
        );

    \I__11488\ : Odrv4
    port map (
            O => \N__52933\,
            I => data_in_3_6
        );

    \I__11487\ : LocalMux
    port map (
            O => \N__52930\,
            I => data_in_3_6
        );

    \I__11486\ : CascadeMux
    port map (
            O => \N__52921\,
            I => \N__52916\
        );

    \I__11485\ : InMux
    port map (
            O => \N__52920\,
            I => \N__52913\
        );

    \I__11484\ : InMux
    port map (
            O => \N__52919\,
            I => \N__52910\
        );

    \I__11483\ : InMux
    port map (
            O => \N__52916\,
            I => \N__52907\
        );

    \I__11482\ : LocalMux
    port map (
            O => \N__52913\,
            I => \N__52904\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__52910\,
            I => \N__52900\
        );

    \I__11480\ : LocalMux
    port map (
            O => \N__52907\,
            I => \N__52895\
        );

    \I__11479\ : Span4Mux_h
    port map (
            O => \N__52904\,
            I => \N__52895\
        );

    \I__11478\ : InMux
    port map (
            O => \N__52903\,
            I => \N__52892\
        );

    \I__11477\ : Span12Mux_h
    port map (
            O => \N__52900\,
            I => \N__52889\
        );

    \I__11476\ : Span4Mux_h
    port map (
            O => \N__52895\,
            I => \N__52886\
        );

    \I__11475\ : LocalMux
    port map (
            O => \N__52892\,
            I => data_in_2_6
        );

    \I__11474\ : Odrv12
    port map (
            O => \N__52889\,
            I => data_in_2_6
        );

    \I__11473\ : Odrv4
    port map (
            O => \N__52886\,
            I => data_in_2_6
        );

    \I__11472\ : InMux
    port map (
            O => \N__52879\,
            I => \N__52876\
        );

    \I__11471\ : LocalMux
    port map (
            O => \N__52876\,
            I => \N__52872\
        );

    \I__11470\ : InMux
    port map (
            O => \N__52875\,
            I => \N__52869\
        );

    \I__11469\ : Odrv4
    port map (
            O => \N__52872\,
            I => \c0.n24_adj_3427\
        );

    \I__11468\ : LocalMux
    port map (
            O => \N__52869\,
            I => \c0.n24_adj_3427\
        );

    \I__11467\ : InMux
    port map (
            O => \N__52864\,
            I => \N__52859\
        );

    \I__11466\ : InMux
    port map (
            O => \N__52863\,
            I => \N__52854\
        );

    \I__11465\ : InMux
    port map (
            O => \N__52862\,
            I => \N__52854\
        );

    \I__11464\ : LocalMux
    port map (
            O => \N__52859\,
            I => \N__52849\
        );

    \I__11463\ : LocalMux
    port map (
            O => \N__52854\,
            I => \N__52849\
        );

    \I__11462\ : Span4Mux_v
    port map (
            O => \N__52849\,
            I => \N__52846\
        );

    \I__11461\ : Odrv4
    port map (
            O => \N__52846\,
            I => \c0.n11714\
        );

    \I__11460\ : InMux
    port map (
            O => \N__52843\,
            I => \N__52840\
        );

    \I__11459\ : LocalMux
    port map (
            O => \N__52840\,
            I => \N__52837\
        );

    \I__11458\ : Span4Mux_h
    port map (
            O => \N__52837\,
            I => \N__52834\
        );

    \I__11457\ : Odrv4
    port map (
            O => \N__52834\,
            I => \c0.n22_adj_3296\
        );

    \I__11456\ : CascadeMux
    port map (
            O => \N__52831\,
            I => \c0.n19159_cascade_\
        );

    \I__11455\ : InMux
    port map (
            O => \N__52828\,
            I => \N__52824\
        );

    \I__11454\ : InMux
    port map (
            O => \N__52827\,
            I => \N__52821\
        );

    \I__11453\ : LocalMux
    port map (
            O => \N__52824\,
            I => \N__52818\
        );

    \I__11452\ : LocalMux
    port map (
            O => \N__52821\,
            I => \N__52815\
        );

    \I__11451\ : Span4Mux_v
    port map (
            O => \N__52818\,
            I => \N__52812\
        );

    \I__11450\ : Span4Mux_h
    port map (
            O => \N__52815\,
            I => \N__52809\
        );

    \I__11449\ : Odrv4
    port map (
            O => \N__52812\,
            I => \c0.n11632\
        );

    \I__11448\ : Odrv4
    port map (
            O => \N__52809\,
            I => \c0.n11632\
        );

    \I__11447\ : InMux
    port map (
            O => \N__52804\,
            I => \N__52801\
        );

    \I__11446\ : LocalMux
    port map (
            O => \N__52801\,
            I => \c0.n19159\
        );

    \I__11445\ : CascadeMux
    port map (
            O => \N__52798\,
            I => \N__52795\
        );

    \I__11444\ : InMux
    port map (
            O => \N__52795\,
            I => \N__52791\
        );

    \I__11443\ : CascadeMux
    port map (
            O => \N__52794\,
            I => \N__52788\
        );

    \I__11442\ : LocalMux
    port map (
            O => \N__52791\,
            I => \N__52785\
        );

    \I__11441\ : InMux
    port map (
            O => \N__52788\,
            I => \N__52782\
        );

    \I__11440\ : Span4Mux_v
    port map (
            O => \N__52785\,
            I => \N__52779\
        );

    \I__11439\ : LocalMux
    port map (
            O => \N__52782\,
            I => \c0.data_in_frame_28_7\
        );

    \I__11438\ : Odrv4
    port map (
            O => \N__52779\,
            I => \c0.data_in_frame_28_7\
        );

    \I__11437\ : InMux
    port map (
            O => \N__52774\,
            I => \N__52771\
        );

    \I__11436\ : LocalMux
    port map (
            O => \N__52771\,
            I => \N__52768\
        );

    \I__11435\ : Span4Mux_h
    port map (
            O => \N__52768\,
            I => \N__52765\
        );

    \I__11434\ : Odrv4
    port map (
            O => \N__52765\,
            I => \c0.n79\
        );

    \I__11433\ : InMux
    port map (
            O => \N__52762\,
            I => \N__52759\
        );

    \I__11432\ : LocalMux
    port map (
            O => \N__52759\,
            I => \N__52755\
        );

    \I__11431\ : InMux
    port map (
            O => \N__52758\,
            I => \N__52752\
        );

    \I__11430\ : Span12Mux_h
    port map (
            O => \N__52755\,
            I => \N__52749\
        );

    \I__11429\ : LocalMux
    port map (
            O => \N__52752\,
            I => \N__52746\
        );

    \I__11428\ : Span12Mux_v
    port map (
            O => \N__52749\,
            I => \N__52743\
        );

    \I__11427\ : Span4Mux_v
    port map (
            O => \N__52746\,
            I => \N__52740\
        );

    \I__11426\ : Odrv12
    port map (
            O => \N__52743\,
            I => \c0.n10_adj_3207\
        );

    \I__11425\ : Odrv4
    port map (
            O => \N__52740\,
            I => \c0.n10_adj_3207\
        );

    \I__11424\ : InMux
    port map (
            O => \N__52735\,
            I => \N__52729\
        );

    \I__11423\ : InMux
    port map (
            O => \N__52734\,
            I => \N__52729\
        );

    \I__11422\ : LocalMux
    port map (
            O => \N__52729\,
            I => \N__52726\
        );

    \I__11421\ : Span4Mux_v
    port map (
            O => \N__52726\,
            I => \N__52723\
        );

    \I__11420\ : Span4Mux_h
    port map (
            O => \N__52723\,
            I => \N__52719\
        );

    \I__11419\ : InMux
    port map (
            O => \N__52722\,
            I => \N__52716\
        );

    \I__11418\ : Odrv4
    port map (
            O => \N__52719\,
            I => \c0.n11_adj_3206\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__52716\,
            I => \c0.n11_adj_3206\
        );

    \I__11416\ : CascadeMux
    port map (
            O => \N__52711\,
            I => \c0.n11776_cascade_\
        );

    \I__11415\ : InMux
    port map (
            O => \N__52708\,
            I => \N__52703\
        );

    \I__11414\ : InMux
    port map (
            O => \N__52707\,
            I => \N__52698\
        );

    \I__11413\ : InMux
    port map (
            O => \N__52706\,
            I => \N__52698\
        );

    \I__11412\ : LocalMux
    port map (
            O => \N__52703\,
            I => \c0.n6_adj_3319\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__52698\,
            I => \c0.n6_adj_3319\
        );

    \I__11410\ : CascadeMux
    port map (
            O => \N__52693\,
            I => \c0.n70_adj_3087_cascade_\
        );

    \I__11409\ : InMux
    port map (
            O => \N__52690\,
            I => \N__52686\
        );

    \I__11408\ : InMux
    port map (
            O => \N__52689\,
            I => \N__52683\
        );

    \I__11407\ : LocalMux
    port map (
            O => \N__52686\,
            I => \N__52678\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__52683\,
            I => \N__52678\
        );

    \I__11405\ : Span4Mux_v
    port map (
            O => \N__52678\,
            I => \N__52675\
        );

    \I__11404\ : Odrv4
    port map (
            O => \N__52675\,
            I => \c0.n20339\
        );

    \I__11403\ : InMux
    port map (
            O => \N__52672\,
            I => \N__52668\
        );

    \I__11402\ : InMux
    port map (
            O => \N__52671\,
            I => \N__52665\
        );

    \I__11401\ : LocalMux
    port map (
            O => \N__52668\,
            I => \N__52662\
        );

    \I__11400\ : LocalMux
    port map (
            O => \N__52665\,
            I => \N__52657\
        );

    \I__11399\ : Span4Mux_h
    port map (
            O => \N__52662\,
            I => \N__52657\
        );

    \I__11398\ : Span4Mux_h
    port map (
            O => \N__52657\,
            I => \N__52654\
        );

    \I__11397\ : Odrv4
    port map (
            O => \N__52654\,
            I => \c0.n27_adj_3311\
        );

    \I__11396\ : InMux
    port map (
            O => \N__52651\,
            I => \N__52648\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__52648\,
            I => \N__52642\
        );

    \I__11394\ : InMux
    port map (
            O => \N__52647\,
            I => \N__52637\
        );

    \I__11393\ : InMux
    port map (
            O => \N__52646\,
            I => \N__52637\
        );

    \I__11392\ : InMux
    port map (
            O => \N__52645\,
            I => \N__52634\
        );

    \I__11391\ : Span4Mux_v
    port map (
            O => \N__52642\,
            I => \N__52629\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__52637\,
            I => \N__52629\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__52634\,
            I => \N__52626\
        );

    \I__11388\ : Span4Mux_h
    port map (
            O => \N__52629\,
            I => \N__52623\
        );

    \I__11387\ : Span4Mux_v
    port map (
            O => \N__52626\,
            I => \N__52620\
        );

    \I__11386\ : Odrv4
    port map (
            O => \N__52623\,
            I => \c0.n7_adj_3094\
        );

    \I__11385\ : Odrv4
    port map (
            O => \N__52620\,
            I => \c0.n7_adj_3094\
        );

    \I__11384\ : InMux
    port map (
            O => \N__52615\,
            I => \N__52612\
        );

    \I__11383\ : LocalMux
    port map (
            O => \N__52612\,
            I => \N__52609\
        );

    \I__11382\ : Odrv4
    port map (
            O => \N__52609\,
            I => \c0.n20_adj_3293\
        );

    \I__11381\ : InMux
    port map (
            O => \N__52606\,
            I => \N__52603\
        );

    \I__11380\ : LocalMux
    port map (
            O => \N__52603\,
            I => \N__52600\
        );

    \I__11379\ : Span4Mux_h
    port map (
            O => \N__52600\,
            I => \N__52596\
        );

    \I__11378\ : InMux
    port map (
            O => \N__52599\,
            I => \N__52593\
        );

    \I__11377\ : Odrv4
    port map (
            O => \N__52596\,
            I => \c0.n33_adj_3279\
        );

    \I__11376\ : LocalMux
    port map (
            O => \N__52593\,
            I => \c0.n33_adj_3279\
        );

    \I__11375\ : InMux
    port map (
            O => \N__52588\,
            I => \N__52585\
        );

    \I__11374\ : LocalMux
    port map (
            O => \N__52585\,
            I => \c0.n30_adj_3295\
        );

    \I__11373\ : CascadeMux
    port map (
            O => \N__52582\,
            I => \c0.n32_adj_3294_cascade_\
        );

    \I__11372\ : InMux
    port map (
            O => \N__52579\,
            I => \N__52576\
        );

    \I__11371\ : LocalMux
    port map (
            O => \N__52576\,
            I => \N__52573\
        );

    \I__11370\ : Span4Mux_v
    port map (
            O => \N__52573\,
            I => \N__52570\
        );

    \I__11369\ : Odrv4
    port map (
            O => \N__52570\,
            I => \c0.n21075\
        );

    \I__11368\ : InMux
    port map (
            O => \N__52567\,
            I => \N__52564\
        );

    \I__11367\ : LocalMux
    port map (
            O => \N__52564\,
            I => \N__52560\
        );

    \I__11366\ : InMux
    port map (
            O => \N__52563\,
            I => \N__52556\
        );

    \I__11365\ : Span4Mux_h
    port map (
            O => \N__52560\,
            I => \N__52553\
        );

    \I__11364\ : InMux
    port map (
            O => \N__52559\,
            I => \N__52550\
        );

    \I__11363\ : LocalMux
    port map (
            O => \N__52556\,
            I => \N__52547\
        );

    \I__11362\ : Span4Mux_v
    port map (
            O => \N__52553\,
            I => \N__52544\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__52550\,
            I => \N__52540\
        );

    \I__11360\ : Span4Mux_v
    port map (
            O => \N__52547\,
            I => \N__52535\
        );

    \I__11359\ : Span4Mux_h
    port map (
            O => \N__52544\,
            I => \N__52535\
        );

    \I__11358\ : InMux
    port map (
            O => \N__52543\,
            I => \N__52532\
        );

    \I__11357\ : Odrv4
    port map (
            O => \N__52540\,
            I => \c0.n7_adj_3079\
        );

    \I__11356\ : Odrv4
    port map (
            O => \N__52535\,
            I => \c0.n7_adj_3079\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__52532\,
            I => \c0.n7_adj_3079\
        );

    \I__11354\ : InMux
    port map (
            O => \N__52525\,
            I => \N__52522\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__52522\,
            I => \c0.n29_adj_3299\
        );

    \I__11352\ : InMux
    port map (
            O => \N__52519\,
            I => \N__52516\
        );

    \I__11351\ : LocalMux
    port map (
            O => \N__52516\,
            I => \N__52513\
        );

    \I__11350\ : Span4Mux_v
    port map (
            O => \N__52513\,
            I => \N__52510\
        );

    \I__11349\ : Odrv4
    port map (
            O => \N__52510\,
            I => \c0.n19_adj_3320\
        );

    \I__11348\ : InMux
    port map (
            O => \N__52507\,
            I => \N__52500\
        );

    \I__11347\ : InMux
    port map (
            O => \N__52506\,
            I => \N__52500\
        );

    \I__11346\ : InMux
    port map (
            O => \N__52505\,
            I => \N__52497\
        );

    \I__11345\ : LocalMux
    port map (
            O => \N__52500\,
            I => \c0.n20336\
        );

    \I__11344\ : LocalMux
    port map (
            O => \N__52497\,
            I => \c0.n20336\
        );

    \I__11343\ : CascadeMux
    port map (
            O => \N__52492\,
            I => \N__52486\
        );

    \I__11342\ : InMux
    port map (
            O => \N__52491\,
            I => \N__52483\
        );

    \I__11341\ : CascadeMux
    port map (
            O => \N__52490\,
            I => \N__52479\
        );

    \I__11340\ : CascadeMux
    port map (
            O => \N__52489\,
            I => \N__52476\
        );

    \I__11339\ : InMux
    port map (
            O => \N__52486\,
            I => \N__52473\
        );

    \I__11338\ : LocalMux
    port map (
            O => \N__52483\,
            I => \N__52470\
        );

    \I__11337\ : InMux
    port map (
            O => \N__52482\,
            I => \N__52467\
        );

    \I__11336\ : InMux
    port map (
            O => \N__52479\,
            I => \N__52462\
        );

    \I__11335\ : InMux
    port map (
            O => \N__52476\,
            I => \N__52462\
        );

    \I__11334\ : LocalMux
    port map (
            O => \N__52473\,
            I => \N__52459\
        );

    \I__11333\ : Span4Mux_h
    port map (
            O => \N__52470\,
            I => \N__52454\
        );

    \I__11332\ : LocalMux
    port map (
            O => \N__52467\,
            I => \N__52454\
        );

    \I__11331\ : LocalMux
    port map (
            O => \N__52462\,
            I => \c0.n18379\
        );

    \I__11330\ : Odrv4
    port map (
            O => \N__52459\,
            I => \c0.n18379\
        );

    \I__11329\ : Odrv4
    port map (
            O => \N__52454\,
            I => \c0.n18379\
        );

    \I__11328\ : InMux
    port map (
            O => \N__52447\,
            I => \N__52441\
        );

    \I__11327\ : InMux
    port map (
            O => \N__52446\,
            I => \N__52438\
        );

    \I__11326\ : InMux
    port map (
            O => \N__52445\,
            I => \N__52435\
        );

    \I__11325\ : InMux
    port map (
            O => \N__52444\,
            I => \N__52432\
        );

    \I__11324\ : LocalMux
    port map (
            O => \N__52441\,
            I => \c0.n21034\
        );

    \I__11323\ : LocalMux
    port map (
            O => \N__52438\,
            I => \c0.n21034\
        );

    \I__11322\ : LocalMux
    port map (
            O => \N__52435\,
            I => \c0.n21034\
        );

    \I__11321\ : LocalMux
    port map (
            O => \N__52432\,
            I => \c0.n21034\
        );

    \I__11320\ : InMux
    port map (
            O => \N__52423\,
            I => \N__52420\
        );

    \I__11319\ : LocalMux
    port map (
            O => \N__52420\,
            I => \N__52417\
        );

    \I__11318\ : Span4Mux_h
    port map (
            O => \N__52417\,
            I => \N__52413\
        );

    \I__11317\ : InMux
    port map (
            O => \N__52416\,
            I => \N__52410\
        );

    \I__11316\ : Odrv4
    port map (
            O => \N__52413\,
            I => \c0.n57\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__52410\,
            I => \c0.n57\
        );

    \I__11314\ : InMux
    port map (
            O => \N__52405\,
            I => \N__52402\
        );

    \I__11313\ : LocalMux
    port map (
            O => \N__52402\,
            I => \c0.n32_adj_3465\
        );

    \I__11312\ : CascadeMux
    port map (
            O => \N__52399\,
            I => \N__52394\
        );

    \I__11311\ : InMux
    port map (
            O => \N__52398\,
            I => \N__52391\
        );

    \I__11310\ : InMux
    port map (
            O => \N__52397\,
            I => \N__52388\
        );

    \I__11309\ : InMux
    port map (
            O => \N__52394\,
            I => \N__52385\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__52391\,
            I => \c0.n33_adj_3315\
        );

    \I__11307\ : LocalMux
    port map (
            O => \N__52388\,
            I => \c0.n33_adj_3315\
        );

    \I__11306\ : LocalMux
    port map (
            O => \N__52385\,
            I => \c0.n33_adj_3315\
        );

    \I__11305\ : InMux
    port map (
            O => \N__52378\,
            I => \N__52375\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__52375\,
            I => \N__52372\
        );

    \I__11303\ : Span4Mux_h
    port map (
            O => \N__52372\,
            I => \N__52369\
        );

    \I__11302\ : Odrv4
    port map (
            O => \N__52369\,
            I => \c0.n49_adj_3316\
        );

    \I__11301\ : InMux
    port map (
            O => \N__52366\,
            I => \N__52363\
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__52363\,
            I => \N__52359\
        );

    \I__11299\ : InMux
    port map (
            O => \N__52362\,
            I => \N__52356\
        );

    \I__11298\ : Odrv4
    port map (
            O => \N__52359\,
            I => \c0.n35_adj_3317\
        );

    \I__11297\ : LocalMux
    port map (
            O => \N__52356\,
            I => \c0.n35_adj_3317\
        );

    \I__11296\ : InMux
    port map (
            O => \N__52351\,
            I => \N__52347\
        );

    \I__11295\ : InMux
    port map (
            O => \N__52350\,
            I => \N__52342\
        );

    \I__11294\ : LocalMux
    port map (
            O => \N__52347\,
            I => \N__52339\
        );

    \I__11293\ : InMux
    port map (
            O => \N__52346\,
            I => \N__52335\
        );

    \I__11292\ : InMux
    port map (
            O => \N__52345\,
            I => \N__52332\
        );

    \I__11291\ : LocalMux
    port map (
            O => \N__52342\,
            I => \N__52328\
        );

    \I__11290\ : Span4Mux_h
    port map (
            O => \N__52339\,
            I => \N__52325\
        );

    \I__11289\ : InMux
    port map (
            O => \N__52338\,
            I => \N__52322\
        );

    \I__11288\ : LocalMux
    port map (
            O => \N__52335\,
            I => \N__52319\
        );

    \I__11287\ : LocalMux
    port map (
            O => \N__52332\,
            I => \N__52316\
        );

    \I__11286\ : CascadeMux
    port map (
            O => \N__52331\,
            I => \N__52313\
        );

    \I__11285\ : Span4Mux_h
    port map (
            O => \N__52328\,
            I => \N__52308\
        );

    \I__11284\ : Span4Mux_v
    port map (
            O => \N__52325\,
            I => \N__52308\
        );

    \I__11283\ : LocalMux
    port map (
            O => \N__52322\,
            I => \N__52305\
        );

    \I__11282\ : Span4Mux_h
    port map (
            O => \N__52319\,
            I => \N__52300\
        );

    \I__11281\ : Span4Mux_h
    port map (
            O => \N__52316\,
            I => \N__52300\
        );

    \I__11280\ : InMux
    port map (
            O => \N__52313\,
            I => \N__52297\
        );

    \I__11279\ : Span4Mux_v
    port map (
            O => \N__52308\,
            I => \N__52294\
        );

    \I__11278\ : Span4Mux_h
    port map (
            O => \N__52305\,
            I => \N__52289\
        );

    \I__11277\ : Span4Mux_v
    port map (
            O => \N__52300\,
            I => \N__52289\
        );

    \I__11276\ : LocalMux
    port map (
            O => \N__52297\,
            I => \c0.data_in_frame_17_1\
        );

    \I__11275\ : Odrv4
    port map (
            O => \N__52294\,
            I => \c0.data_in_frame_17_1\
        );

    \I__11274\ : Odrv4
    port map (
            O => \N__52289\,
            I => \c0.data_in_frame_17_1\
        );

    \I__11273\ : InMux
    port map (
            O => \N__52282\,
            I => \N__52279\
        );

    \I__11272\ : LocalMux
    port map (
            O => \N__52279\,
            I => \N__52276\
        );

    \I__11271\ : Span4Mux_v
    port map (
            O => \N__52276\,
            I => \N__52272\
        );

    \I__11270\ : InMux
    port map (
            O => \N__52275\,
            I => \N__52269\
        );

    \I__11269\ : Span4Mux_h
    port map (
            O => \N__52272\,
            I => \N__52264\
        );

    \I__11268\ : LocalMux
    port map (
            O => \N__52269\,
            I => \N__52264\
        );

    \I__11267\ : Odrv4
    port map (
            O => \N__52264\,
            I => \c0.n17871\
        );

    \I__11266\ : InMux
    port map (
            O => \N__52261\,
            I => \N__52258\
        );

    \I__11265\ : LocalMux
    port map (
            O => \N__52258\,
            I => \N__52255\
        );

    \I__11264\ : Odrv4
    port map (
            O => \N__52255\,
            I => \c0.n22_adj_3363\
        );

    \I__11263\ : CascadeMux
    port map (
            O => \N__52252\,
            I => \c0.n22_adj_3363_cascade_\
        );

    \I__11262\ : InMux
    port map (
            O => \N__52249\,
            I => \N__52246\
        );

    \I__11261\ : LocalMux
    port map (
            O => \N__52246\,
            I => \N__52243\
        );

    \I__11260\ : Odrv4
    port map (
            O => \N__52243\,
            I => \c0.n30_adj_3468\
        );

    \I__11259\ : InMux
    port map (
            O => \N__52240\,
            I => \N__52237\
        );

    \I__11258\ : LocalMux
    port map (
            O => \N__52237\,
            I => \N__52234\
        );

    \I__11257\ : Odrv12
    port map (
            O => \N__52234\,
            I => \c0.n65\
        );

    \I__11256\ : InMux
    port map (
            O => \N__52231\,
            I => \N__52228\
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__52228\,
            I => \N__52225\
        );

    \I__11254\ : Sp12to4
    port map (
            O => \N__52225\,
            I => \N__52222\
        );

    \I__11253\ : Span12Mux_v
    port map (
            O => \N__52222\,
            I => \N__52219\
        );

    \I__11252\ : Odrv12
    port map (
            O => \N__52219\,
            I => \c0.n19223\
        );

    \I__11251\ : InMux
    port map (
            O => \N__52216\,
            I => \N__52213\
        );

    \I__11250\ : LocalMux
    port map (
            O => \N__52213\,
            I => \N__52210\
        );

    \I__11249\ : Span4Mux_h
    port map (
            O => \N__52210\,
            I => \N__52207\
        );

    \I__11248\ : Span4Mux_v
    port map (
            O => \N__52207\,
            I => \N__52203\
        );

    \I__11247\ : InMux
    port map (
            O => \N__52206\,
            I => \N__52200\
        );

    \I__11246\ : Odrv4
    port map (
            O => \N__52203\,
            I => \c0.n12218\
        );

    \I__11245\ : LocalMux
    port map (
            O => \N__52200\,
            I => \c0.n12218\
        );

    \I__11244\ : CascadeMux
    port map (
            O => \N__52195\,
            I => \c0.n7_adj_3047_cascade_\
        );

    \I__11243\ : CascadeMux
    port map (
            O => \N__52192\,
            I => \c0.n28_adj_3059_cascade_\
        );

    \I__11242\ : InMux
    port map (
            O => \N__52189\,
            I => \N__52186\
        );

    \I__11241\ : LocalMux
    port map (
            O => \N__52186\,
            I => \N__52181\
        );

    \I__11240\ : InMux
    port map (
            O => \N__52185\,
            I => \N__52176\
        );

    \I__11239\ : InMux
    port map (
            O => \N__52184\,
            I => \N__52176\
        );

    \I__11238\ : Odrv4
    port map (
            O => \N__52181\,
            I => \c0.n36_adj_3452\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__52176\,
            I => \c0.n36_adj_3452\
        );

    \I__11236\ : InMux
    port map (
            O => \N__52171\,
            I => \N__52168\
        );

    \I__11235\ : LocalMux
    port map (
            O => \N__52168\,
            I => \N__52163\
        );

    \I__11234\ : InMux
    port map (
            O => \N__52167\,
            I => \N__52160\
        );

    \I__11233\ : InMux
    port map (
            O => \N__52166\,
            I => \N__52155\
        );

    \I__11232\ : Span4Mux_h
    port map (
            O => \N__52163\,
            I => \N__52152\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__52160\,
            I => \N__52149\
        );

    \I__11230\ : InMux
    port map (
            O => \N__52159\,
            I => \N__52144\
        );

    \I__11229\ : InMux
    port map (
            O => \N__52158\,
            I => \N__52144\
        );

    \I__11228\ : LocalMux
    port map (
            O => \N__52155\,
            I => \c0.n47\
        );

    \I__11227\ : Odrv4
    port map (
            O => \N__52152\,
            I => \c0.n47\
        );

    \I__11226\ : Odrv4
    port map (
            O => \N__52149\,
            I => \c0.n47\
        );

    \I__11225\ : LocalMux
    port map (
            O => \N__52144\,
            I => \c0.n47\
        );

    \I__11224\ : InMux
    port map (
            O => \N__52135\,
            I => \N__52131\
        );

    \I__11223\ : InMux
    port map (
            O => \N__52134\,
            I => \N__52127\
        );

    \I__11222\ : LocalMux
    port map (
            O => \N__52131\,
            I => \N__52124\
        );

    \I__11221\ : InMux
    port map (
            O => \N__52130\,
            I => \N__52121\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__52127\,
            I => \N__52118\
        );

    \I__11219\ : Span4Mux_h
    port map (
            O => \N__52124\,
            I => \N__52115\
        );

    \I__11218\ : LocalMux
    port map (
            O => \N__52121\,
            I => \c0.n17819\
        );

    \I__11217\ : Odrv4
    port map (
            O => \N__52118\,
            I => \c0.n17819\
        );

    \I__11216\ : Odrv4
    port map (
            O => \N__52115\,
            I => \c0.n17819\
        );

    \I__11215\ : InMux
    port map (
            O => \N__52108\,
            I => \N__52104\
        );

    \I__11214\ : InMux
    port map (
            O => \N__52107\,
            I => \N__52100\
        );

    \I__11213\ : LocalMux
    port map (
            O => \N__52104\,
            I => \N__52097\
        );

    \I__11212\ : InMux
    port map (
            O => \N__52103\,
            I => \N__52094\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__52100\,
            I => \N__52089\
        );

    \I__11210\ : Span4Mux_h
    port map (
            O => \N__52097\,
            I => \N__52084\
        );

    \I__11209\ : LocalMux
    port map (
            O => \N__52094\,
            I => \N__52084\
        );

    \I__11208\ : InMux
    port map (
            O => \N__52093\,
            I => \N__52081\
        );

    \I__11207\ : InMux
    port map (
            O => \N__52092\,
            I => \N__52078\
        );

    \I__11206\ : Span4Mux_h
    port map (
            O => \N__52089\,
            I => \N__52075\
        );

    \I__11205\ : Span4Mux_v
    port map (
            O => \N__52084\,
            I => \N__52070\
        );

    \I__11204\ : LocalMux
    port map (
            O => \N__52081\,
            I => \N__52070\
        );

    \I__11203\ : LocalMux
    port map (
            O => \N__52078\,
            I => \N__52067\
        );

    \I__11202\ : Odrv4
    port map (
            O => \N__52075\,
            I => \c0.n20321\
        );

    \I__11201\ : Odrv4
    port map (
            O => \N__52070\,
            I => \c0.n20321\
        );

    \I__11200\ : Odrv4
    port map (
            O => \N__52067\,
            I => \c0.n20321\
        );

    \I__11199\ : InMux
    port map (
            O => \N__52060\,
            I => \N__52057\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__52057\,
            I => \c0.n19824\
        );

    \I__11197\ : InMux
    port map (
            O => \N__52054\,
            I => \N__52050\
        );

    \I__11196\ : InMux
    port map (
            O => \N__52053\,
            I => \N__52047\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__52050\,
            I => \N__52044\
        );

    \I__11194\ : LocalMux
    port map (
            O => \N__52047\,
            I => \N__52041\
        );

    \I__11193\ : Span4Mux_v
    port map (
            O => \N__52044\,
            I => \N__52037\
        );

    \I__11192\ : Span4Mux_v
    port map (
            O => \N__52041\,
            I => \N__52034\
        );

    \I__11191\ : InMux
    port map (
            O => \N__52040\,
            I => \N__52031\
        );

    \I__11190\ : Odrv4
    port map (
            O => \N__52037\,
            I => \c0.n12_adj_3469\
        );

    \I__11189\ : Odrv4
    port map (
            O => \N__52034\,
            I => \c0.n12_adj_3469\
        );

    \I__11188\ : LocalMux
    port map (
            O => \N__52031\,
            I => \c0.n12_adj_3469\
        );

    \I__11187\ : CascadeMux
    port map (
            O => \N__52024\,
            I => \c0.n29_adj_3461_cascade_\
        );

    \I__11186\ : InMux
    port map (
            O => \N__52021\,
            I => \N__52016\
        );

    \I__11185\ : InMux
    port map (
            O => \N__52020\,
            I => \N__52012\
        );

    \I__11184\ : InMux
    port map (
            O => \N__52019\,
            I => \N__52009\
        );

    \I__11183\ : LocalMux
    port map (
            O => \N__52016\,
            I => \N__52006\
        );

    \I__11182\ : InMux
    port map (
            O => \N__52015\,
            I => \N__52003\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__52012\,
            I => \N__52000\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__52009\,
            I => \N__51997\
        );

    \I__11179\ : Span4Mux_v
    port map (
            O => \N__52006\,
            I => \N__51992\
        );

    \I__11178\ : LocalMux
    port map (
            O => \N__52003\,
            I => \N__51992\
        );

    \I__11177\ : Span4Mux_v
    port map (
            O => \N__52000\,
            I => \N__51986\
        );

    \I__11176\ : Span4Mux_v
    port map (
            O => \N__51997\,
            I => \N__51986\
        );

    \I__11175\ : Span4Mux_h
    port map (
            O => \N__51992\,
            I => \N__51983\
        );

    \I__11174\ : InMux
    port map (
            O => \N__51991\,
            I => \N__51980\
        );

    \I__11173\ : Odrv4
    port map (
            O => \N__51986\,
            I => \c0.n25_adj_3035\
        );

    \I__11172\ : Odrv4
    port map (
            O => \N__51983\,
            I => \c0.n25_adj_3035\
        );

    \I__11171\ : LocalMux
    port map (
            O => \N__51980\,
            I => \c0.n25_adj_3035\
        );

    \I__11170\ : InMux
    port map (
            O => \N__51973\,
            I => \N__51969\
        );

    \I__11169\ : InMux
    port map (
            O => \N__51972\,
            I => \N__51966\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__51969\,
            I => \N__51963\
        );

    \I__11167\ : LocalMux
    port map (
            O => \N__51966\,
            I => \N__51960\
        );

    \I__11166\ : Sp12to4
    port map (
            O => \N__51963\,
            I => \N__51957\
        );

    \I__11165\ : Span4Mux_v
    port map (
            O => \N__51960\,
            I => \N__51954\
        );

    \I__11164\ : Span12Mux_h
    port map (
            O => \N__51957\,
            I => \N__51951\
        );

    \I__11163\ : Odrv4
    port map (
            O => \N__51954\,
            I => \c0.n23_adj_3364\
        );

    \I__11162\ : Odrv12
    port map (
            O => \N__51951\,
            I => \c0.n23_adj_3364\
        );

    \I__11161\ : InMux
    port map (
            O => \N__51946\,
            I => \N__51943\
        );

    \I__11160\ : LocalMux
    port map (
            O => \N__51943\,
            I => \N__51939\
        );

    \I__11159\ : InMux
    port map (
            O => \N__51942\,
            I => \N__51936\
        );

    \I__11158\ : Span4Mux_v
    port map (
            O => \N__51939\,
            I => \N__51933\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__51936\,
            I => \N__51930\
        );

    \I__11156\ : Span4Mux_h
    port map (
            O => \N__51933\,
            I => \N__51927\
        );

    \I__11155\ : Span4Mux_v
    port map (
            O => \N__51930\,
            I => \N__51924\
        );

    \I__11154\ : Odrv4
    port map (
            O => \N__51927\,
            I => \c0.n24_adj_3335\
        );

    \I__11153\ : Odrv4
    port map (
            O => \N__51924\,
            I => \c0.n24_adj_3335\
        );

    \I__11152\ : CascadeMux
    port map (
            O => \N__51919\,
            I => \c0.n36_adj_3470_cascade_\
        );

    \I__11151\ : InMux
    port map (
            O => \N__51916\,
            I => \N__51913\
        );

    \I__11150\ : LocalMux
    port map (
            O => \N__51913\,
            I => \N__51909\
        );

    \I__11149\ : InMux
    port map (
            O => \N__51912\,
            I => \N__51906\
        );

    \I__11148\ : Span4Mux_v
    port map (
            O => \N__51909\,
            I => \N__51903\
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__51906\,
            I => \N__51900\
        );

    \I__11146\ : Odrv4
    port map (
            O => \N__51903\,
            I => \c0.n22_adj_3341\
        );

    \I__11145\ : Odrv4
    port map (
            O => \N__51900\,
            I => \c0.n22_adj_3341\
        );

    \I__11144\ : CascadeMux
    port map (
            O => \N__51895\,
            I => \c0.n11_adj_3124_cascade_\
        );

    \I__11143\ : InMux
    port map (
            O => \N__51892\,
            I => \N__51889\
        );

    \I__11142\ : LocalMux
    port map (
            O => \N__51889\,
            I => \N__51886\
        );

    \I__11141\ : Span4Mux_h
    port map (
            O => \N__51886\,
            I => \N__51882\
        );

    \I__11140\ : InMux
    port map (
            O => \N__51885\,
            I => \N__51879\
        );

    \I__11139\ : Odrv4
    port map (
            O => \N__51882\,
            I => \c0.n22_adj_3287\
        );

    \I__11138\ : LocalMux
    port map (
            O => \N__51879\,
            I => \c0.n22_adj_3287\
        );

    \I__11137\ : CascadeMux
    port map (
            O => \N__51874\,
            I => \c0.n47_adj_3286_cascade_\
        );

    \I__11136\ : InMux
    port map (
            O => \N__51871\,
            I => \N__51868\
        );

    \I__11135\ : LocalMux
    port map (
            O => \N__51868\,
            I => \c0.n51_adj_3290\
        );

    \I__11134\ : CascadeMux
    port map (
            O => \N__51865\,
            I => \c0.n52_adj_3288_cascade_\
        );

    \I__11133\ : InMux
    port map (
            O => \N__51862\,
            I => \N__51859\
        );

    \I__11132\ : LocalMux
    port map (
            O => \N__51859\,
            I => \N__51856\
        );

    \I__11131\ : Span4Mux_h
    port map (
            O => \N__51856\,
            I => \N__51853\
        );

    \I__11130\ : Span4Mux_v
    port map (
            O => \N__51853\,
            I => \N__51850\
        );

    \I__11129\ : Odrv4
    port map (
            O => \N__51850\,
            I => \c0.n6_adj_3291\
        );

    \I__11128\ : CascadeMux
    port map (
            O => \N__51847\,
            I => \N__51843\
        );

    \I__11127\ : CascadeMux
    port map (
            O => \N__51846\,
            I => \N__51840\
        );

    \I__11126\ : InMux
    port map (
            O => \N__51843\,
            I => \N__51837\
        );

    \I__11125\ : InMux
    port map (
            O => \N__51840\,
            I => \N__51834\
        );

    \I__11124\ : LocalMux
    port map (
            O => \N__51837\,
            I => \N__51830\
        );

    \I__11123\ : LocalMux
    port map (
            O => \N__51834\,
            I => \N__51827\
        );

    \I__11122\ : InMux
    port map (
            O => \N__51833\,
            I => \N__51824\
        );

    \I__11121\ : Span4Mux_h
    port map (
            O => \N__51830\,
            I => \N__51821\
        );

    \I__11120\ : Span4Mux_h
    port map (
            O => \N__51827\,
            I => \N__51818\
        );

    \I__11119\ : LocalMux
    port map (
            O => \N__51824\,
            I => \c0.data_in_frame_11_6\
        );

    \I__11118\ : Odrv4
    port map (
            O => \N__51821\,
            I => \c0.data_in_frame_11_6\
        );

    \I__11117\ : Odrv4
    port map (
            O => \N__51818\,
            I => \c0.data_in_frame_11_6\
        );

    \I__11116\ : CascadeMux
    port map (
            O => \N__51811\,
            I => \c0.n19909_cascade_\
        );

    \I__11115\ : InMux
    port map (
            O => \N__51808\,
            I => \N__51804\
        );

    \I__11114\ : InMux
    port map (
            O => \N__51807\,
            I => \N__51801\
        );

    \I__11113\ : LocalMux
    port map (
            O => \N__51804\,
            I => \N__51798\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__51801\,
            I => \N__51795\
        );

    \I__11111\ : Span4Mux_h
    port map (
            O => \N__51798\,
            I => \N__51792\
        );

    \I__11110\ : Odrv4
    port map (
            O => \N__51795\,
            I => \c0.n87\
        );

    \I__11109\ : Odrv4
    port map (
            O => \N__51792\,
            I => \c0.n87\
        );

    \I__11108\ : InMux
    port map (
            O => \N__51787\,
            I => \N__51782\
        );

    \I__11107\ : InMux
    port map (
            O => \N__51786\,
            I => \N__51777\
        );

    \I__11106\ : InMux
    port map (
            O => \N__51785\,
            I => \N__51777\
        );

    \I__11105\ : LocalMux
    port map (
            O => \N__51782\,
            I => \N__51770\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__51777\,
            I => \N__51770\
        );

    \I__11103\ : InMux
    port map (
            O => \N__51776\,
            I => \N__51765\
        );

    \I__11102\ : InMux
    port map (
            O => \N__51775\,
            I => \N__51765\
        );

    \I__11101\ : Odrv12
    port map (
            O => \N__51770\,
            I => \c0.n6_adj_3137\
        );

    \I__11100\ : LocalMux
    port map (
            O => \N__51765\,
            I => \c0.n6_adj_3137\
        );

    \I__11099\ : InMux
    port map (
            O => \N__51760\,
            I => \N__51756\
        );

    \I__11098\ : CascadeMux
    port map (
            O => \N__51759\,
            I => \N__51753\
        );

    \I__11097\ : LocalMux
    port map (
            O => \N__51756\,
            I => \N__51750\
        );

    \I__11096\ : InMux
    port map (
            O => \N__51753\,
            I => \N__51747\
        );

    \I__11095\ : Span4Mux_v
    port map (
            O => \N__51750\,
            I => \N__51744\
        );

    \I__11094\ : LocalMux
    port map (
            O => \N__51747\,
            I => \N__51741\
        );

    \I__11093\ : Span4Mux_h
    port map (
            O => \N__51744\,
            I => \N__51736\
        );

    \I__11092\ : Span4Mux_h
    port map (
            O => \N__51741\,
            I => \N__51736\
        );

    \I__11091\ : Span4Mux_v
    port map (
            O => \N__51736\,
            I => \N__51733\
        );

    \I__11090\ : Odrv4
    port map (
            O => \N__51733\,
            I => \c0.n35_adj_3098\
        );

    \I__11089\ : InMux
    port map (
            O => \N__51730\,
            I => \N__51726\
        );

    \I__11088\ : InMux
    port map (
            O => \N__51729\,
            I => \N__51723\
        );

    \I__11087\ : LocalMux
    port map (
            O => \N__51726\,
            I => \c0.n19909\
        );

    \I__11086\ : LocalMux
    port map (
            O => \N__51723\,
            I => \c0.n19909\
        );

    \I__11085\ : CascadeMux
    port map (
            O => \N__51718\,
            I => \N__51715\
        );

    \I__11084\ : InMux
    port map (
            O => \N__51715\,
            I => \N__51712\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__51712\,
            I => \N__51708\
        );

    \I__11082\ : InMux
    port map (
            O => \N__51711\,
            I => \N__51703\
        );

    \I__11081\ : Span4Mux_h
    port map (
            O => \N__51708\,
            I => \N__51700\
        );

    \I__11080\ : InMux
    port map (
            O => \N__51707\,
            I => \N__51695\
        );

    \I__11079\ : InMux
    port map (
            O => \N__51706\,
            I => \N__51695\
        );

    \I__11078\ : LocalMux
    port map (
            O => \N__51703\,
            I => \c0.data_in_frame_13_5\
        );

    \I__11077\ : Odrv4
    port map (
            O => \N__51700\,
            I => \c0.data_in_frame_13_5\
        );

    \I__11076\ : LocalMux
    port map (
            O => \N__51695\,
            I => \c0.data_in_frame_13_5\
        );

    \I__11075\ : InMux
    port map (
            O => \N__51688\,
            I => \N__51682\
        );

    \I__11074\ : InMux
    port map (
            O => \N__51687\,
            I => \N__51675\
        );

    \I__11073\ : InMux
    port map (
            O => \N__51686\,
            I => \N__51675\
        );

    \I__11072\ : InMux
    port map (
            O => \N__51685\,
            I => \N__51675\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__51682\,
            I => \N__51669\
        );

    \I__11070\ : LocalMux
    port map (
            O => \N__51675\,
            I => \N__51666\
        );

    \I__11069\ : InMux
    port map (
            O => \N__51674\,
            I => \N__51663\
        );

    \I__11068\ : InMux
    port map (
            O => \N__51673\,
            I => \N__51658\
        );

    \I__11067\ : InMux
    port map (
            O => \N__51672\,
            I => \N__51658\
        );

    \I__11066\ : Odrv4
    port map (
            O => \N__51669\,
            I => \c0.n20826\
        );

    \I__11065\ : Odrv4
    port map (
            O => \N__51666\,
            I => \c0.n20826\
        );

    \I__11064\ : LocalMux
    port map (
            O => \N__51663\,
            I => \c0.n20826\
        );

    \I__11063\ : LocalMux
    port map (
            O => \N__51658\,
            I => \c0.n20826\
        );

    \I__11062\ : InMux
    port map (
            O => \N__51649\,
            I => \N__51646\
        );

    \I__11061\ : LocalMux
    port map (
            O => \N__51646\,
            I => \N__51643\
        );

    \I__11060\ : Odrv12
    port map (
            O => \N__51643\,
            I => \c0.n54_adj_3234\
        );

    \I__11059\ : CascadeMux
    port map (
            O => \N__51640\,
            I => \c0.n43_adj_3232_cascade_\
        );

    \I__11058\ : InMux
    port map (
            O => \N__51637\,
            I => \N__51633\
        );

    \I__11057\ : InMux
    port map (
            O => \N__51636\,
            I => \N__51630\
        );

    \I__11056\ : LocalMux
    port map (
            O => \N__51633\,
            I => \N__51627\
        );

    \I__11055\ : LocalMux
    port map (
            O => \N__51630\,
            I => \N__51624\
        );

    \I__11054\ : Span4Mux_v
    port map (
            O => \N__51627\,
            I => \N__51618\
        );

    \I__11053\ : Span4Mux_h
    port map (
            O => \N__51624\,
            I => \N__51618\
        );

    \I__11052\ : InMux
    port map (
            O => \N__51623\,
            I => \N__51614\
        );

    \I__11051\ : Span4Mux_h
    port map (
            O => \N__51618\,
            I => \N__51611\
        );

    \I__11050\ : InMux
    port map (
            O => \N__51617\,
            I => \N__51608\
        );

    \I__11049\ : LocalMux
    port map (
            O => \N__51614\,
            I => \c0.n17849\
        );

    \I__11048\ : Odrv4
    port map (
            O => \N__51611\,
            I => \c0.n17849\
        );

    \I__11047\ : LocalMux
    port map (
            O => \N__51608\,
            I => \c0.n17849\
        );

    \I__11046\ : InMux
    port map (
            O => \N__51601\,
            I => \N__51598\
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__51598\,
            I => \c0.n49_adj_3237\
        );

    \I__11044\ : CascadeMux
    port map (
            O => \N__51595\,
            I => \c0.n7_adj_3225_cascade_\
        );

    \I__11043\ : CascadeMux
    port map (
            O => \N__51592\,
            I => \N__51589\
        );

    \I__11042\ : InMux
    port map (
            O => \N__51589\,
            I => \N__51583\
        );

    \I__11041\ : InMux
    port map (
            O => \N__51588\,
            I => \N__51583\
        );

    \I__11040\ : LocalMux
    port map (
            O => \N__51583\,
            I => \N__51579\
        );

    \I__11039\ : CascadeMux
    port map (
            O => \N__51582\,
            I => \N__51576\
        );

    \I__11038\ : Span4Mux_h
    port map (
            O => \N__51579\,
            I => \N__51573\
        );

    \I__11037\ : InMux
    port map (
            O => \N__51576\,
            I => \N__51570\
        );

    \I__11036\ : Span4Mux_h
    port map (
            O => \N__51573\,
            I => \N__51567\
        );

    \I__11035\ : LocalMux
    port map (
            O => \N__51570\,
            I => \N__51562\
        );

    \I__11034\ : Span4Mux_v
    port map (
            O => \N__51567\,
            I => \N__51562\
        );

    \I__11033\ : Odrv4
    port map (
            O => \N__51562\,
            I => \c0.data_in_frame_15_4\
        );

    \I__11032\ : InMux
    port map (
            O => \N__51559\,
            I => \N__51556\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__51556\,
            I => \c0.n7_adj_3225\
        );

    \I__11030\ : InMux
    port map (
            O => \N__51553\,
            I => \N__51550\
        );

    \I__11029\ : LocalMux
    port map (
            O => \N__51550\,
            I => \N__51547\
        );

    \I__11028\ : Odrv4
    port map (
            O => \N__51547\,
            I => \c0.n44_adj_3226\
        );

    \I__11027\ : InMux
    port map (
            O => \N__51544\,
            I => \N__51541\
        );

    \I__11026\ : LocalMux
    port map (
            O => \N__51541\,
            I => \N__51535\
        );

    \I__11025\ : InMux
    port map (
            O => \N__51540\,
            I => \N__51532\
        );

    \I__11024\ : InMux
    port map (
            O => \N__51539\,
            I => \N__51527\
        );

    \I__11023\ : InMux
    port map (
            O => \N__51538\,
            I => \N__51527\
        );

    \I__11022\ : Odrv12
    port map (
            O => \N__51535\,
            I => \c0.data_in_frame_10_4\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__51532\,
            I => \c0.data_in_frame_10_4\
        );

    \I__11020\ : LocalMux
    port map (
            O => \N__51527\,
            I => \c0.data_in_frame_10_4\
        );

    \I__11019\ : CascadeMux
    port map (
            O => \N__51520\,
            I => \N__51515\
        );

    \I__11018\ : CascadeMux
    port map (
            O => \N__51519\,
            I => \N__51510\
        );

    \I__11017\ : CascadeMux
    port map (
            O => \N__51518\,
            I => \N__51507\
        );

    \I__11016\ : InMux
    port map (
            O => \N__51515\,
            I => \N__51504\
        );

    \I__11015\ : InMux
    port map (
            O => \N__51514\,
            I => \N__51501\
        );

    \I__11014\ : InMux
    port map (
            O => \N__51513\,
            I => \N__51498\
        );

    \I__11013\ : InMux
    port map (
            O => \N__51510\,
            I => \N__51495\
        );

    \I__11012\ : InMux
    port map (
            O => \N__51507\,
            I => \N__51492\
        );

    \I__11011\ : LocalMux
    port map (
            O => \N__51504\,
            I => \N__51489\
        );

    \I__11010\ : LocalMux
    port map (
            O => \N__51501\,
            I => \N__51484\
        );

    \I__11009\ : LocalMux
    port map (
            O => \N__51498\,
            I => \N__51484\
        );

    \I__11008\ : LocalMux
    port map (
            O => \N__51495\,
            I => \N__51479\
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__51492\,
            I => \N__51479\
        );

    \I__11006\ : Span4Mux_v
    port map (
            O => \N__51489\,
            I => \N__51475\
        );

    \I__11005\ : Span4Mux_v
    port map (
            O => \N__51484\,
            I => \N__51472\
        );

    \I__11004\ : Span4Mux_v
    port map (
            O => \N__51479\,
            I => \N__51469\
        );

    \I__11003\ : InMux
    port map (
            O => \N__51478\,
            I => \N__51466\
        );

    \I__11002\ : Odrv4
    port map (
            O => \N__51475\,
            I => \c0.data_in_frame_8_1\
        );

    \I__11001\ : Odrv4
    port map (
            O => \N__51472\,
            I => \c0.data_in_frame_8_1\
        );

    \I__11000\ : Odrv4
    port map (
            O => \N__51469\,
            I => \c0.data_in_frame_8_1\
        );

    \I__10999\ : LocalMux
    port map (
            O => \N__51466\,
            I => \c0.data_in_frame_8_1\
        );

    \I__10998\ : CascadeMux
    port map (
            O => \N__51457\,
            I => \N__51453\
        );

    \I__10997\ : CascadeMux
    port map (
            O => \N__51456\,
            I => \N__51450\
        );

    \I__10996\ : InMux
    port map (
            O => \N__51453\,
            I => \N__51445\
        );

    \I__10995\ : InMux
    port map (
            O => \N__51450\,
            I => \N__51445\
        );

    \I__10994\ : LocalMux
    port map (
            O => \N__51445\,
            I => \N__51442\
        );

    \I__10993\ : Span4Mux_h
    port map (
            O => \N__51442\,
            I => \N__51439\
        );

    \I__10992\ : Odrv4
    port map (
            O => \N__51439\,
            I => \c0.n41_adj_3365\
        );

    \I__10991\ : InMux
    port map (
            O => \N__51436\,
            I => \N__51433\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__51433\,
            I => \N__51429\
        );

    \I__10989\ : InMux
    port map (
            O => \N__51432\,
            I => \N__51426\
        );

    \I__10988\ : Odrv4
    port map (
            O => \N__51429\,
            I => \c0.n16_adj_3218\
        );

    \I__10987\ : LocalMux
    port map (
            O => \N__51426\,
            I => \c0.n16_adj_3218\
        );

    \I__10986\ : InMux
    port map (
            O => \N__51421\,
            I => \N__51418\
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__51418\,
            I => \c0.n48\
        );

    \I__10984\ : InMux
    port map (
            O => \N__51415\,
            I => \N__51411\
        );

    \I__10983\ : CascadeMux
    port map (
            O => \N__51414\,
            I => \N__51407\
        );

    \I__10982\ : LocalMux
    port map (
            O => \N__51411\,
            I => \N__51403\
        );

    \I__10981\ : InMux
    port map (
            O => \N__51410\,
            I => \N__51400\
        );

    \I__10980\ : InMux
    port map (
            O => \N__51407\,
            I => \N__51396\
        );

    \I__10979\ : CascadeMux
    port map (
            O => \N__51406\,
            I => \N__51393\
        );

    \I__10978\ : Span4Mux_v
    port map (
            O => \N__51403\,
            I => \N__51390\
        );

    \I__10977\ : LocalMux
    port map (
            O => \N__51400\,
            I => \N__51387\
        );

    \I__10976\ : InMux
    port map (
            O => \N__51399\,
            I => \N__51383\
        );

    \I__10975\ : LocalMux
    port map (
            O => \N__51396\,
            I => \N__51380\
        );

    \I__10974\ : InMux
    port map (
            O => \N__51393\,
            I => \N__51377\
        );

    \I__10973\ : Span4Mux_h
    port map (
            O => \N__51390\,
            I => \N__51374\
        );

    \I__10972\ : Span12Mux_s10_v
    port map (
            O => \N__51387\,
            I => \N__51371\
        );

    \I__10971\ : InMux
    port map (
            O => \N__51386\,
            I => \N__51368\
        );

    \I__10970\ : LocalMux
    port map (
            O => \N__51383\,
            I => \N__51365\
        );

    \I__10969\ : Span4Mux_h
    port map (
            O => \N__51380\,
            I => \N__51362\
        );

    \I__10968\ : LocalMux
    port map (
            O => \N__51377\,
            I => \c0.data_in_frame_5_1\
        );

    \I__10967\ : Odrv4
    port map (
            O => \N__51374\,
            I => \c0.data_in_frame_5_1\
        );

    \I__10966\ : Odrv12
    port map (
            O => \N__51371\,
            I => \c0.data_in_frame_5_1\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__51368\,
            I => \c0.data_in_frame_5_1\
        );

    \I__10964\ : Odrv4
    port map (
            O => \N__51365\,
            I => \c0.data_in_frame_5_1\
        );

    \I__10963\ : Odrv4
    port map (
            O => \N__51362\,
            I => \c0.data_in_frame_5_1\
        );

    \I__10962\ : InMux
    port map (
            O => \N__51349\,
            I => \N__51346\
        );

    \I__10961\ : LocalMux
    port map (
            O => \N__51346\,
            I => \N__51342\
        );

    \I__10960\ : InMux
    port map (
            O => \N__51345\,
            I => \N__51339\
        );

    \I__10959\ : Span4Mux_v
    port map (
            O => \N__51342\,
            I => \N__51335\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__51339\,
            I => \N__51332\
        );

    \I__10957\ : InMux
    port map (
            O => \N__51338\,
            I => \N__51327\
        );

    \I__10956\ : Span4Mux_v
    port map (
            O => \N__51335\,
            I => \N__51324\
        );

    \I__10955\ : Span4Mux_v
    port map (
            O => \N__51332\,
            I => \N__51321\
        );

    \I__10954\ : InMux
    port map (
            O => \N__51331\,
            I => \N__51318\
        );

    \I__10953\ : InMux
    port map (
            O => \N__51330\,
            I => \N__51315\
        );

    \I__10952\ : LocalMux
    port map (
            O => \N__51327\,
            I => \N__51312\
        );

    \I__10951\ : Odrv4
    port map (
            O => \N__51324\,
            I => \c0.n20224\
        );

    \I__10950\ : Odrv4
    port map (
            O => \N__51321\,
            I => \c0.n20224\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__51318\,
            I => \c0.n20224\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__51315\,
            I => \c0.n20224\
        );

    \I__10947\ : Odrv12
    port map (
            O => \N__51312\,
            I => \c0.n20224\
        );

    \I__10946\ : CascadeMux
    port map (
            O => \N__51301\,
            I => \N__51298\
        );

    \I__10945\ : InMux
    port map (
            O => \N__51298\,
            I => \N__51295\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__51295\,
            I => \c0.n5_adj_3549\
        );

    \I__10943\ : InMux
    port map (
            O => \N__51292\,
            I => \N__51288\
        );

    \I__10942\ : InMux
    port map (
            O => \N__51291\,
            I => \N__51284\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__51288\,
            I => \N__51279\
        );

    \I__10940\ : InMux
    port map (
            O => \N__51287\,
            I => \N__51276\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__51284\,
            I => \N__51273\
        );

    \I__10938\ : InMux
    port map (
            O => \N__51283\,
            I => \N__51270\
        );

    \I__10937\ : CascadeMux
    port map (
            O => \N__51282\,
            I => \N__51267\
        );

    \I__10936\ : Span4Mux_v
    port map (
            O => \N__51279\,
            I => \N__51261\
        );

    \I__10935\ : LocalMux
    port map (
            O => \N__51276\,
            I => \N__51261\
        );

    \I__10934\ : Span4Mux_h
    port map (
            O => \N__51273\,
            I => \N__51252\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__51270\,
            I => \N__51249\
        );

    \I__10932\ : InMux
    port map (
            O => \N__51267\,
            I => \N__51244\
        );

    \I__10931\ : InMux
    port map (
            O => \N__51266\,
            I => \N__51244\
        );

    \I__10930\ : Span4Mux_h
    port map (
            O => \N__51261\,
            I => \N__51241\
        );

    \I__10929\ : InMux
    port map (
            O => \N__51260\,
            I => \N__51234\
        );

    \I__10928\ : InMux
    port map (
            O => \N__51259\,
            I => \N__51234\
        );

    \I__10927\ : InMux
    port map (
            O => \N__51258\,
            I => \N__51234\
        );

    \I__10926\ : InMux
    port map (
            O => \N__51257\,
            I => \N__51227\
        );

    \I__10925\ : InMux
    port map (
            O => \N__51256\,
            I => \N__51227\
        );

    \I__10924\ : InMux
    port map (
            O => \N__51255\,
            I => \N__51227\
        );

    \I__10923\ : Odrv4
    port map (
            O => \N__51252\,
            I => \c0.data_in_frame_4_7\
        );

    \I__10922\ : Odrv4
    port map (
            O => \N__51249\,
            I => \c0.data_in_frame_4_7\
        );

    \I__10921\ : LocalMux
    port map (
            O => \N__51244\,
            I => \c0.data_in_frame_4_7\
        );

    \I__10920\ : Odrv4
    port map (
            O => \N__51241\,
            I => \c0.data_in_frame_4_7\
        );

    \I__10919\ : LocalMux
    port map (
            O => \N__51234\,
            I => \c0.data_in_frame_4_7\
        );

    \I__10918\ : LocalMux
    port map (
            O => \N__51227\,
            I => \c0.data_in_frame_4_7\
        );

    \I__10917\ : InMux
    port map (
            O => \N__51214\,
            I => \N__51211\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__51211\,
            I => \c0.n11613\
        );

    \I__10915\ : InMux
    port map (
            O => \N__51208\,
            I => \N__51204\
        );

    \I__10914\ : InMux
    port map (
            O => \N__51207\,
            I => \N__51201\
        );

    \I__10913\ : LocalMux
    port map (
            O => \N__51204\,
            I => \N__51197\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__51201\,
            I => \N__51194\
        );

    \I__10911\ : InMux
    port map (
            O => \N__51200\,
            I => \N__51191\
        );

    \I__10910\ : Span4Mux_h
    port map (
            O => \N__51197\,
            I => \N__51188\
        );

    \I__10909\ : Span4Mux_h
    port map (
            O => \N__51194\,
            I => \N__51185\
        );

    \I__10908\ : LocalMux
    port map (
            O => \N__51191\,
            I => \c0.data_in_frame_17_6\
        );

    \I__10907\ : Odrv4
    port map (
            O => \N__51188\,
            I => \c0.data_in_frame_17_6\
        );

    \I__10906\ : Odrv4
    port map (
            O => \N__51185\,
            I => \c0.data_in_frame_17_6\
        );

    \I__10905\ : InMux
    port map (
            O => \N__51178\,
            I => \N__51175\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__51175\,
            I => \N__51172\
        );

    \I__10903\ : Span4Mux_v
    port map (
            O => \N__51172\,
            I => \N__51168\
        );

    \I__10902\ : InMux
    port map (
            O => \N__51171\,
            I => \N__51165\
        );

    \I__10901\ : Span4Mux_h
    port map (
            O => \N__51168\,
            I => \N__51162\
        );

    \I__10900\ : LocalMux
    port map (
            O => \N__51165\,
            I => data_in_frame_18_0
        );

    \I__10899\ : Odrv4
    port map (
            O => \N__51162\,
            I => data_in_frame_18_0
        );

    \I__10898\ : CascadeMux
    port map (
            O => \N__51157\,
            I => \c0.n11613_cascade_\
        );

    \I__10897\ : InMux
    port map (
            O => \N__51154\,
            I => \N__51150\
        );

    \I__10896\ : InMux
    port map (
            O => \N__51153\,
            I => \N__51147\
        );

    \I__10895\ : LocalMux
    port map (
            O => \N__51150\,
            I => \N__51142\
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__51147\,
            I => \N__51142\
        );

    \I__10893\ : Odrv4
    port map (
            O => \N__51142\,
            I => \c0.n19477\
        );

    \I__10892\ : InMux
    port map (
            O => \N__51139\,
            I => \N__51136\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__51136\,
            I => \c0.n17_adj_3482\
        );

    \I__10890\ : InMux
    port map (
            O => \N__51133\,
            I => \N__51130\
        );

    \I__10889\ : LocalMux
    port map (
            O => \N__51130\,
            I => \N__51126\
        );

    \I__10888\ : CascadeMux
    port map (
            O => \N__51129\,
            I => \N__51123\
        );

    \I__10887\ : Span4Mux_h
    port map (
            O => \N__51126\,
            I => \N__51119\
        );

    \I__10886\ : InMux
    port map (
            O => \N__51123\,
            I => \N__51114\
        );

    \I__10885\ : InMux
    port map (
            O => \N__51122\,
            I => \N__51114\
        );

    \I__10884\ : Odrv4
    port map (
            O => \N__51119\,
            I => \c0.data_in_frame_13_6\
        );

    \I__10883\ : LocalMux
    port map (
            O => \N__51114\,
            I => \c0.data_in_frame_13_6\
        );

    \I__10882\ : InMux
    port map (
            O => \N__51109\,
            I => \N__51105\
        );

    \I__10881\ : InMux
    port map (
            O => \N__51108\,
            I => \N__51101\
        );

    \I__10880\ : LocalMux
    port map (
            O => \N__51105\,
            I => \N__51098\
        );

    \I__10879\ : CascadeMux
    port map (
            O => \N__51104\,
            I => \N__51094\
        );

    \I__10878\ : LocalMux
    port map (
            O => \N__51101\,
            I => \N__51091\
        );

    \I__10877\ : Span4Mux_v
    port map (
            O => \N__51098\,
            I => \N__51087\
        );

    \I__10876\ : InMux
    port map (
            O => \N__51097\,
            I => \N__51084\
        );

    \I__10875\ : InMux
    port map (
            O => \N__51094\,
            I => \N__51081\
        );

    \I__10874\ : Span4Mux_h
    port map (
            O => \N__51091\,
            I => \N__51078\
        );

    \I__10873\ : InMux
    port map (
            O => \N__51090\,
            I => \N__51075\
        );

    \I__10872\ : Span4Mux_h
    port map (
            O => \N__51087\,
            I => \N__51070\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__51084\,
            I => \N__51070\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__51081\,
            I => \c0.data_in_frame_7_4\
        );

    \I__10869\ : Odrv4
    port map (
            O => \N__51078\,
            I => \c0.data_in_frame_7_4\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__51075\,
            I => \c0.data_in_frame_7_4\
        );

    \I__10867\ : Odrv4
    port map (
            O => \N__51070\,
            I => \c0.data_in_frame_7_4\
        );

    \I__10866\ : InMux
    port map (
            O => \N__51061\,
            I => \N__51058\
        );

    \I__10865\ : LocalMux
    port map (
            O => \N__51058\,
            I => \N__51055\
        );

    \I__10864\ : Span4Mux_v
    port map (
            O => \N__51055\,
            I => \N__51051\
        );

    \I__10863\ : InMux
    port map (
            O => \N__51054\,
            I => \N__51048\
        );

    \I__10862\ : Odrv4
    port map (
            O => \N__51051\,
            I => \c0.n20391\
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__51048\,
            I => \c0.n20391\
        );

    \I__10860\ : InMux
    port map (
            O => \N__51043\,
            I => \N__51040\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__51040\,
            I => \c0.n4\
        );

    \I__10858\ : InMux
    port map (
            O => \N__51037\,
            I => \N__51034\
        );

    \I__10857\ : LocalMux
    port map (
            O => \N__51034\,
            I => \N__51030\
        );

    \I__10856\ : InMux
    port map (
            O => \N__51033\,
            I => \N__51027\
        );

    \I__10855\ : Span4Mux_v
    port map (
            O => \N__51030\,
            I => \N__51022\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__51027\,
            I => \N__51022\
        );

    \I__10853\ : Span4Mux_h
    port map (
            O => \N__51022\,
            I => \N__51019\
        );

    \I__10852\ : Odrv4
    port map (
            O => \N__51019\,
            I => \c0.n12026\
        );

    \I__10851\ : InMux
    port map (
            O => \N__51016\,
            I => \N__51012\
        );

    \I__10850\ : InMux
    port map (
            O => \N__51015\,
            I => \N__51009\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__51012\,
            I => \N__51006\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__51009\,
            I => \N__51003\
        );

    \I__10847\ : Span4Mux_v
    port map (
            O => \N__51006\,
            I => \N__51000\
        );

    \I__10846\ : Span4Mux_v
    port map (
            O => \N__51003\,
            I => \N__50997\
        );

    \I__10845\ : Odrv4
    port map (
            O => \N__51000\,
            I => \c0.n5\
        );

    \I__10844\ : Odrv4
    port map (
            O => \N__50997\,
            I => \c0.n5\
        );

    \I__10843\ : CascadeMux
    port map (
            O => \N__50992\,
            I => \c0.n4_cascade_\
        );

    \I__10842\ : InMux
    port map (
            O => \N__50989\,
            I => \N__50985\
        );

    \I__10841\ : InMux
    port map (
            O => \N__50988\,
            I => \N__50981\
        );

    \I__10840\ : LocalMux
    port map (
            O => \N__50985\,
            I => \N__50978\
        );

    \I__10839\ : CascadeMux
    port map (
            O => \N__50984\,
            I => \N__50974\
        );

    \I__10838\ : LocalMux
    port map (
            O => \N__50981\,
            I => \N__50971\
        );

    \I__10837\ : Span4Mux_h
    port map (
            O => \N__50978\,
            I => \N__50968\
        );

    \I__10836\ : InMux
    port map (
            O => \N__50977\,
            I => \N__50965\
        );

    \I__10835\ : InMux
    port map (
            O => \N__50974\,
            I => \N__50962\
        );

    \I__10834\ : Span4Mux_h
    port map (
            O => \N__50971\,
            I => \N__50959\
        );

    \I__10833\ : Span4Mux_v
    port map (
            O => \N__50968\,
            I => \N__50956\
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__50965\,
            I => \N__50953\
        );

    \I__10831\ : LocalMux
    port map (
            O => \N__50962\,
            I => \c0.data_in_frame_11_4\
        );

    \I__10830\ : Odrv4
    port map (
            O => \N__50959\,
            I => \c0.data_in_frame_11_4\
        );

    \I__10829\ : Odrv4
    port map (
            O => \N__50956\,
            I => \c0.data_in_frame_11_4\
        );

    \I__10828\ : Odrv12
    port map (
            O => \N__50953\,
            I => \c0.data_in_frame_11_4\
        );

    \I__10827\ : CascadeMux
    port map (
            O => \N__50944\,
            I => \N__50941\
        );

    \I__10826\ : InMux
    port map (
            O => \N__50941\,
            I => \N__50938\
        );

    \I__10825\ : LocalMux
    port map (
            O => \N__50938\,
            I => \N__50934\
        );

    \I__10824\ : CascadeMux
    port map (
            O => \N__50937\,
            I => \N__50930\
        );

    \I__10823\ : Span4Mux_v
    port map (
            O => \N__50934\,
            I => \N__50927\
        );

    \I__10822\ : InMux
    port map (
            O => \N__50933\,
            I => \N__50924\
        );

    \I__10821\ : InMux
    port map (
            O => \N__50930\,
            I => \N__50921\
        );

    \I__10820\ : Span4Mux_h
    port map (
            O => \N__50927\,
            I => \N__50918\
        );

    \I__10819\ : LocalMux
    port map (
            O => \N__50924\,
            I => \N__50915\
        );

    \I__10818\ : LocalMux
    port map (
            O => \N__50921\,
            I => \c0.data_in_frame_10_0\
        );

    \I__10817\ : Odrv4
    port map (
            O => \N__50918\,
            I => \c0.data_in_frame_10_0\
        );

    \I__10816\ : Odrv4
    port map (
            O => \N__50915\,
            I => \c0.data_in_frame_10_0\
        );

    \I__10815\ : InMux
    port map (
            O => \N__50908\,
            I => \N__50905\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__50905\,
            I => \N__50900\
        );

    \I__10813\ : InMux
    port map (
            O => \N__50904\,
            I => \N__50897\
        );

    \I__10812\ : CascadeMux
    port map (
            O => \N__50903\,
            I => \N__50894\
        );

    \I__10811\ : Span4Mux_v
    port map (
            O => \N__50900\,
            I => \N__50891\
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__50897\,
            I => \N__50888\
        );

    \I__10809\ : InMux
    port map (
            O => \N__50894\,
            I => \N__50885\
        );

    \I__10808\ : Span4Mux_h
    port map (
            O => \N__50891\,
            I => \N__50882\
        );

    \I__10807\ : Span4Mux_h
    port map (
            O => \N__50888\,
            I => \N__50879\
        );

    \I__10806\ : LocalMux
    port map (
            O => \N__50885\,
            I => \c0.data_in_frame_21_0\
        );

    \I__10805\ : Odrv4
    port map (
            O => \N__50882\,
            I => \c0.data_in_frame_21_0\
        );

    \I__10804\ : Odrv4
    port map (
            O => \N__50879\,
            I => \c0.data_in_frame_21_0\
        );

    \I__10803\ : CascadeMux
    port map (
            O => \N__50872\,
            I => \c0.n36_adj_3212_cascade_\
        );

    \I__10802\ : InMux
    port map (
            O => \N__50869\,
            I => \N__50866\
        );

    \I__10801\ : LocalMux
    port map (
            O => \N__50866\,
            I => \c0.n41_adj_3213\
        );

    \I__10800\ : InMux
    port map (
            O => \N__50863\,
            I => \N__50860\
        );

    \I__10799\ : LocalMux
    port map (
            O => \N__50860\,
            I => \N__50857\
        );

    \I__10798\ : Span4Mux_v
    port map (
            O => \N__50857\,
            I => \N__50854\
        );

    \I__10797\ : Span4Mux_h
    port map (
            O => \N__50854\,
            I => \N__50849\
        );

    \I__10796\ : InMux
    port map (
            O => \N__50853\,
            I => \N__50844\
        );

    \I__10795\ : InMux
    port map (
            O => \N__50852\,
            I => \N__50844\
        );

    \I__10794\ : Odrv4
    port map (
            O => \N__50849\,
            I => \c0.n20340\
        );

    \I__10793\ : LocalMux
    port map (
            O => \N__50844\,
            I => \c0.n20340\
        );

    \I__10792\ : CascadeMux
    port map (
            O => \N__50839\,
            I => \c0.n11651_cascade_\
        );

    \I__10791\ : InMux
    port map (
            O => \N__50836\,
            I => \N__50833\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__50833\,
            I => \c0.n27_adj_3082\
        );

    \I__10789\ : InMux
    port map (
            O => \N__50830\,
            I => \N__50826\
        );

    \I__10788\ : InMux
    port map (
            O => \N__50829\,
            I => \N__50823\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__50826\,
            I => \N__50819\
        );

    \I__10786\ : LocalMux
    port map (
            O => \N__50823\,
            I => \N__50816\
        );

    \I__10785\ : InMux
    port map (
            O => \N__50822\,
            I => \N__50813\
        );

    \I__10784\ : Span4Mux_h
    port map (
            O => \N__50819\,
            I => \N__50810\
        );

    \I__10783\ : Span4Mux_h
    port map (
            O => \N__50816\,
            I => \N__50807\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__50813\,
            I => \N__50804\
        );

    \I__10781\ : Odrv4
    port map (
            O => \N__50810\,
            I => \c0.n11800\
        );

    \I__10780\ : Odrv4
    port map (
            O => \N__50807\,
            I => \c0.n11800\
        );

    \I__10779\ : Odrv4
    port map (
            O => \N__50804\,
            I => \c0.n11800\
        );

    \I__10778\ : InMux
    port map (
            O => \N__50797\,
            I => \N__50793\
        );

    \I__10777\ : InMux
    port map (
            O => \N__50796\,
            I => \N__50790\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__50793\,
            I => \c0.n31\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__50790\,
            I => \c0.n31\
        );

    \I__10774\ : CascadeMux
    port map (
            O => \N__50785\,
            I => \N__50781\
        );

    \I__10773\ : CascadeMux
    port map (
            O => \N__50784\,
            I => \N__50778\
        );

    \I__10772\ : InMux
    port map (
            O => \N__50781\,
            I => \N__50775\
        );

    \I__10771\ : InMux
    port map (
            O => \N__50778\,
            I => \N__50772\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__50775\,
            I => \N__50769\
        );

    \I__10769\ : LocalMux
    port map (
            O => \N__50772\,
            I => \N__50766\
        );

    \I__10768\ : Span4Mux_v
    port map (
            O => \N__50769\,
            I => \N__50763\
        );

    \I__10767\ : Span4Mux_v
    port map (
            O => \N__50766\,
            I => \N__50760\
        );

    \I__10766\ : Span4Mux_h
    port map (
            O => \N__50763\,
            I => \N__50757\
        );

    \I__10765\ : Span4Mux_h
    port map (
            O => \N__50760\,
            I => \N__50754\
        );

    \I__10764\ : Odrv4
    port map (
            O => \N__50757\,
            I => \c0.n37_adj_3153\
        );

    \I__10763\ : Odrv4
    port map (
            O => \N__50754\,
            I => \c0.n37_adj_3153\
        );

    \I__10762\ : InMux
    port map (
            O => \N__50749\,
            I => \N__50746\
        );

    \I__10761\ : LocalMux
    port map (
            O => \N__50746\,
            I => \N__50743\
        );

    \I__10760\ : Odrv12
    port map (
            O => \N__50743\,
            I => \c0.n35_adj_3233\
        );

    \I__10759\ : InMux
    port map (
            O => \N__50740\,
            I => \N__50736\
        );

    \I__10758\ : InMux
    port map (
            O => \N__50739\,
            I => \N__50733\
        );

    \I__10757\ : LocalMux
    port map (
            O => \N__50736\,
            I => \N__50730\
        );

    \I__10756\ : LocalMux
    port map (
            O => \N__50733\,
            I => \N__50727\
        );

    \I__10755\ : Span4Mux_h
    port map (
            O => \N__50730\,
            I => \N__50722\
        );

    \I__10754\ : Span4Mux_v
    port map (
            O => \N__50727\,
            I => \N__50722\
        );

    \I__10753\ : Span4Mux_v
    port map (
            O => \N__50722\,
            I => \N__50719\
        );

    \I__10752\ : Odrv4
    port map (
            O => \N__50719\,
            I => \c0.n60\
        );

    \I__10751\ : CascadeMux
    port map (
            O => \N__50716\,
            I => \c0.n52_adj_3223_cascade_\
        );

    \I__10750\ : CascadeMux
    port map (
            O => \N__50713\,
            I => \N__50710\
        );

    \I__10749\ : InMux
    port map (
            O => \N__50710\,
            I => \N__50707\
        );

    \I__10748\ : LocalMux
    port map (
            O => \N__50707\,
            I => \N__50704\
        );

    \I__10747\ : Span4Mux_h
    port map (
            O => \N__50704\,
            I => \N__50701\
        );

    \I__10746\ : Odrv4
    port map (
            O => \N__50701\,
            I => \c0.n60_adj_3503\
        );

    \I__10745\ : InMux
    port map (
            O => \N__50698\,
            I => \N__50695\
        );

    \I__10744\ : LocalMux
    port map (
            O => \N__50695\,
            I => \N__50692\
        );

    \I__10743\ : Span4Mux_h
    port map (
            O => \N__50692\,
            I => \N__50688\
        );

    \I__10742\ : InMux
    port map (
            O => \N__50691\,
            I => \N__50685\
        );

    \I__10741\ : Odrv4
    port map (
            O => \N__50688\,
            I => \c0.n52_adj_3402\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__50685\,
            I => \c0.n52_adj_3402\
        );

    \I__10739\ : CascadeMux
    port map (
            O => \N__50680\,
            I => \N__50675\
        );

    \I__10738\ : CascadeMux
    port map (
            O => \N__50679\,
            I => \N__50669\
        );

    \I__10737\ : InMux
    port map (
            O => \N__50678\,
            I => \N__50666\
        );

    \I__10736\ : InMux
    port map (
            O => \N__50675\,
            I => \N__50663\
        );

    \I__10735\ : InMux
    port map (
            O => \N__50674\,
            I => \N__50660\
        );

    \I__10734\ : InMux
    port map (
            O => \N__50673\,
            I => \N__50654\
        );

    \I__10733\ : InMux
    port map (
            O => \N__50672\,
            I => \N__50654\
        );

    \I__10732\ : InMux
    port map (
            O => \N__50669\,
            I => \N__50651\
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__50666\,
            I => \N__50648\
        );

    \I__10730\ : LocalMux
    port map (
            O => \N__50663\,
            I => \N__50645\
        );

    \I__10729\ : LocalMux
    port map (
            O => \N__50660\,
            I => \N__50642\
        );

    \I__10728\ : InMux
    port map (
            O => \N__50659\,
            I => \N__50636\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__50654\,
            I => \N__50633\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__50651\,
            I => \N__50624\
        );

    \I__10725\ : Span4Mux_v
    port map (
            O => \N__50648\,
            I => \N__50624\
        );

    \I__10724\ : Span4Mux_v
    port map (
            O => \N__50645\,
            I => \N__50624\
        );

    \I__10723\ : Span4Mux_h
    port map (
            O => \N__50642\,
            I => \N__50624\
        );

    \I__10722\ : InMux
    port map (
            O => \N__50641\,
            I => \N__50621\
        );

    \I__10721\ : InMux
    port map (
            O => \N__50640\,
            I => \N__50616\
        );

    \I__10720\ : InMux
    port map (
            O => \N__50639\,
            I => \N__50616\
        );

    \I__10719\ : LocalMux
    port map (
            O => \N__50636\,
            I => \c0.data_in_frame_3_1\
        );

    \I__10718\ : Odrv12
    port map (
            O => \N__50633\,
            I => \c0.data_in_frame_3_1\
        );

    \I__10717\ : Odrv4
    port map (
            O => \N__50624\,
            I => \c0.data_in_frame_3_1\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__50621\,
            I => \c0.data_in_frame_3_1\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__50616\,
            I => \c0.data_in_frame_3_1\
        );

    \I__10714\ : InMux
    port map (
            O => \N__50605\,
            I => \N__50596\
        );

    \I__10713\ : InMux
    port map (
            O => \N__50604\,
            I => \N__50593\
        );

    \I__10712\ : InMux
    port map (
            O => \N__50603\,
            I => \N__50589\
        );

    \I__10711\ : InMux
    port map (
            O => \N__50602\,
            I => \N__50586\
        );

    \I__10710\ : InMux
    port map (
            O => \N__50601\,
            I => \N__50583\
        );

    \I__10709\ : CascadeMux
    port map (
            O => \N__50600\,
            I => \N__50579\
        );

    \I__10708\ : CascadeMux
    port map (
            O => \N__50599\,
            I => \N__50576\
        );

    \I__10707\ : LocalMux
    port map (
            O => \N__50596\,
            I => \N__50573\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__50593\,
            I => \N__50570\
        );

    \I__10705\ : InMux
    port map (
            O => \N__50592\,
            I => \N__50567\
        );

    \I__10704\ : LocalMux
    port map (
            O => \N__50589\,
            I => \N__50563\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__50586\,
            I => \N__50558\
        );

    \I__10702\ : LocalMux
    port map (
            O => \N__50583\,
            I => \N__50558\
        );

    \I__10701\ : CascadeMux
    port map (
            O => \N__50582\,
            I => \N__50555\
        );

    \I__10700\ : InMux
    port map (
            O => \N__50579\,
            I => \N__50545\
        );

    \I__10699\ : InMux
    port map (
            O => \N__50576\,
            I => \N__50545\
        );

    \I__10698\ : Span4Mux_h
    port map (
            O => \N__50573\,
            I => \N__50538\
        );

    \I__10697\ : Span4Mux_h
    port map (
            O => \N__50570\,
            I => \N__50538\
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__50567\,
            I => \N__50538\
        );

    \I__10695\ : InMux
    port map (
            O => \N__50566\,
            I => \N__50535\
        );

    \I__10694\ : Span4Mux_h
    port map (
            O => \N__50563\,
            I => \N__50530\
        );

    \I__10693\ : Span4Mux_v
    port map (
            O => \N__50558\,
            I => \N__50530\
        );

    \I__10692\ : InMux
    port map (
            O => \N__50555\,
            I => \N__50525\
        );

    \I__10691\ : InMux
    port map (
            O => \N__50554\,
            I => \N__50525\
        );

    \I__10690\ : InMux
    port map (
            O => \N__50553\,
            I => \N__50518\
        );

    \I__10689\ : InMux
    port map (
            O => \N__50552\,
            I => \N__50518\
        );

    \I__10688\ : InMux
    port map (
            O => \N__50551\,
            I => \N__50518\
        );

    \I__10687\ : InMux
    port map (
            O => \N__50550\,
            I => \N__50515\
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__50545\,
            I => data_in_frame_0_5
        );

    \I__10685\ : Odrv4
    port map (
            O => \N__50538\,
            I => data_in_frame_0_5
        );

    \I__10684\ : LocalMux
    port map (
            O => \N__50535\,
            I => data_in_frame_0_5
        );

    \I__10683\ : Odrv4
    port map (
            O => \N__50530\,
            I => data_in_frame_0_5
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__50525\,
            I => data_in_frame_0_5
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__50518\,
            I => data_in_frame_0_5
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__50515\,
            I => data_in_frame_0_5
        );

    \I__10679\ : InMux
    port map (
            O => \N__50500\,
            I => \N__50497\
        );

    \I__10678\ : LocalMux
    port map (
            O => \N__50497\,
            I => \N__50493\
        );

    \I__10677\ : InMux
    port map (
            O => \N__50496\,
            I => \N__50490\
        );

    \I__10676\ : Span4Mux_h
    port map (
            O => \N__50493\,
            I => \N__50487\
        );

    \I__10675\ : LocalMux
    port map (
            O => \N__50490\,
            I => \N__50482\
        );

    \I__10674\ : Span4Mux_h
    port map (
            O => \N__50487\,
            I => \N__50479\
        );

    \I__10673\ : InMux
    port map (
            O => \N__50486\,
            I => \N__50474\
        );

    \I__10672\ : InMux
    port map (
            O => \N__50485\,
            I => \N__50474\
        );

    \I__10671\ : Odrv12
    port map (
            O => \N__50482\,
            I => \c0.n33_adj_3088\
        );

    \I__10670\ : Odrv4
    port map (
            O => \N__50479\,
            I => \c0.n33_adj_3088\
        );

    \I__10669\ : LocalMux
    port map (
            O => \N__50474\,
            I => \c0.n33_adj_3088\
        );

    \I__10668\ : InMux
    port map (
            O => \N__50467\,
            I => \N__50464\
        );

    \I__10667\ : LocalMux
    port map (
            O => \N__50464\,
            I => \c0.n15_adj_3545\
        );

    \I__10666\ : InMux
    port map (
            O => \N__50461\,
            I => \N__50458\
        );

    \I__10665\ : LocalMux
    port map (
            O => \N__50458\,
            I => \N__50453\
        );

    \I__10664\ : InMux
    port map (
            O => \N__50457\,
            I => \N__50450\
        );

    \I__10663\ : CascadeMux
    port map (
            O => \N__50456\,
            I => \N__50447\
        );

    \I__10662\ : Span4Mux_v
    port map (
            O => \N__50453\,
            I => \N__50442\
        );

    \I__10661\ : LocalMux
    port map (
            O => \N__50450\,
            I => \N__50442\
        );

    \I__10660\ : InMux
    port map (
            O => \N__50447\,
            I => \N__50439\
        );

    \I__10659\ : Odrv4
    port map (
            O => \N__50442\,
            I => \c0.n24_adj_3013\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__50439\,
            I => \c0.n24_adj_3013\
        );

    \I__10657\ : CascadeMux
    port map (
            O => \N__50434\,
            I => \N__50429\
        );

    \I__10656\ : CascadeMux
    port map (
            O => \N__50433\,
            I => \N__50426\
        );

    \I__10655\ : CascadeMux
    port map (
            O => \N__50432\,
            I => \N__50422\
        );

    \I__10654\ : InMux
    port map (
            O => \N__50429\,
            I => \N__50419\
        );

    \I__10653\ : InMux
    port map (
            O => \N__50426\,
            I => \N__50412\
        );

    \I__10652\ : InMux
    port map (
            O => \N__50425\,
            I => \N__50412\
        );

    \I__10651\ : InMux
    port map (
            O => \N__50422\,
            I => \N__50412\
        );

    \I__10650\ : LocalMux
    port map (
            O => \N__50419\,
            I => \c0.data_in_frame_3_3\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__50412\,
            I => \c0.data_in_frame_3_3\
        );

    \I__10648\ : InMux
    port map (
            O => \N__50407\,
            I => \N__50402\
        );

    \I__10647\ : CascadeMux
    port map (
            O => \N__50406\,
            I => \N__50399\
        );

    \I__10646\ : InMux
    port map (
            O => \N__50405\,
            I => \N__50396\
        );

    \I__10645\ : LocalMux
    port map (
            O => \N__50402\,
            I => \N__50390\
        );

    \I__10644\ : InMux
    port map (
            O => \N__50399\,
            I => \N__50387\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__50396\,
            I => \N__50384\
        );

    \I__10642\ : InMux
    port map (
            O => \N__50395\,
            I => \N__50379\
        );

    \I__10641\ : InMux
    port map (
            O => \N__50394\,
            I => \N__50379\
        );

    \I__10640\ : InMux
    port map (
            O => \N__50393\,
            I => \N__50376\
        );

    \I__10639\ : Span4Mux_v
    port map (
            O => \N__50390\,
            I => \N__50371\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__50387\,
            I => \N__50371\
        );

    \I__10637\ : Odrv4
    port map (
            O => \N__50384\,
            I => \c0.data_in_frame_3_2\
        );

    \I__10636\ : LocalMux
    port map (
            O => \N__50379\,
            I => \c0.data_in_frame_3_2\
        );

    \I__10635\ : LocalMux
    port map (
            O => \N__50376\,
            I => \c0.data_in_frame_3_2\
        );

    \I__10634\ : Odrv4
    port map (
            O => \N__50371\,
            I => \c0.data_in_frame_3_2\
        );

    \I__10633\ : InMux
    port map (
            O => \N__50362\,
            I => \N__50356\
        );

    \I__10632\ : InMux
    port map (
            O => \N__50361\,
            I => \N__50353\
        );

    \I__10631\ : InMux
    port map (
            O => \N__50360\,
            I => \N__50350\
        );

    \I__10630\ : CascadeMux
    port map (
            O => \N__50359\,
            I => \N__50343\
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__50356\,
            I => \N__50340\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__50353\,
            I => \N__50336\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__50350\,
            I => \N__50333\
        );

    \I__10626\ : InMux
    port map (
            O => \N__50349\,
            I => \N__50329\
        );

    \I__10625\ : InMux
    port map (
            O => \N__50348\,
            I => \N__50326\
        );

    \I__10624\ : InMux
    port map (
            O => \N__50347\,
            I => \N__50321\
        );

    \I__10623\ : InMux
    port map (
            O => \N__50346\,
            I => \N__50321\
        );

    \I__10622\ : InMux
    port map (
            O => \N__50343\,
            I => \N__50318\
        );

    \I__10621\ : Span12Mux_v
    port map (
            O => \N__50340\,
            I => \N__50314\
        );

    \I__10620\ : InMux
    port map (
            O => \N__50339\,
            I => \N__50310\
        );

    \I__10619\ : Span4Mux_h
    port map (
            O => \N__50336\,
            I => \N__50305\
        );

    \I__10618\ : Span4Mux_v
    port map (
            O => \N__50333\,
            I => \N__50305\
        );

    \I__10617\ : InMux
    port map (
            O => \N__50332\,
            I => \N__50302\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__50329\,
            I => \N__50297\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__50326\,
            I => \N__50290\
        );

    \I__10614\ : LocalMux
    port map (
            O => \N__50321\,
            I => \N__50290\
        );

    \I__10613\ : LocalMux
    port map (
            O => \N__50318\,
            I => \N__50290\
        );

    \I__10612\ : InMux
    port map (
            O => \N__50317\,
            I => \N__50287\
        );

    \I__10611\ : Span12Mux_h
    port map (
            O => \N__50314\,
            I => \N__50282\
        );

    \I__10610\ : InMux
    port map (
            O => \N__50313\,
            I => \N__50279\
        );

    \I__10609\ : LocalMux
    port map (
            O => \N__50310\,
            I => \N__50272\
        );

    \I__10608\ : Span4Mux_h
    port map (
            O => \N__50305\,
            I => \N__50272\
        );

    \I__10607\ : LocalMux
    port map (
            O => \N__50302\,
            I => \N__50272\
        );

    \I__10606\ : InMux
    port map (
            O => \N__50301\,
            I => \N__50267\
        );

    \I__10605\ : InMux
    port map (
            O => \N__50300\,
            I => \N__50267\
        );

    \I__10604\ : Span4Mux_v
    port map (
            O => \N__50297\,
            I => \N__50260\
        );

    \I__10603\ : Span4Mux_v
    port map (
            O => \N__50290\,
            I => \N__50260\
        );

    \I__10602\ : LocalMux
    port map (
            O => \N__50287\,
            I => \N__50260\
        );

    \I__10601\ : InMux
    port map (
            O => \N__50286\,
            I => \N__50257\
        );

    \I__10600\ : InMux
    port map (
            O => \N__50285\,
            I => \N__50254\
        );

    \I__10599\ : Odrv12
    port map (
            O => \N__50282\,
            I => \data_out_frame_29__3__N_647\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__50279\,
            I => \data_out_frame_29__3__N_647\
        );

    \I__10597\ : Odrv4
    port map (
            O => \N__50272\,
            I => \data_out_frame_29__3__N_647\
        );

    \I__10596\ : LocalMux
    port map (
            O => \N__50267\,
            I => \data_out_frame_29__3__N_647\
        );

    \I__10595\ : Odrv4
    port map (
            O => \N__50260\,
            I => \data_out_frame_29__3__N_647\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__50257\,
            I => \data_out_frame_29__3__N_647\
        );

    \I__10593\ : LocalMux
    port map (
            O => \N__50254\,
            I => \data_out_frame_29__3__N_647\
        );

    \I__10592\ : InMux
    port map (
            O => \N__50239\,
            I => \N__50236\
        );

    \I__10591\ : LocalMux
    port map (
            O => \N__50236\,
            I => \N__50233\
        );

    \I__10590\ : Odrv12
    port map (
            O => \N__50233\,
            I => \c0.n29_adj_3216\
        );

    \I__10589\ : InMux
    port map (
            O => \N__50230\,
            I => \N__50227\
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__50227\,
            I => \N__50223\
        );

    \I__10587\ : InMux
    port map (
            O => \N__50226\,
            I => \N__50220\
        );

    \I__10586\ : Span4Mux_v
    port map (
            O => \N__50223\,
            I => \N__50217\
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__50220\,
            I => \N__50214\
        );

    \I__10584\ : Odrv4
    port map (
            O => \N__50217\,
            I => \c0.n78\
        );

    \I__10583\ : Odrv12
    port map (
            O => \N__50214\,
            I => \c0.n78\
        );

    \I__10582\ : InMux
    port map (
            O => \N__50209\,
            I => \N__50206\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__50206\,
            I => \N__50203\
        );

    \I__10580\ : Span4Mux_v
    port map (
            O => \N__50203\,
            I => \N__50200\
        );

    \I__10579\ : Sp12to4
    port map (
            O => \N__50200\,
            I => \N__50197\
        );

    \I__10578\ : Odrv12
    port map (
            O => \N__50197\,
            I => \c0.n37_adj_3215\
        );

    \I__10577\ : CascadeMux
    port map (
            O => \N__50194\,
            I => \c0.n29_adj_3216_cascade_\
        );

    \I__10576\ : InMux
    port map (
            O => \N__50191\,
            I => \N__50188\
        );

    \I__10575\ : LocalMux
    port map (
            O => \N__50188\,
            I => \c0.n44_adj_3217\
        );

    \I__10574\ : CascadeMux
    port map (
            O => \N__50185\,
            I => \c0.n8_adj_3066_cascade_\
        );

    \I__10573\ : InMux
    port map (
            O => \N__50182\,
            I => \N__50179\
        );

    \I__10572\ : LocalMux
    port map (
            O => \N__50179\,
            I => \N__50176\
        );

    \I__10571\ : Span4Mux_v
    port map (
            O => \N__50176\,
            I => \N__50172\
        );

    \I__10570\ : InMux
    port map (
            O => \N__50175\,
            I => \N__50169\
        );

    \I__10569\ : Span4Mux_h
    port map (
            O => \N__50172\,
            I => \N__50164\
        );

    \I__10568\ : LocalMux
    port map (
            O => \N__50169\,
            I => \N__50164\
        );

    \I__10567\ : Odrv4
    port map (
            O => \N__50164\,
            I => \c0.n19170\
        );

    \I__10566\ : CascadeMux
    port map (
            O => \N__50161\,
            I => \c0.n19170_cascade_\
        );

    \I__10565\ : CascadeMux
    port map (
            O => \N__50158\,
            I => \N__50154\
        );

    \I__10564\ : InMux
    port map (
            O => \N__50157\,
            I => \N__50151\
        );

    \I__10563\ : InMux
    port map (
            O => \N__50154\,
            I => \N__50146\
        );

    \I__10562\ : LocalMux
    port map (
            O => \N__50151\,
            I => \N__50143\
        );

    \I__10561\ : InMux
    port map (
            O => \N__50150\,
            I => \N__50140\
        );

    \I__10560\ : CascadeMux
    port map (
            O => \N__50149\,
            I => \N__50137\
        );

    \I__10559\ : LocalMux
    port map (
            O => \N__50146\,
            I => \N__50134\
        );

    \I__10558\ : Span4Mux_v
    port map (
            O => \N__50143\,
            I => \N__50129\
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__50140\,
            I => \N__50129\
        );

    \I__10556\ : InMux
    port map (
            O => \N__50137\,
            I => \N__50126\
        );

    \I__10555\ : Span4Mux_v
    port map (
            O => \N__50134\,
            I => \N__50123\
        );

    \I__10554\ : Span4Mux_h
    port map (
            O => \N__50129\,
            I => \N__50120\
        );

    \I__10553\ : LocalMux
    port map (
            O => \N__50126\,
            I => \c0.data_in_frame_8_2\
        );

    \I__10552\ : Odrv4
    port map (
            O => \N__50123\,
            I => \c0.data_in_frame_8_2\
        );

    \I__10551\ : Odrv4
    port map (
            O => \N__50120\,
            I => \c0.data_in_frame_8_2\
        );

    \I__10550\ : InMux
    port map (
            O => \N__50113\,
            I => \N__50110\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__50110\,
            I => \N__50105\
        );

    \I__10548\ : InMux
    port map (
            O => \N__50109\,
            I => \N__50102\
        );

    \I__10547\ : InMux
    port map (
            O => \N__50108\,
            I => \N__50099\
        );

    \I__10546\ : Span4Mux_v
    port map (
            O => \N__50105\,
            I => \N__50092\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__50102\,
            I => \N__50092\
        );

    \I__10544\ : LocalMux
    port map (
            O => \N__50099\,
            I => \N__50092\
        );

    \I__10543\ : Span4Mux_h
    port map (
            O => \N__50092\,
            I => \N__50089\
        );

    \I__10542\ : Odrv4
    port map (
            O => \N__50089\,
            I => \c0.n21_adj_3053\
        );

    \I__10541\ : CascadeMux
    port map (
            O => \N__50086\,
            I => \N__50083\
        );

    \I__10540\ : InMux
    port map (
            O => \N__50083\,
            I => \N__50078\
        );

    \I__10539\ : InMux
    port map (
            O => \N__50082\,
            I => \N__50073\
        );

    \I__10538\ : CascadeMux
    port map (
            O => \N__50081\,
            I => \N__50070\
        );

    \I__10537\ : LocalMux
    port map (
            O => \N__50078\,
            I => \N__50067\
        );

    \I__10536\ : InMux
    port map (
            O => \N__50077\,
            I => \N__50064\
        );

    \I__10535\ : InMux
    port map (
            O => \N__50076\,
            I => \N__50060\
        );

    \I__10534\ : LocalMux
    port map (
            O => \N__50073\,
            I => \N__50057\
        );

    \I__10533\ : InMux
    port map (
            O => \N__50070\,
            I => \N__50054\
        );

    \I__10532\ : Span4Mux_v
    port map (
            O => \N__50067\,
            I => \N__50049\
        );

    \I__10531\ : LocalMux
    port map (
            O => \N__50064\,
            I => \N__50049\
        );

    \I__10530\ : InMux
    port map (
            O => \N__50063\,
            I => \N__50046\
        );

    \I__10529\ : LocalMux
    port map (
            O => \N__50060\,
            I => \N__50043\
        );

    \I__10528\ : Span4Mux_h
    port map (
            O => \N__50057\,
            I => \N__50038\
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__50054\,
            I => \N__50038\
        );

    \I__10526\ : Span4Mux_v
    port map (
            O => \N__50049\,
            I => \N__50033\
        );

    \I__10525\ : LocalMux
    port map (
            O => \N__50046\,
            I => \N__50033\
        );

    \I__10524\ : Span4Mux_h
    port map (
            O => \N__50043\,
            I => \N__50026\
        );

    \I__10523\ : Span4Mux_v
    port map (
            O => \N__50038\,
            I => \N__50026\
        );

    \I__10522\ : Span4Mux_h
    port map (
            O => \N__50033\,
            I => \N__50026\
        );

    \I__10521\ : Odrv4
    port map (
            O => \N__50026\,
            I => \c0.n21\
        );

    \I__10520\ : CascadeMux
    port map (
            O => \N__50023\,
            I => \N__50019\
        );

    \I__10519\ : InMux
    port map (
            O => \N__50022\,
            I => \N__50016\
        );

    \I__10518\ : InMux
    port map (
            O => \N__50019\,
            I => \N__50013\
        );

    \I__10517\ : LocalMux
    port map (
            O => \N__50016\,
            I => \N__50010\
        );

    \I__10516\ : LocalMux
    port map (
            O => \N__50013\,
            I => \c0.data_in_frame_5_4\
        );

    \I__10515\ : Odrv4
    port map (
            O => \N__50010\,
            I => \c0.data_in_frame_5_4\
        );

    \I__10514\ : CascadeMux
    port map (
            O => \N__50005\,
            I => \N__50001\
        );

    \I__10513\ : InMux
    port map (
            O => \N__50004\,
            I => \N__49998\
        );

    \I__10512\ : InMux
    port map (
            O => \N__50001\,
            I => \N__49995\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__49998\,
            I => \c0.n25\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__49995\,
            I => \c0.n25\
        );

    \I__10509\ : InMux
    port map (
            O => \N__49990\,
            I => \N__49987\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__49987\,
            I => \c0.n89\
        );

    \I__10507\ : CascadeMux
    port map (
            O => \N__49984\,
            I => \N__49981\
        );

    \I__10506\ : InMux
    port map (
            O => \N__49981\,
            I => \N__49976\
        );

    \I__10505\ : InMux
    port map (
            O => \N__49980\,
            I => \N__49971\
        );

    \I__10504\ : InMux
    port map (
            O => \N__49979\,
            I => \N__49968\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__49976\,
            I => \N__49965\
        );

    \I__10502\ : InMux
    port map (
            O => \N__49975\,
            I => \N__49960\
        );

    \I__10501\ : InMux
    port map (
            O => \N__49974\,
            I => \N__49960\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__49971\,
            I => \c0.data_in_frame_4_0\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__49968\,
            I => \c0.data_in_frame_4_0\
        );

    \I__10498\ : Odrv4
    port map (
            O => \N__49965\,
            I => \c0.data_in_frame_4_0\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__49960\,
            I => \c0.data_in_frame_4_0\
        );

    \I__10496\ : InMux
    port map (
            O => \N__49951\,
            I => \N__49948\
        );

    \I__10495\ : LocalMux
    port map (
            O => \N__49948\,
            I => \N__49945\
        );

    \I__10494\ : Span4Mux_v
    port map (
            O => \N__49945\,
            I => \N__49942\
        );

    \I__10493\ : Odrv4
    port map (
            O => \N__49942\,
            I => \c0.n17_adj_3113\
        );

    \I__10492\ : InMux
    port map (
            O => \N__49939\,
            I => \N__49936\
        );

    \I__10491\ : LocalMux
    port map (
            O => \N__49936\,
            I => \c0.n5_adj_3030\
        );

    \I__10490\ : CascadeMux
    port map (
            O => \N__49933\,
            I => \c0.n60_cascade_\
        );

    \I__10489\ : InMux
    port map (
            O => \N__49930\,
            I => \N__49927\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__49927\,
            I => \N__49924\
        );

    \I__10487\ : Odrv4
    port map (
            O => \N__49924\,
            I => \c0.n93\
        );

    \I__10486\ : InMux
    port map (
            O => \N__49921\,
            I => \N__49918\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__49918\,
            I => \N__49913\
        );

    \I__10484\ : InMux
    port map (
            O => \N__49917\,
            I => \N__49910\
        );

    \I__10483\ : InMux
    port map (
            O => \N__49916\,
            I => \N__49907\
        );

    \I__10482\ : Span4Mux_v
    port map (
            O => \N__49913\,
            I => \N__49903\
        );

    \I__10481\ : LocalMux
    port map (
            O => \N__49910\,
            I => \N__49900\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__49907\,
            I => \N__49897\
        );

    \I__10479\ : InMux
    port map (
            O => \N__49906\,
            I => \N__49894\
        );

    \I__10478\ : Span4Mux_v
    port map (
            O => \N__49903\,
            I => \N__49891\
        );

    \I__10477\ : Span4Mux_h
    port map (
            O => \N__49900\,
            I => \N__49886\
        );

    \I__10476\ : Span4Mux_h
    port map (
            O => \N__49897\,
            I => \N__49886\
        );

    \I__10475\ : LocalMux
    port map (
            O => \N__49894\,
            I => \c0.data_in_frame_6_1\
        );

    \I__10474\ : Odrv4
    port map (
            O => \N__49891\,
            I => \c0.data_in_frame_6_1\
        );

    \I__10473\ : Odrv4
    port map (
            O => \N__49886\,
            I => \c0.data_in_frame_6_1\
        );

    \I__10472\ : InMux
    port map (
            O => \N__49879\,
            I => \N__49876\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__49876\,
            I => \N__49872\
        );

    \I__10470\ : CascadeMux
    port map (
            O => \N__49875\,
            I => \N__49869\
        );

    \I__10469\ : Span4Mux_v
    port map (
            O => \N__49872\,
            I => \N__49866\
        );

    \I__10468\ : InMux
    port map (
            O => \N__49869\,
            I => \N__49863\
        );

    \I__10467\ : Odrv4
    port map (
            O => \N__49866\,
            I => \c0.n5_adj_3028\
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__49863\,
            I => \c0.n5_adj_3028\
        );

    \I__10465\ : InMux
    port map (
            O => \N__49858\,
            I => \N__49855\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__49855\,
            I => \N__49852\
        );

    \I__10463\ : Span4Mux_h
    port map (
            O => \N__49852\,
            I => \N__49848\
        );

    \I__10462\ : InMux
    port map (
            O => \N__49851\,
            I => \N__49844\
        );

    \I__10461\ : Span4Mux_v
    port map (
            O => \N__49848\,
            I => \N__49841\
        );

    \I__10460\ : InMux
    port map (
            O => \N__49847\,
            I => \N__49838\
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__49844\,
            I => \N__49835\
        );

    \I__10458\ : Odrv4
    port map (
            O => \N__49841\,
            I => \c0.n19443\
        );

    \I__10457\ : LocalMux
    port map (
            O => \N__49838\,
            I => \c0.n19443\
        );

    \I__10456\ : Odrv4
    port map (
            O => \N__49835\,
            I => \c0.n19443\
        );

    \I__10455\ : InMux
    port map (
            O => \N__49828\,
            I => \N__49825\
        );

    \I__10454\ : LocalMux
    port map (
            O => \N__49825\,
            I => \N__49822\
        );

    \I__10453\ : Span4Mux_v
    port map (
            O => \N__49822\,
            I => \N__49819\
        );

    \I__10452\ : Span4Mux_h
    port map (
            O => \N__49819\,
            I => \N__49816\
        );

    \I__10451\ : Odrv4
    port map (
            O => \N__49816\,
            I => \c0.n11687\
        );

    \I__10450\ : InMux
    port map (
            O => \N__49813\,
            I => \N__49810\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__49810\,
            I => \N__49806\
        );

    \I__10448\ : CascadeMux
    port map (
            O => \N__49809\,
            I => \N__49803\
        );

    \I__10447\ : Span4Mux_v
    port map (
            O => \N__49806\,
            I => \N__49799\
        );

    \I__10446\ : InMux
    port map (
            O => \N__49803\,
            I => \N__49794\
        );

    \I__10445\ : InMux
    port map (
            O => \N__49802\,
            I => \N__49794\
        );

    \I__10444\ : Odrv4
    port map (
            O => \N__49799\,
            I => \c0.n20313\
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__49794\,
            I => \c0.n20313\
        );

    \I__10442\ : InMux
    port map (
            O => \N__49789\,
            I => \N__49786\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__49786\,
            I => \N__49782\
        );

    \I__10440\ : CascadeMux
    port map (
            O => \N__49785\,
            I => \N__49778\
        );

    \I__10439\ : Span4Mux_h
    port map (
            O => \N__49782\,
            I => \N__49775\
        );

    \I__10438\ : InMux
    port map (
            O => \N__49781\,
            I => \N__49770\
        );

    \I__10437\ : InMux
    port map (
            O => \N__49778\,
            I => \N__49770\
        );

    \I__10436\ : Odrv4
    port map (
            O => \N__49775\,
            I => \c0.data_in_frame_26_5\
        );

    \I__10435\ : LocalMux
    port map (
            O => \N__49770\,
            I => \c0.data_in_frame_26_5\
        );

    \I__10434\ : InMux
    port map (
            O => \N__49765\,
            I => \N__49762\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__49762\,
            I => \N__49759\
        );

    \I__10432\ : Odrv4
    port map (
            O => \N__49759\,
            I => \c0.n17840\
        );

    \I__10431\ : InMux
    port map (
            O => \N__49756\,
            I => \N__49751\
        );

    \I__10430\ : InMux
    port map (
            O => \N__49755\,
            I => \N__49748\
        );

    \I__10429\ : InMux
    port map (
            O => \N__49754\,
            I => \N__49745\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__49751\,
            I => \N__49741\
        );

    \I__10427\ : LocalMux
    port map (
            O => \N__49748\,
            I => \N__49738\
        );

    \I__10426\ : LocalMux
    port map (
            O => \N__49745\,
            I => \N__49735\
        );

    \I__10425\ : CascadeMux
    port map (
            O => \N__49744\,
            I => \N__49731\
        );

    \I__10424\ : Span4Mux_v
    port map (
            O => \N__49741\,
            I => \N__49723\
        );

    \I__10423\ : Span4Mux_v
    port map (
            O => \N__49738\,
            I => \N__49723\
        );

    \I__10422\ : Span4Mux_v
    port map (
            O => \N__49735\,
            I => \N__49723\
        );

    \I__10421\ : InMux
    port map (
            O => \N__49734\,
            I => \N__49720\
        );

    \I__10420\ : InMux
    port map (
            O => \N__49731\,
            I => \N__49717\
        );

    \I__10419\ : InMux
    port map (
            O => \N__49730\,
            I => \N__49714\
        );

    \I__10418\ : Span4Mux_h
    port map (
            O => \N__49723\,
            I => \N__49711\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__49720\,
            I => \N__49706\
        );

    \I__10416\ : LocalMux
    port map (
            O => \N__49717\,
            I => \N__49706\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__49714\,
            I => data_in_3_0
        );

    \I__10414\ : Odrv4
    port map (
            O => \N__49711\,
            I => data_in_3_0
        );

    \I__10413\ : Odrv12
    port map (
            O => \N__49706\,
            I => data_in_3_0
        );

    \I__10412\ : InMux
    port map (
            O => \N__49699\,
            I => \N__49696\
        );

    \I__10411\ : LocalMux
    port map (
            O => \N__49696\,
            I => \N__49693\
        );

    \I__10410\ : Span4Mux_v
    port map (
            O => \N__49693\,
            I => \N__49688\
        );

    \I__10409\ : InMux
    port map (
            O => \N__49692\,
            I => \N__49683\
        );

    \I__10408\ : InMux
    port map (
            O => \N__49691\,
            I => \N__49683\
        );

    \I__10407\ : Odrv4
    port map (
            O => \N__49688\,
            I => \c0.n12_adj_3498\
        );

    \I__10406\ : LocalMux
    port map (
            O => \N__49683\,
            I => \c0.n12_adj_3498\
        );

    \I__10405\ : CascadeMux
    port map (
            O => \N__49678\,
            I => \N__49673\
        );

    \I__10404\ : InMux
    port map (
            O => \N__49677\,
            I => \N__49669\
        );

    \I__10403\ : InMux
    port map (
            O => \N__49676\,
            I => \N__49666\
        );

    \I__10402\ : InMux
    port map (
            O => \N__49673\,
            I => \N__49662\
        );

    \I__10401\ : InMux
    port map (
            O => \N__49672\,
            I => \N__49659\
        );

    \I__10400\ : LocalMux
    port map (
            O => \N__49669\,
            I => \N__49656\
        );

    \I__10399\ : LocalMux
    port map (
            O => \N__49666\,
            I => \N__49652\
        );

    \I__10398\ : InMux
    port map (
            O => \N__49665\,
            I => \N__49649\
        );

    \I__10397\ : LocalMux
    port map (
            O => \N__49662\,
            I => \N__49644\
        );

    \I__10396\ : LocalMux
    port map (
            O => \N__49659\,
            I => \N__49644\
        );

    \I__10395\ : Span4Mux_v
    port map (
            O => \N__49656\,
            I => \N__49641\
        );

    \I__10394\ : InMux
    port map (
            O => \N__49655\,
            I => \N__49638\
        );

    \I__10393\ : Span4Mux_h
    port map (
            O => \N__49652\,
            I => \N__49633\
        );

    \I__10392\ : LocalMux
    port map (
            O => \N__49649\,
            I => \N__49633\
        );

    \I__10391\ : Span4Mux_v
    port map (
            O => \N__49644\,
            I => \N__49630\
        );

    \I__10390\ : Span4Mux_v
    port map (
            O => \N__49641\,
            I => \N__49627\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__49638\,
            I => \N__49624\
        );

    \I__10388\ : Span4Mux_h
    port map (
            O => \N__49633\,
            I => \N__49619\
        );

    \I__10387\ : Span4Mux_v
    port map (
            O => \N__49630\,
            I => \N__49619\
        );

    \I__10386\ : Span4Mux_v
    port map (
            O => \N__49627\,
            I => \N__49615\
        );

    \I__10385\ : Span4Mux_h
    port map (
            O => \N__49624\,
            I => \N__49612\
        );

    \I__10384\ : Span4Mux_v
    port map (
            O => \N__49619\,
            I => \N__49609\
        );

    \I__10383\ : InMux
    port map (
            O => \N__49618\,
            I => \N__49606\
        );

    \I__10382\ : Odrv4
    port map (
            O => \N__49615\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__10381\ : Odrv4
    port map (
            O => \N__49612\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__10380\ : Odrv4
    port map (
            O => \N__49609\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__10379\ : LocalMux
    port map (
            O => \N__49606\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__10378\ : SRMux
    port map (
            O => \N__49597\,
            I => \N__49594\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__49594\,
            I => \N__49591\
        );

    \I__10376\ : Sp12to4
    port map (
            O => \N__49591\,
            I => \N__49588\
        );

    \I__10375\ : Span12Mux_s7_v
    port map (
            O => \N__49588\,
            I => \N__49585\
        );

    \I__10374\ : Odrv12
    port map (
            O => \N__49585\,
            I => \c0.n6_adj_3149\
        );

    \I__10373\ : CascadeMux
    port map (
            O => \N__49582\,
            I => \N__49578\
        );

    \I__10372\ : CascadeMux
    port map (
            O => \N__49581\,
            I => \N__49574\
        );

    \I__10371\ : InMux
    port map (
            O => \N__49578\,
            I => \N__49571\
        );

    \I__10370\ : InMux
    port map (
            O => \N__49577\,
            I => \N__49566\
        );

    \I__10369\ : InMux
    port map (
            O => \N__49574\,
            I => \N__49566\
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__49571\,
            I => \N__49563\
        );

    \I__10367\ : LocalMux
    port map (
            O => \N__49566\,
            I => \N__49560\
        );

    \I__10366\ : Span4Mux_h
    port map (
            O => \N__49563\,
            I => \N__49553\
        );

    \I__10365\ : Span4Mux_v
    port map (
            O => \N__49560\,
            I => \N__49553\
        );

    \I__10364\ : InMux
    port map (
            O => \N__49559\,
            I => \N__49548\
        );

    \I__10363\ : InMux
    port map (
            O => \N__49558\,
            I => \N__49548\
        );

    \I__10362\ : Odrv4
    port map (
            O => \N__49553\,
            I => \c0.data_in_frame_8_6\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__49548\,
            I => \c0.data_in_frame_8_6\
        );

    \I__10360\ : InMux
    port map (
            O => \N__49543\,
            I => \N__49540\
        );

    \I__10359\ : LocalMux
    port map (
            O => \N__49540\,
            I => \N__49537\
        );

    \I__10358\ : Span4Mux_h
    port map (
            O => \N__49537\,
            I => \N__49532\
        );

    \I__10357\ : InMux
    port map (
            O => \N__49536\,
            I => \N__49527\
        );

    \I__10356\ : InMux
    port map (
            O => \N__49535\,
            I => \N__49527\
        );

    \I__10355\ : Odrv4
    port map (
            O => \N__49532\,
            I => \c0.n11936\
        );

    \I__10354\ : LocalMux
    port map (
            O => \N__49527\,
            I => \c0.n11936\
        );

    \I__10353\ : CascadeMux
    port map (
            O => \N__49522\,
            I => \N__49519\
        );

    \I__10352\ : InMux
    port map (
            O => \N__49519\,
            I => \N__49516\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__49516\,
            I => \N__49513\
        );

    \I__10350\ : Span4Mux_h
    port map (
            O => \N__49513\,
            I => \N__49510\
        );

    \I__10349\ : Odrv4
    port map (
            O => \N__49510\,
            I => \c0.n12_adj_3141\
        );

    \I__10348\ : InMux
    port map (
            O => \N__49507\,
            I => \N__49502\
        );

    \I__10347\ : InMux
    port map (
            O => \N__49506\,
            I => \N__49499\
        );

    \I__10346\ : InMux
    port map (
            O => \N__49505\,
            I => \N__49495\
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__49502\,
            I => \N__49492\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__49499\,
            I => \N__49488\
        );

    \I__10343\ : InMux
    port map (
            O => \N__49498\,
            I => \N__49484\
        );

    \I__10342\ : LocalMux
    port map (
            O => \N__49495\,
            I => \N__49479\
        );

    \I__10341\ : Span4Mux_v
    port map (
            O => \N__49492\,
            I => \N__49479\
        );

    \I__10340\ : InMux
    port map (
            O => \N__49491\,
            I => \N__49476\
        );

    \I__10339\ : Span4Mux_v
    port map (
            O => \N__49488\,
            I => \N__49473\
        );

    \I__10338\ : InMux
    port map (
            O => \N__49487\,
            I => \N__49470\
        );

    \I__10337\ : LocalMux
    port map (
            O => \N__49484\,
            I => data_in_frame_24_6
        );

    \I__10336\ : Odrv4
    port map (
            O => \N__49479\,
            I => data_in_frame_24_6
        );

    \I__10335\ : LocalMux
    port map (
            O => \N__49476\,
            I => data_in_frame_24_6
        );

    \I__10334\ : Odrv4
    port map (
            O => \N__49473\,
            I => data_in_frame_24_6
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__49470\,
            I => data_in_frame_24_6
        );

    \I__10332\ : InMux
    port map (
            O => \N__49459\,
            I => \N__49455\
        );

    \I__10331\ : InMux
    port map (
            O => \N__49458\,
            I => \N__49451\
        );

    \I__10330\ : LocalMux
    port map (
            O => \N__49455\,
            I => \N__49448\
        );

    \I__10329\ : InMux
    port map (
            O => \N__49454\,
            I => \N__49445\
        );

    \I__10328\ : LocalMux
    port map (
            O => \N__49451\,
            I => \N__49441\
        );

    \I__10327\ : Span4Mux_v
    port map (
            O => \N__49448\,
            I => \N__49436\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__49445\,
            I => \N__49436\
        );

    \I__10325\ : InMux
    port map (
            O => \N__49444\,
            I => \N__49432\
        );

    \I__10324\ : Span4Mux_h
    port map (
            O => \N__49441\,
            I => \N__49429\
        );

    \I__10323\ : Span4Mux_h
    port map (
            O => \N__49436\,
            I => \N__49426\
        );

    \I__10322\ : InMux
    port map (
            O => \N__49435\,
            I => \N__49423\
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__49432\,
            I => data_in_frame_24_4
        );

    \I__10320\ : Odrv4
    port map (
            O => \N__49429\,
            I => data_in_frame_24_4
        );

    \I__10319\ : Odrv4
    port map (
            O => \N__49426\,
            I => data_in_frame_24_4
        );

    \I__10318\ : LocalMux
    port map (
            O => \N__49423\,
            I => data_in_frame_24_4
        );

    \I__10317\ : CascadeMux
    port map (
            O => \N__49414\,
            I => \c0.n19465_cascade_\
        );

    \I__10316\ : InMux
    port map (
            O => \N__49411\,
            I => \N__49408\
        );

    \I__10315\ : LocalMux
    port map (
            O => \N__49408\,
            I => \N__49405\
        );

    \I__10314\ : Odrv4
    port map (
            O => \N__49405\,
            I => \c0.n17\
        );

    \I__10313\ : InMux
    port map (
            O => \N__49402\,
            I => \N__49398\
        );

    \I__10312\ : InMux
    port map (
            O => \N__49401\,
            I => \N__49393\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__49398\,
            I => \N__49390\
        );

    \I__10310\ : InMux
    port map (
            O => \N__49397\,
            I => \N__49387\
        );

    \I__10309\ : InMux
    port map (
            O => \N__49396\,
            I => \N__49384\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__49393\,
            I => \c0.n21044\
        );

    \I__10307\ : Odrv4
    port map (
            O => \N__49390\,
            I => \c0.n21044\
        );

    \I__10306\ : LocalMux
    port map (
            O => \N__49387\,
            I => \c0.n21044\
        );

    \I__10305\ : LocalMux
    port map (
            O => \N__49384\,
            I => \c0.n21044\
        );

    \I__10304\ : InMux
    port map (
            O => \N__49375\,
            I => \N__49372\
        );

    \I__10303\ : LocalMux
    port map (
            O => \N__49372\,
            I => \N__49368\
        );

    \I__10302\ : InMux
    port map (
            O => \N__49371\,
            I => \N__49365\
        );

    \I__10301\ : Span4Mux_h
    port map (
            O => \N__49368\,
            I => \N__49362\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__49365\,
            I => \c0.n19703\
        );

    \I__10299\ : Odrv4
    port map (
            O => \N__49362\,
            I => \c0.n19703\
        );

    \I__10298\ : CascadeMux
    port map (
            O => \N__49357\,
            I => \c0.n19703_cascade_\
        );

    \I__10297\ : InMux
    port map (
            O => \N__49354\,
            I => \N__49351\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__49351\,
            I => \c0.n44_adj_3278\
        );

    \I__10295\ : CascadeMux
    port map (
            O => \N__49348\,
            I => \N__49343\
        );

    \I__10294\ : InMux
    port map (
            O => \N__49347\,
            I => \N__49340\
        );

    \I__10293\ : InMux
    port map (
            O => \N__49346\,
            I => \N__49337\
        );

    \I__10292\ : InMux
    port map (
            O => \N__49343\,
            I => \N__49334\
        );

    \I__10291\ : LocalMux
    port map (
            O => \N__49340\,
            I => \N__49329\
        );

    \I__10290\ : LocalMux
    port map (
            O => \N__49337\,
            I => \N__49329\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__49334\,
            I => \N__49323\
        );

    \I__10288\ : Span4Mux_h
    port map (
            O => \N__49329\,
            I => \N__49320\
        );

    \I__10287\ : InMux
    port map (
            O => \N__49328\,
            I => \N__49317\
        );

    \I__10286\ : InMux
    port map (
            O => \N__49327\,
            I => \N__49312\
        );

    \I__10285\ : InMux
    port map (
            O => \N__49326\,
            I => \N__49312\
        );

    \I__10284\ : Odrv4
    port map (
            O => \N__49323\,
            I => \c0.data_in_frame_25_1\
        );

    \I__10283\ : Odrv4
    port map (
            O => \N__49320\,
            I => \c0.data_in_frame_25_1\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__49317\,
            I => \c0.data_in_frame_25_1\
        );

    \I__10281\ : LocalMux
    port map (
            O => \N__49312\,
            I => \c0.data_in_frame_25_1\
        );

    \I__10280\ : CascadeMux
    port map (
            O => \N__49303\,
            I => \N__49298\
        );

    \I__10279\ : InMux
    port map (
            O => \N__49302\,
            I => \N__49295\
        );

    \I__10278\ : InMux
    port map (
            O => \N__49301\,
            I => \N__49292\
        );

    \I__10277\ : InMux
    port map (
            O => \N__49298\,
            I => \N__49289\
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__49295\,
            I => \N__49285\
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__49292\,
            I => \N__49282\
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__49289\,
            I => \N__49279\
        );

    \I__10273\ : InMux
    port map (
            O => \N__49288\,
            I => \N__49276\
        );

    \I__10272\ : Span4Mux_h
    port map (
            O => \N__49285\,
            I => \N__49269\
        );

    \I__10271\ : Span4Mux_v
    port map (
            O => \N__49282\,
            I => \N__49269\
        );

    \I__10270\ : Span4Mux_h
    port map (
            O => \N__49279\,
            I => \N__49269\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__49276\,
            I => \N__49266\
        );

    \I__10268\ : Odrv4
    port map (
            O => \N__49269\,
            I => \c0.n18377\
        );

    \I__10267\ : Odrv4
    port map (
            O => \N__49266\,
            I => \c0.n18377\
        );

    \I__10266\ : InMux
    port map (
            O => \N__49261\,
            I => \N__49252\
        );

    \I__10265\ : InMux
    port map (
            O => \N__49260\,
            I => \N__49252\
        );

    \I__10264\ : InMux
    port map (
            O => \N__49259\,
            I => \N__49249\
        );

    \I__10263\ : InMux
    port map (
            O => \N__49258\,
            I => \N__49246\
        );

    \I__10262\ : InMux
    port map (
            O => \N__49257\,
            I => \N__49243\
        );

    \I__10261\ : LocalMux
    port map (
            O => \N__49252\,
            I => \N__49240\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__49249\,
            I => \c0.data_in_frame_25_2\
        );

    \I__10259\ : LocalMux
    port map (
            O => \N__49246\,
            I => \c0.data_in_frame_25_2\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__49243\,
            I => \c0.data_in_frame_25_2\
        );

    \I__10257\ : Odrv4
    port map (
            O => \N__49240\,
            I => \c0.data_in_frame_25_2\
        );

    \I__10256\ : InMux
    port map (
            O => \N__49231\,
            I => \N__49222\
        );

    \I__10255\ : InMux
    port map (
            O => \N__49230\,
            I => \N__49222\
        );

    \I__10254\ : InMux
    port map (
            O => \N__49229\,
            I => \N__49219\
        );

    \I__10253\ : InMux
    port map (
            O => \N__49228\,
            I => \N__49214\
        );

    \I__10252\ : InMux
    port map (
            O => \N__49227\,
            I => \N__49214\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__49222\,
            I => \N__49210\
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__49219\,
            I => \N__49205\
        );

    \I__10249\ : LocalMux
    port map (
            O => \N__49214\,
            I => \N__49205\
        );

    \I__10248\ : CascadeMux
    port map (
            O => \N__49213\,
            I => \N__49202\
        );

    \I__10247\ : Span4Mux_v
    port map (
            O => \N__49210\,
            I => \N__49199\
        );

    \I__10246\ : Span4Mux_v
    port map (
            O => \N__49205\,
            I => \N__49196\
        );

    \I__10245\ : InMux
    port map (
            O => \N__49202\,
            I => \N__49193\
        );

    \I__10244\ : Span4Mux_h
    port map (
            O => \N__49199\,
            I => \N__49188\
        );

    \I__10243\ : Span4Mux_v
    port map (
            O => \N__49196\,
            I => \N__49188\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__49193\,
            I => \c0.data_in_frame_25_3\
        );

    \I__10241\ : Odrv4
    port map (
            O => \N__49188\,
            I => \c0.data_in_frame_25_3\
        );

    \I__10240\ : CascadeMux
    port map (
            O => \N__49183\,
            I => \N__49179\
        );

    \I__10239\ : CascadeMux
    port map (
            O => \N__49182\,
            I => \N__49175\
        );

    \I__10238\ : InMux
    port map (
            O => \N__49179\,
            I => \N__49172\
        );

    \I__10237\ : InMux
    port map (
            O => \N__49178\,
            I => \N__49169\
        );

    \I__10236\ : InMux
    port map (
            O => \N__49175\,
            I => \N__49166\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__49172\,
            I => \N__49161\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__49169\,
            I => \N__49161\
        );

    \I__10233\ : LocalMux
    port map (
            O => \N__49166\,
            I => \N__49155\
        );

    \I__10232\ : Span4Mux_h
    port map (
            O => \N__49161\,
            I => \N__49155\
        );

    \I__10231\ : InMux
    port map (
            O => \N__49160\,
            I => \N__49152\
        );

    \I__10230\ : Odrv4
    port map (
            O => \N__49155\,
            I => \c0.n19400\
        );

    \I__10229\ : LocalMux
    port map (
            O => \N__49152\,
            I => \c0.n19400\
        );

    \I__10228\ : InMux
    port map (
            O => \N__49147\,
            I => \N__49144\
        );

    \I__10227\ : LocalMux
    port map (
            O => \N__49144\,
            I => \N__49140\
        );

    \I__10226\ : InMux
    port map (
            O => \N__49143\,
            I => \N__49137\
        );

    \I__10225\ : Span4Mux_h
    port map (
            O => \N__49140\,
            I => \N__49133\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__49137\,
            I => \N__49130\
        );

    \I__10223\ : InMux
    port map (
            O => \N__49136\,
            I => \N__49127\
        );

    \I__10222\ : Span4Mux_v
    port map (
            O => \N__49133\,
            I => \N__49124\
        );

    \I__10221\ : Span4Mux_h
    port map (
            O => \N__49130\,
            I => \N__49121\
        );

    \I__10220\ : LocalMux
    port map (
            O => \N__49127\,
            I => \N__49118\
        );

    \I__10219\ : Odrv4
    port map (
            O => \N__49124\,
            I => \c0.n12134\
        );

    \I__10218\ : Odrv4
    port map (
            O => \N__49121\,
            I => \c0.n12134\
        );

    \I__10217\ : Odrv12
    port map (
            O => \N__49118\,
            I => \c0.n12134\
        );

    \I__10216\ : InMux
    port map (
            O => \N__49111\,
            I => \N__49108\
        );

    \I__10215\ : LocalMux
    port map (
            O => \N__49108\,
            I => \c0.n58_adj_3381\
        );

    \I__10214\ : InMux
    port map (
            O => \N__49105\,
            I => \N__49102\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__49102\,
            I => \N__49099\
        );

    \I__10212\ : Span4Mux_v
    port map (
            O => \N__49099\,
            I => \N__49095\
        );

    \I__10211\ : InMux
    port map (
            O => \N__49098\,
            I => \N__49092\
        );

    \I__10210\ : Odrv4
    port map (
            O => \N__49095\,
            I => \c0.n43_adj_3330\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__49092\,
            I => \c0.n43_adj_3330\
        );

    \I__10208\ : InMux
    port map (
            O => \N__49087\,
            I => \N__49084\
        );

    \I__10207\ : LocalMux
    port map (
            O => \N__49084\,
            I => \c0.n50_adj_3331\
        );

    \I__10206\ : InMux
    port map (
            O => \N__49081\,
            I => \N__49076\
        );

    \I__10205\ : InMux
    port map (
            O => \N__49080\,
            I => \N__49073\
        );

    \I__10204\ : InMux
    port map (
            O => \N__49079\,
            I => \N__49070\
        );

    \I__10203\ : LocalMux
    port map (
            O => \N__49076\,
            I => \N__49065\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__49073\,
            I => \N__49062\
        );

    \I__10201\ : LocalMux
    port map (
            O => \N__49070\,
            I => \N__49059\
        );

    \I__10200\ : InMux
    port map (
            O => \N__49069\,
            I => \N__49056\
        );

    \I__10199\ : InMux
    port map (
            O => \N__49068\,
            I => \N__49053\
        );

    \I__10198\ : Span4Mux_v
    port map (
            O => \N__49065\,
            I => \N__49050\
        );

    \I__10197\ : Span4Mux_v
    port map (
            O => \N__49062\,
            I => \N__49045\
        );

    \I__10196\ : Span4Mux_h
    port map (
            O => \N__49059\,
            I => \N__49045\
        );

    \I__10195\ : LocalMux
    port map (
            O => \N__49056\,
            I => \N__49040\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__49053\,
            I => \N__49040\
        );

    \I__10193\ : Span4Mux_h
    port map (
            O => \N__49050\,
            I => \N__49037\
        );

    \I__10192\ : Span4Mux_v
    port map (
            O => \N__49045\,
            I => \N__49034\
        );

    \I__10191\ : Span4Mux_h
    port map (
            O => \N__49040\,
            I => \N__49031\
        );

    \I__10190\ : Odrv4
    port map (
            O => \N__49037\,
            I => \c0.n35_adj_3266\
        );

    \I__10189\ : Odrv4
    port map (
            O => \N__49034\,
            I => \c0.n35_adj_3266\
        );

    \I__10188\ : Odrv4
    port map (
            O => \N__49031\,
            I => \c0.n35_adj_3266\
        );

    \I__10187\ : InMux
    port map (
            O => \N__49024\,
            I => \N__49021\
        );

    \I__10186\ : LocalMux
    port map (
            O => \N__49021\,
            I => \N__49018\
        );

    \I__10185\ : Span4Mux_v
    port map (
            O => \N__49018\,
            I => \N__49014\
        );

    \I__10184\ : InMux
    port map (
            O => \N__49017\,
            I => \N__49011\
        );

    \I__10183\ : Odrv4
    port map (
            O => \N__49014\,
            I => \c0.n33_adj_3097\
        );

    \I__10182\ : LocalMux
    port map (
            O => \N__49011\,
            I => \c0.n33_adj_3097\
        );

    \I__10181\ : CascadeMux
    port map (
            O => \N__49006\,
            I => \N__49003\
        );

    \I__10180\ : InMux
    port map (
            O => \N__49003\,
            I => \N__49000\
        );

    \I__10179\ : LocalMux
    port map (
            O => \N__49000\,
            I => \N__48997\
        );

    \I__10178\ : Span4Mux_v
    port map (
            O => \N__48997\,
            I => \N__48994\
        );

    \I__10177\ : Odrv4
    port map (
            O => \N__48994\,
            I => \c0.n9_adj_3240\
        );

    \I__10176\ : InMux
    port map (
            O => \N__48991\,
            I => \N__48988\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__48988\,
            I => \N__48985\
        );

    \I__10174\ : Span4Mux_v
    port map (
            O => \N__48985\,
            I => \N__48982\
        );

    \I__10173\ : Odrv4
    port map (
            O => \N__48982\,
            I => \c0.n20112\
        );

    \I__10172\ : InMux
    port map (
            O => \N__48979\,
            I => \N__48976\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__48976\,
            I => \N__48973\
        );

    \I__10170\ : Span4Mux_h
    port map (
            O => \N__48973\,
            I => \N__48970\
        );

    \I__10169\ : Span4Mux_v
    port map (
            O => \N__48970\,
            I => \N__48967\
        );

    \I__10168\ : Odrv4
    port map (
            O => \N__48967\,
            I => \c0.n32_adj_3236\
        );

    \I__10167\ : InMux
    port map (
            O => \N__48964\,
            I => \N__48961\
        );

    \I__10166\ : LocalMux
    port map (
            O => \N__48961\,
            I => \N__48957\
        );

    \I__10165\ : InMux
    port map (
            O => \N__48960\,
            I => \N__48954\
        );

    \I__10164\ : Span4Mux_v
    port map (
            O => \N__48957\,
            I => \N__48949\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__48954\,
            I => \N__48949\
        );

    \I__10162\ : Span4Mux_v
    port map (
            O => \N__48949\,
            I => \N__48946\
        );

    \I__10161\ : Odrv4
    port map (
            O => \N__48946\,
            I => \c0.n28_adj_3245\
        );

    \I__10160\ : CascadeMux
    port map (
            O => \N__48943\,
            I => \c0.n27_adj_3241_cascade_\
        );

    \I__10159\ : InMux
    port map (
            O => \N__48940\,
            I => \N__48937\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__48937\,
            I => \N__48934\
        );

    \I__10157\ : Span4Mux_v
    port map (
            O => \N__48934\,
            I => \N__48927\
        );

    \I__10156\ : InMux
    port map (
            O => \N__48933\,
            I => \N__48924\
        );

    \I__10155\ : InMux
    port map (
            O => \N__48932\,
            I => \N__48921\
        );

    \I__10154\ : InMux
    port map (
            O => \N__48931\,
            I => \N__48916\
        );

    \I__10153\ : InMux
    port map (
            O => \N__48930\,
            I => \N__48916\
        );

    \I__10152\ : Odrv4
    port map (
            O => \N__48927\,
            I => \c0.n13_adj_3244\
        );

    \I__10151\ : LocalMux
    port map (
            O => \N__48924\,
            I => \c0.n13_adj_3244\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__48921\,
            I => \c0.n13_adj_3244\
        );

    \I__10149\ : LocalMux
    port map (
            O => \N__48916\,
            I => \c0.n13_adj_3244\
        );

    \I__10148\ : InMux
    port map (
            O => \N__48907\,
            I => \N__48904\
        );

    \I__10147\ : LocalMux
    port map (
            O => \N__48904\,
            I => \c0.n19_adj_3135\
        );

    \I__10146\ : CascadeMux
    port map (
            O => \N__48901\,
            I => \c0.n19_adj_3135_cascade_\
        );

    \I__10145\ : InMux
    port map (
            O => \N__48898\,
            I => \N__48895\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__48895\,
            I => \N__48891\
        );

    \I__10143\ : InMux
    port map (
            O => \N__48894\,
            I => \N__48888\
        );

    \I__10142\ : Span4Mux_h
    port map (
            O => \N__48891\,
            I => \N__48885\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__48888\,
            I => \c0.n24_adj_3134\
        );

    \I__10140\ : Odrv4
    port map (
            O => \N__48885\,
            I => \c0.n24_adj_3134\
        );

    \I__10139\ : InMux
    port map (
            O => \N__48880\,
            I => \N__48877\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__48877\,
            I => \N__48873\
        );

    \I__10137\ : InMux
    port map (
            O => \N__48876\,
            I => \N__48870\
        );

    \I__10136\ : Span4Mux_v
    port map (
            O => \N__48873\,
            I => \N__48864\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__48870\,
            I => \N__48864\
        );

    \I__10134\ : InMux
    port map (
            O => \N__48869\,
            I => \N__48861\
        );

    \I__10133\ : Span4Mux_v
    port map (
            O => \N__48864\,
            I => \N__48855\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__48861\,
            I => \N__48855\
        );

    \I__10131\ : InMux
    port map (
            O => \N__48860\,
            I => \N__48852\
        );

    \I__10130\ : Span4Mux_h
    port map (
            O => \N__48855\,
            I => \N__48849\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__48852\,
            I => \c0.n86\
        );

    \I__10128\ : Odrv4
    port map (
            O => \N__48849\,
            I => \c0.n86\
        );

    \I__10127\ : CascadeMux
    port map (
            O => \N__48844\,
            I => \c0.n22_adj_3136_cascade_\
        );

    \I__10126\ : CascadeMux
    port map (
            O => \N__48841\,
            I => \c0.n11936_cascade_\
        );

    \I__10125\ : InMux
    port map (
            O => \N__48838\,
            I => \N__48834\
        );

    \I__10124\ : InMux
    port map (
            O => \N__48837\,
            I => \N__48831\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__48834\,
            I => \N__48826\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__48831\,
            I => \N__48823\
        );

    \I__10121\ : CascadeMux
    port map (
            O => \N__48830\,
            I => \N__48820\
        );

    \I__10120\ : InMux
    port map (
            O => \N__48829\,
            I => \N__48817\
        );

    \I__10119\ : Span4Mux_h
    port map (
            O => \N__48826\,
            I => \N__48814\
        );

    \I__10118\ : Span4Mux_h
    port map (
            O => \N__48823\,
            I => \N__48811\
        );

    \I__10117\ : InMux
    port map (
            O => \N__48820\,
            I => \N__48808\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__48817\,
            I => \N__48805\
        );

    \I__10115\ : Span4Mux_h
    port map (
            O => \N__48814\,
            I => \N__48802\
        );

    \I__10114\ : Span4Mux_h
    port map (
            O => \N__48811\,
            I => \N__48799\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__48808\,
            I => \c0.data_in_frame_27_4\
        );

    \I__10112\ : Odrv4
    port map (
            O => \N__48805\,
            I => \c0.data_in_frame_27_4\
        );

    \I__10111\ : Odrv4
    port map (
            O => \N__48802\,
            I => \c0.data_in_frame_27_4\
        );

    \I__10110\ : Odrv4
    port map (
            O => \N__48799\,
            I => \c0.data_in_frame_27_4\
        );

    \I__10109\ : InMux
    port map (
            O => \N__48790\,
            I => \N__48786\
        );

    \I__10108\ : InMux
    port map (
            O => \N__48789\,
            I => \N__48782\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__48786\,
            I => \N__48779\
        );

    \I__10106\ : CascadeMux
    port map (
            O => \N__48785\,
            I => \N__48775\
        );

    \I__10105\ : LocalMux
    port map (
            O => \N__48782\,
            I => \N__48772\
        );

    \I__10104\ : Span4Mux_v
    port map (
            O => \N__48779\,
            I => \N__48769\
        );

    \I__10103\ : CascadeMux
    port map (
            O => \N__48778\,
            I => \N__48766\
        );

    \I__10102\ : InMux
    port map (
            O => \N__48775\,
            I => \N__48763\
        );

    \I__10101\ : Span4Mux_h
    port map (
            O => \N__48772\,
            I => \N__48760\
        );

    \I__10100\ : Sp12to4
    port map (
            O => \N__48769\,
            I => \N__48757\
        );

    \I__10099\ : InMux
    port map (
            O => \N__48766\,
            I => \N__48754\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__48763\,
            I => \N__48751\
        );

    \I__10097\ : Span4Mux_v
    port map (
            O => \N__48760\,
            I => \N__48748\
        );

    \I__10096\ : Span12Mux_h
    port map (
            O => \N__48757\,
            I => \N__48743\
        );

    \I__10095\ : LocalMux
    port map (
            O => \N__48754\,
            I => \N__48743\
        );

    \I__10094\ : Odrv4
    port map (
            O => \N__48751\,
            I => \c0.data_in_frame_27_5\
        );

    \I__10093\ : Odrv4
    port map (
            O => \N__48748\,
            I => \c0.data_in_frame_27_5\
        );

    \I__10092\ : Odrv12
    port map (
            O => \N__48743\,
            I => \c0.data_in_frame_27_5\
        );

    \I__10091\ : InMux
    port map (
            O => \N__48736\,
            I => \N__48733\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__48733\,
            I => \N__48730\
        );

    \I__10089\ : Odrv4
    port map (
            O => \N__48730\,
            I => \c0.n17_adj_3318\
        );

    \I__10088\ : CascadeMux
    port map (
            O => \N__48727\,
            I => \c0.n32_adj_3057_cascade_\
        );

    \I__10087\ : InMux
    port map (
            O => \N__48724\,
            I => \N__48716\
        );

    \I__10086\ : InMux
    port map (
            O => \N__48723\,
            I => \N__48716\
        );

    \I__10085\ : InMux
    port map (
            O => \N__48722\,
            I => \N__48711\
        );

    \I__10084\ : InMux
    port map (
            O => \N__48721\,
            I => \N__48711\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__48716\,
            I => \N__48708\
        );

    \I__10082\ : LocalMux
    port map (
            O => \N__48711\,
            I => \N__48703\
        );

    \I__10081\ : Span4Mux_v
    port map (
            O => \N__48708\,
            I => \N__48703\
        );

    \I__10080\ : Span4Mux_v
    port map (
            O => \N__48703\,
            I => \N__48700\
        );

    \I__10079\ : Odrv4
    port map (
            O => \N__48700\,
            I => \c0.n33_adj_3289\
        );

    \I__10078\ : InMux
    port map (
            O => \N__48697\,
            I => \N__48694\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__48694\,
            I => \N__48691\
        );

    \I__10076\ : Odrv4
    port map (
            O => \N__48691\,
            I => \c0.n10_adj_3555\
        );

    \I__10075\ : CascadeMux
    port map (
            O => \N__48688\,
            I => \N__48685\
        );

    \I__10074\ : InMux
    port map (
            O => \N__48685\,
            I => \N__48682\
        );

    \I__10073\ : LocalMux
    port map (
            O => \N__48682\,
            I => \N__48679\
        );

    \I__10072\ : Span4Mux_v
    port map (
            O => \N__48679\,
            I => \N__48676\
        );

    \I__10071\ : Span4Mux_h
    port map (
            O => \N__48676\,
            I => \N__48673\
        );

    \I__10070\ : Sp12to4
    port map (
            O => \N__48673\,
            I => \N__48670\
        );

    \I__10069\ : Odrv12
    port map (
            O => \N__48670\,
            I => \c0.n4_adj_3522\
        );

    \I__10068\ : InMux
    port map (
            O => \N__48667\,
            I => \N__48661\
        );

    \I__10067\ : InMux
    port map (
            O => \N__48666\,
            I => \N__48661\
        );

    \I__10066\ : LocalMux
    port map (
            O => \N__48661\,
            I => \c0.n55_adj_3273\
        );

    \I__10065\ : InMux
    port map (
            O => \N__48658\,
            I => \N__48655\
        );

    \I__10064\ : LocalMux
    port map (
            O => \N__48655\,
            I => \N__48651\
        );

    \I__10063\ : InMux
    port map (
            O => \N__48654\,
            I => \N__48647\
        );

    \I__10062\ : Span4Mux_v
    port map (
            O => \N__48651\,
            I => \N__48644\
        );

    \I__10061\ : InMux
    port map (
            O => \N__48650\,
            I => \N__48641\
        );

    \I__10060\ : LocalMux
    port map (
            O => \N__48647\,
            I => \c0.n19514\
        );

    \I__10059\ : Odrv4
    port map (
            O => \N__48644\,
            I => \c0.n19514\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__48641\,
            I => \c0.n19514\
        );

    \I__10057\ : CascadeMux
    port map (
            O => \N__48634\,
            I => \c0.n20965_cascade_\
        );

    \I__10056\ : InMux
    port map (
            O => \N__48631\,
            I => \N__48628\
        );

    \I__10055\ : LocalMux
    port map (
            O => \N__48628\,
            I => \N__48625\
        );

    \I__10054\ : Span4Mux_h
    port map (
            O => \N__48625\,
            I => \N__48622\
        );

    \I__10053\ : Odrv4
    port map (
            O => \N__48622\,
            I => \c0.n40_adj_3323\
        );

    \I__10052\ : InMux
    port map (
            O => \N__48619\,
            I => \N__48614\
        );

    \I__10051\ : InMux
    port map (
            O => \N__48618\,
            I => \N__48611\
        );

    \I__10050\ : CascadeMux
    port map (
            O => \N__48617\,
            I => \N__48608\
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__48614\,
            I => \N__48605\
        );

    \I__10048\ : LocalMux
    port map (
            O => \N__48611\,
            I => \N__48602\
        );

    \I__10047\ : InMux
    port map (
            O => \N__48608\,
            I => \N__48599\
        );

    \I__10046\ : Span4Mux_v
    port map (
            O => \N__48605\,
            I => \N__48596\
        );

    \I__10045\ : Span4Mux_v
    port map (
            O => \N__48602\,
            I => \N__48592\
        );

    \I__10044\ : LocalMux
    port map (
            O => \N__48599\,
            I => \N__48587\
        );

    \I__10043\ : Span4Mux_v
    port map (
            O => \N__48596\,
            I => \N__48587\
        );

    \I__10042\ : InMux
    port map (
            O => \N__48595\,
            I => \N__48584\
        );

    \I__10041\ : Span4Mux_h
    port map (
            O => \N__48592\,
            I => \N__48581\
        );

    \I__10040\ : Odrv4
    port map (
            O => \N__48587\,
            I => \c0.data_in_frame_27_3\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__48584\,
            I => \c0.data_in_frame_27_3\
        );

    \I__10038\ : Odrv4
    port map (
            O => \N__48581\,
            I => \c0.data_in_frame_27_3\
        );

    \I__10037\ : CascadeMux
    port map (
            O => \N__48574\,
            I => \c0.n20336_cascade_\
        );

    \I__10036\ : InMux
    port map (
            O => \N__48571\,
            I => \N__48568\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__48568\,
            I => \N__48565\
        );

    \I__10034\ : Span4Mux_v
    port map (
            O => \N__48565\,
            I => \N__48562\
        );

    \I__10033\ : Odrv4
    port map (
            O => \N__48562\,
            I => \c0.n61_adj_3387\
        );

    \I__10032\ : InMux
    port map (
            O => \N__48559\,
            I => \N__48556\
        );

    \I__10031\ : LocalMux
    port map (
            O => \N__48556\,
            I => \N__48553\
        );

    \I__10030\ : Odrv4
    port map (
            O => \N__48553\,
            I => \c0.n63_adj_3391\
        );

    \I__10029\ : CascadeMux
    port map (
            O => \N__48550\,
            I => \c0.n21034_cascade_\
        );

    \I__10028\ : CascadeMux
    port map (
            O => \N__48547\,
            I => \c0.n35_adj_3274_cascade_\
        );

    \I__10027\ : InMux
    port map (
            O => \N__48544\,
            I => \N__48541\
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__48541\,
            I => \c0.n59\
        );

    \I__10025\ : InMux
    port map (
            O => \N__48538\,
            I => \N__48535\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__48535\,
            I => \N__48531\
        );

    \I__10023\ : InMux
    port map (
            O => \N__48534\,
            I => \N__48528\
        );

    \I__10022\ : Span4Mux_h
    port map (
            O => \N__48531\,
            I => \N__48524\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__48528\,
            I => \N__48521\
        );

    \I__10020\ : InMux
    port map (
            O => \N__48527\,
            I => \N__48518\
        );

    \I__10019\ : Odrv4
    port map (
            O => \N__48524\,
            I => \c0.n30_adj_3392\
        );

    \I__10018\ : Odrv12
    port map (
            O => \N__48521\,
            I => \c0.n30_adj_3392\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__48518\,
            I => \c0.n30_adj_3392\
        );

    \I__10016\ : InMux
    port map (
            O => \N__48511\,
            I => \N__48507\
        );

    \I__10015\ : InMux
    port map (
            O => \N__48510\,
            I => \N__48504\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__48507\,
            I => \N__48501\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__48504\,
            I => \N__48496\
        );

    \I__10012\ : Span4Mux_v
    port map (
            O => \N__48501\,
            I => \N__48496\
        );

    \I__10011\ : Span4Mux_v
    port map (
            O => \N__48496\,
            I => \N__48493\
        );

    \I__10010\ : Odrv4
    port map (
            O => \N__48493\,
            I => \c0.n21047\
        );

    \I__10009\ : InMux
    port map (
            O => \N__48490\,
            I => \N__48486\
        );

    \I__10008\ : InMux
    port map (
            O => \N__48489\,
            I => \N__48483\
        );

    \I__10007\ : LocalMux
    port map (
            O => \N__48486\,
            I => \N__48480\
        );

    \I__10006\ : LocalMux
    port map (
            O => \N__48483\,
            I => \N__48477\
        );

    \I__10005\ : Span4Mux_h
    port map (
            O => \N__48480\,
            I => \N__48474\
        );

    \I__10004\ : Span4Mux_v
    port map (
            O => \N__48477\,
            I => \N__48471\
        );

    \I__10003\ : Sp12to4
    port map (
            O => \N__48474\,
            I => \N__48468\
        );

    \I__10002\ : Span4Mux_v
    port map (
            O => \N__48471\,
            I => \N__48465\
        );

    \I__10001\ : Odrv12
    port map (
            O => \N__48468\,
            I => \c0.n12_adj_3049\
        );

    \I__10000\ : Odrv4
    port map (
            O => \N__48465\,
            I => \c0.n12_adj_3049\
        );

    \I__9999\ : InMux
    port map (
            O => \N__48460\,
            I => \N__48457\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__48457\,
            I => \N__48454\
        );

    \I__9997\ : Odrv12
    port map (
            O => \N__48454\,
            I => \c0.n91\
        );

    \I__9996\ : CascadeMux
    port map (
            O => \N__48451\,
            I => \N__48447\
        );

    \I__9995\ : InMux
    port map (
            O => \N__48450\,
            I => \N__48444\
        );

    \I__9994\ : InMux
    port map (
            O => \N__48447\,
            I => \N__48441\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__48444\,
            I => \c0.n35_adj_3274\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__48441\,
            I => \c0.n35_adj_3274\
        );

    \I__9991\ : InMux
    port map (
            O => \N__48436\,
            I => \N__48433\
        );

    \I__9990\ : LocalMux
    port map (
            O => \N__48433\,
            I => \N__48430\
        );

    \I__9989\ : Span4Mux_v
    port map (
            O => \N__48430\,
            I => \N__48426\
        );

    \I__9988\ : InMux
    port map (
            O => \N__48429\,
            I => \N__48423\
        );

    \I__9987\ : Span4Mux_h
    port map (
            O => \N__48426\,
            I => \N__48420\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__48423\,
            I => \N__48417\
        );

    \I__9985\ : Odrv4
    port map (
            O => \N__48420\,
            I => \c0.n17_adj_3451\
        );

    \I__9984\ : Odrv4
    port map (
            O => \N__48417\,
            I => \c0.n17_adj_3451\
        );

    \I__9983\ : InMux
    port map (
            O => \N__48412\,
            I => \N__48409\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__48409\,
            I => \N__48406\
        );

    \I__9981\ : Span4Mux_v
    port map (
            O => \N__48406\,
            I => \N__48403\
        );

    \I__9980\ : Span4Mux_h
    port map (
            O => \N__48403\,
            I => \N__48399\
        );

    \I__9979\ : InMux
    port map (
            O => \N__48402\,
            I => \N__48396\
        );

    \I__9978\ : Odrv4
    port map (
            O => \N__48399\,
            I => \c0.n20403\
        );

    \I__9977\ : LocalMux
    port map (
            O => \N__48396\,
            I => \c0.n20403\
        );

    \I__9976\ : InMux
    port map (
            O => \N__48391\,
            I => \N__48388\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__48388\,
            I => \c0.n22_adj_3450\
        );

    \I__9974\ : CascadeMux
    port map (
            O => \N__48385\,
            I => \c0.n24_adj_3427_cascade_\
        );

    \I__9973\ : InMux
    port map (
            O => \N__48382\,
            I => \N__48378\
        );

    \I__9972\ : InMux
    port map (
            O => \N__48381\,
            I => \N__48374\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__48378\,
            I => \N__48370\
        );

    \I__9970\ : InMux
    port map (
            O => \N__48377\,
            I => \N__48367\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__48374\,
            I => \N__48363\
        );

    \I__9968\ : InMux
    port map (
            O => \N__48373\,
            I => \N__48360\
        );

    \I__9967\ : Span4Mux_v
    port map (
            O => \N__48370\,
            I => \N__48355\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__48367\,
            I => \N__48355\
        );

    \I__9965\ : CascadeMux
    port map (
            O => \N__48366\,
            I => \N__48352\
        );

    \I__9964\ : Span4Mux_v
    port map (
            O => \N__48363\,
            I => \N__48345\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__48360\,
            I => \N__48345\
        );

    \I__9962\ : Span4Mux_h
    port map (
            O => \N__48355\,
            I => \N__48345\
        );

    \I__9961\ : InMux
    port map (
            O => \N__48352\,
            I => \N__48342\
        );

    \I__9960\ : Span4Mux_v
    port map (
            O => \N__48345\,
            I => \N__48339\
        );

    \I__9959\ : LocalMux
    port map (
            O => \N__48342\,
            I => \c0.data_in_frame_17_0\
        );

    \I__9958\ : Odrv4
    port map (
            O => \N__48339\,
            I => \c0.data_in_frame_17_0\
        );

    \I__9957\ : InMux
    port map (
            O => \N__48334\,
            I => \N__48330\
        );

    \I__9956\ : InMux
    port map (
            O => \N__48333\,
            I => \N__48327\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__48330\,
            I => \N__48322\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__48327\,
            I => \N__48319\
        );

    \I__9953\ : InMux
    port map (
            O => \N__48326\,
            I => \N__48314\
        );

    \I__9952\ : InMux
    port map (
            O => \N__48325\,
            I => \N__48314\
        );

    \I__9951\ : Span12Mux_v
    port map (
            O => \N__48322\,
            I => \N__48311\
        );

    \I__9950\ : Odrv4
    port map (
            O => \N__48319\,
            I => \c0.data_in_frame_13_1\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__48314\,
            I => \c0.data_in_frame_13_1\
        );

    \I__9948\ : Odrv12
    port map (
            O => \N__48311\,
            I => \c0.data_in_frame_13_1\
        );

    \I__9947\ : CascadeMux
    port map (
            O => \N__48304\,
            I => \c0.n18398_cascade_\
        );

    \I__9946\ : CascadeMux
    port map (
            O => \N__48301\,
            I => \c0.n37_adj_3390_cascade_\
        );

    \I__9945\ : InMux
    port map (
            O => \N__48298\,
            I => \N__48295\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__48295\,
            I => \c0.n37_adj_3390\
        );

    \I__9943\ : CascadeMux
    port map (
            O => \N__48292\,
            I => \c0.n60_adj_3368_cascade_\
        );

    \I__9942\ : InMux
    port map (
            O => \N__48289\,
            I => \N__48286\
        );

    \I__9941\ : LocalMux
    port map (
            O => \N__48286\,
            I => \c0.n51_adj_3376\
        );

    \I__9940\ : InMux
    port map (
            O => \N__48283\,
            I => \N__48280\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__48280\,
            I => \N__48276\
        );

    \I__9938\ : InMux
    port map (
            O => \N__48279\,
            I => \N__48273\
        );

    \I__9937\ : Span4Mux_v
    port map (
            O => \N__48276\,
            I => \N__48270\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__48273\,
            I => \c0.n19916\
        );

    \I__9935\ : Odrv4
    port map (
            O => \N__48270\,
            I => \c0.n19916\
        );

    \I__9934\ : InMux
    port map (
            O => \N__48265\,
            I => \N__48262\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__48262\,
            I => \N__48257\
        );

    \I__9932\ : InMux
    port map (
            O => \N__48261\,
            I => \N__48254\
        );

    \I__9931\ : InMux
    port map (
            O => \N__48260\,
            I => \N__48251\
        );

    \I__9930\ : Span4Mux_h
    port map (
            O => \N__48257\,
            I => \N__48248\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__48254\,
            I => \N__48243\
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__48251\,
            I => \N__48243\
        );

    \I__9927\ : Span4Mux_v
    port map (
            O => \N__48248\,
            I => \N__48240\
        );

    \I__9926\ : Span4Mux_v
    port map (
            O => \N__48243\,
            I => \N__48237\
        );

    \I__9925\ : Odrv4
    port map (
            O => \N__48240\,
            I => \c0.n18443\
        );

    \I__9924\ : Odrv4
    port map (
            O => \N__48237\,
            I => \c0.n18443\
        );

    \I__9923\ : InMux
    port map (
            O => \N__48232\,
            I => \N__48229\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__48229\,
            I => \c0.n39_adj_3334\
        );

    \I__9921\ : InMux
    port map (
            O => \N__48226\,
            I => \N__48220\
        );

    \I__9920\ : InMux
    port map (
            O => \N__48225\,
            I => \N__48220\
        );

    \I__9919\ : LocalMux
    port map (
            O => \N__48220\,
            I => \N__48216\
        );

    \I__9918\ : CascadeMux
    port map (
            O => \N__48219\,
            I => \N__48213\
        );

    \I__9917\ : Span4Mux_v
    port map (
            O => \N__48216\,
            I => \N__48210\
        );

    \I__9916\ : InMux
    port map (
            O => \N__48213\,
            I => \N__48207\
        );

    \I__9915\ : Odrv4
    port map (
            O => \N__48210\,
            I => \c0.n19_adj_3336\
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__48207\,
            I => \c0.n19_adj_3336\
        );

    \I__9913\ : CascadeMux
    port map (
            O => \N__48202\,
            I => \c0.n39_adj_3334_cascade_\
        );

    \I__9912\ : InMux
    port map (
            O => \N__48199\,
            I => \N__48196\
        );

    \I__9911\ : LocalMux
    port map (
            O => \N__48196\,
            I => \c0.n25_adj_3431\
        );

    \I__9910\ : InMux
    port map (
            O => \N__48193\,
            I => \N__48187\
        );

    \I__9909\ : InMux
    port map (
            O => \N__48192\,
            I => \N__48187\
        );

    \I__9908\ : LocalMux
    port map (
            O => \N__48187\,
            I => \N__48184\
        );

    \I__9907\ : Odrv12
    port map (
            O => \N__48184\,
            I => \c0.n42_adj_3367\
        );

    \I__9906\ : InMux
    port map (
            O => \N__48181\,
            I => \N__48178\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__48178\,
            I => \N__48174\
        );

    \I__9904\ : InMux
    port map (
            O => \N__48177\,
            I => \N__48171\
        );

    \I__9903\ : Span4Mux_v
    port map (
            O => \N__48174\,
            I => \N__48168\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__48171\,
            I => \c0.n43_adj_3386\
        );

    \I__9901\ : Odrv4
    port map (
            O => \N__48168\,
            I => \c0.n43_adj_3386\
        );

    \I__9900\ : InMux
    port map (
            O => \N__48163\,
            I => \N__48157\
        );

    \I__9899\ : InMux
    port map (
            O => \N__48162\,
            I => \N__48157\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__48157\,
            I => \N__48154\
        );

    \I__9897\ : Span4Mux_v
    port map (
            O => \N__48154\,
            I => \N__48151\
        );

    \I__9896\ : Span4Mux_h
    port map (
            O => \N__48151\,
            I => \N__48148\
        );

    \I__9895\ : Odrv4
    port map (
            O => \N__48148\,
            I => \c0.n40_adj_3366\
        );

    \I__9894\ : InMux
    port map (
            O => \N__48145\,
            I => \N__48142\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__48142\,
            I => \c0.n30_adj_3429\
        );

    \I__9892\ : InMux
    port map (
            O => \N__48139\,
            I => \N__48136\
        );

    \I__9891\ : LocalMux
    port map (
            O => \N__48136\,
            I => \c0.n46\
        );

    \I__9890\ : InMux
    port map (
            O => \N__48133\,
            I => \N__48127\
        );

    \I__9889\ : InMux
    port map (
            O => \N__48132\,
            I => \N__48120\
        );

    \I__9888\ : InMux
    port map (
            O => \N__48131\,
            I => \N__48120\
        );

    \I__9887\ : InMux
    port map (
            O => \N__48130\,
            I => \N__48120\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__48127\,
            I => \N__48117\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__48120\,
            I => \N__48114\
        );

    \I__9884\ : Span4Mux_v
    port map (
            O => \N__48117\,
            I => \N__48111\
        );

    \I__9883\ : Span4Mux_h
    port map (
            O => \N__48114\,
            I => \N__48108\
        );

    \I__9882\ : Odrv4
    port map (
            O => \N__48111\,
            I => \c0.n8\
        );

    \I__9881\ : Odrv4
    port map (
            O => \N__48108\,
            I => \c0.n8\
        );

    \I__9880\ : InMux
    port map (
            O => \N__48103\,
            I => \N__48099\
        );

    \I__9879\ : CascadeMux
    port map (
            O => \N__48102\,
            I => \N__48096\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__48099\,
            I => \N__48093\
        );

    \I__9877\ : InMux
    port map (
            O => \N__48096\,
            I => \N__48090\
        );

    \I__9876\ : Odrv12
    port map (
            O => \N__48093\,
            I => \c0.n84\
        );

    \I__9875\ : LocalMux
    port map (
            O => \N__48090\,
            I => \c0.n84\
        );

    \I__9874\ : CascadeMux
    port map (
            O => \N__48085\,
            I => \c0.n19824_cascade_\
        );

    \I__9873\ : InMux
    port map (
            O => \N__48082\,
            I => \N__48078\
        );

    \I__9872\ : InMux
    port map (
            O => \N__48081\,
            I => \N__48075\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__48078\,
            I => \N__48072\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__48075\,
            I => \N__48069\
        );

    \I__9869\ : Span4Mux_h
    port map (
            O => \N__48072\,
            I => \N__48065\
        );

    \I__9868\ : Span4Mux_v
    port map (
            O => \N__48069\,
            I => \N__48062\
        );

    \I__9867\ : InMux
    port map (
            O => \N__48068\,
            I => \N__48059\
        );

    \I__9866\ : Odrv4
    port map (
            O => \N__48065\,
            I => \c0.n29\
        );

    \I__9865\ : Odrv4
    port map (
            O => \N__48062\,
            I => \c0.n29\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__48059\,
            I => \c0.n29\
        );

    \I__9863\ : CascadeMux
    port map (
            O => \N__48052\,
            I => \c0.n18_adj_3360_cascade_\
        );

    \I__9862\ : CascadeMux
    port map (
            O => \N__48049\,
            I => \c0.n32_adj_3362_cascade_\
        );

    \I__9861\ : CascadeMux
    port map (
            O => \N__48046\,
            I => \c0.n20112_cascade_\
        );

    \I__9860\ : CascadeMux
    port map (
            O => \N__48043\,
            I => \c0.n12_adj_3249_cascade_\
        );

    \I__9859\ : InMux
    port map (
            O => \N__48040\,
            I => \N__48037\
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__48037\,
            I => \c0.n12056\
        );

    \I__9857\ : InMux
    port map (
            O => \N__48034\,
            I => \N__48027\
        );

    \I__9856\ : InMux
    port map (
            O => \N__48033\,
            I => \N__48027\
        );

    \I__9855\ : CascadeMux
    port map (
            O => \N__48032\,
            I => \N__48024\
        );

    \I__9854\ : LocalMux
    port map (
            O => \N__48027\,
            I => \N__48021\
        );

    \I__9853\ : InMux
    port map (
            O => \N__48024\,
            I => \N__48018\
        );

    \I__9852\ : Sp12to4
    port map (
            O => \N__48021\,
            I => \N__48015\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__48018\,
            I => \N__48012\
        );

    \I__9850\ : Odrv12
    port map (
            O => \N__48015\,
            I => \c0.n19301\
        );

    \I__9849\ : Odrv12
    port map (
            O => \N__48012\,
            I => \c0.n19301\
        );

    \I__9848\ : CascadeMux
    port map (
            O => \N__48007\,
            I => \c0.n19301_cascade_\
        );

    \I__9847\ : CascadeMux
    port map (
            O => \N__48004\,
            I => \c0.n31_adj_3126_cascade_\
        );

    \I__9846\ : CascadeMux
    port map (
            O => \N__48001\,
            I => \N__47997\
        );

    \I__9845\ : CascadeMux
    port map (
            O => \N__48000\,
            I => \N__47994\
        );

    \I__9844\ : InMux
    port map (
            O => \N__47997\,
            I => \N__47989\
        );

    \I__9843\ : InMux
    port map (
            O => \N__47994\,
            I => \N__47989\
        );

    \I__9842\ : LocalMux
    port map (
            O => \N__47989\,
            I => \N__47986\
        );

    \I__9841\ : Span4Mux_h
    port map (
            O => \N__47986\,
            I => \N__47983\
        );

    \I__9840\ : Odrv4
    port map (
            O => \N__47983\,
            I => \c0.n19427\
        );

    \I__9839\ : InMux
    port map (
            O => \N__47980\,
            I => \N__47977\
        );

    \I__9838\ : LocalMux
    port map (
            O => \N__47977\,
            I => \N__47972\
        );

    \I__9837\ : InMux
    port map (
            O => \N__47976\,
            I => \N__47967\
        );

    \I__9836\ : InMux
    port map (
            O => \N__47975\,
            I => \N__47967\
        );

    \I__9835\ : Span4Mux_h
    port map (
            O => \N__47972\,
            I => \N__47964\
        );

    \I__9834\ : LocalMux
    port map (
            O => \N__47967\,
            I => \N__47961\
        );

    \I__9833\ : Odrv4
    port map (
            O => \N__47964\,
            I => \c0.n19551\
        );

    \I__9832\ : Odrv12
    port map (
            O => \N__47961\,
            I => \c0.n19551\
        );

    \I__9831\ : InMux
    port map (
            O => \N__47956\,
            I => \N__47953\
        );

    \I__9830\ : LocalMux
    port map (
            O => \N__47953\,
            I => \N__47950\
        );

    \I__9829\ : Span4Mux_h
    port map (
            O => \N__47950\,
            I => \N__47947\
        );

    \I__9828\ : Odrv4
    port map (
            O => \N__47947\,
            I => \c0.n27_adj_3455\
        );

    \I__9827\ : CascadeMux
    port map (
            O => \N__47944\,
            I => \c0.n46_cascade_\
        );

    \I__9826\ : InMux
    port map (
            O => \N__47941\,
            I => \N__47938\
        );

    \I__9825\ : LocalMux
    port map (
            O => \N__47938\,
            I => \N__47935\
        );

    \I__9824\ : Span4Mux_h
    port map (
            O => \N__47935\,
            I => \N__47932\
        );

    \I__9823\ : Span4Mux_v
    port map (
            O => \N__47932\,
            I => \N__47929\
        );

    \I__9822\ : Odrv4
    port map (
            O => \N__47929\,
            I => \c0.n31_adj_3532\
        );

    \I__9821\ : InMux
    port map (
            O => \N__47926\,
            I => \N__47922\
        );

    \I__9820\ : InMux
    port map (
            O => \N__47925\,
            I => \N__47918\
        );

    \I__9819\ : LocalMux
    port map (
            O => \N__47922\,
            I => \N__47915\
        );

    \I__9818\ : InMux
    port map (
            O => \N__47921\,
            I => \N__47912\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__47918\,
            I => \N__47908\
        );

    \I__9816\ : Span4Mux_v
    port map (
            O => \N__47915\,
            I => \N__47903\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__47912\,
            I => \N__47903\
        );

    \I__9814\ : InMux
    port map (
            O => \N__47911\,
            I => \N__47900\
        );

    \I__9813\ : Span4Mux_v
    port map (
            O => \N__47908\,
            I => \N__47897\
        );

    \I__9812\ : Span4Mux_h
    port map (
            O => \N__47903\,
            I => \N__47894\
        );

    \I__9811\ : LocalMux
    port map (
            O => \N__47900\,
            I => \c0.n11537\
        );

    \I__9810\ : Odrv4
    port map (
            O => \N__47897\,
            I => \c0.n11537\
        );

    \I__9809\ : Odrv4
    port map (
            O => \N__47894\,
            I => \c0.n11537\
        );

    \I__9808\ : InMux
    port map (
            O => \N__47887\,
            I => \N__47882\
        );

    \I__9807\ : CascadeMux
    port map (
            O => \N__47886\,
            I => \N__47879\
        );

    \I__9806\ : InMux
    port map (
            O => \N__47885\,
            I => \N__47876\
        );

    \I__9805\ : LocalMux
    port map (
            O => \N__47882\,
            I => \N__47873\
        );

    \I__9804\ : InMux
    port map (
            O => \N__47879\,
            I => \N__47870\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__47876\,
            I => \N__47867\
        );

    \I__9802\ : Span12Mux_h
    port map (
            O => \N__47873\,
            I => \N__47864\
        );

    \I__9801\ : LocalMux
    port map (
            O => \N__47870\,
            I => \c0.data_in_frame_15_6\
        );

    \I__9800\ : Odrv4
    port map (
            O => \N__47867\,
            I => \c0.data_in_frame_15_6\
        );

    \I__9799\ : Odrv12
    port map (
            O => \N__47864\,
            I => \c0.data_in_frame_15_6\
        );

    \I__9798\ : CascadeMux
    port map (
            O => \N__47857\,
            I => \c0.n16_adj_3481_cascade_\
        );

    \I__9797\ : CascadeMux
    port map (
            O => \N__47854\,
            I => \c0.n11815_cascade_\
        );

    \I__9796\ : InMux
    port map (
            O => \N__47851\,
            I => \N__47845\
        );

    \I__9795\ : InMux
    port map (
            O => \N__47850\,
            I => \N__47845\
        );

    \I__9794\ : LocalMux
    port map (
            O => \N__47845\,
            I => \N__47842\
        );

    \I__9793\ : Span12Mux_v
    port map (
            O => \N__47842\,
            I => \N__47839\
        );

    \I__9792\ : Odrv12
    port map (
            O => \N__47839\,
            I => \c0.n19291\
        );

    \I__9791\ : CascadeMux
    port map (
            O => \N__47836\,
            I => \N__47831\
        );

    \I__9790\ : InMux
    port map (
            O => \N__47835\,
            I => \N__47827\
        );

    \I__9789\ : InMux
    port map (
            O => \N__47834\,
            I => \N__47824\
        );

    \I__9788\ : InMux
    port map (
            O => \N__47831\,
            I => \N__47821\
        );

    \I__9787\ : InMux
    port map (
            O => \N__47830\,
            I => \N__47818\
        );

    \I__9786\ : LocalMux
    port map (
            O => \N__47827\,
            I => \N__47815\
        );

    \I__9785\ : LocalMux
    port map (
            O => \N__47824\,
            I => \N__47812\
        );

    \I__9784\ : LocalMux
    port map (
            O => \N__47821\,
            I => \N__47809\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__47818\,
            I => \N__47804\
        );

    \I__9782\ : Span4Mux_h
    port map (
            O => \N__47815\,
            I => \N__47804\
        );

    \I__9781\ : Span4Mux_v
    port map (
            O => \N__47812\,
            I => \N__47799\
        );

    \I__9780\ : Span4Mux_v
    port map (
            O => \N__47809\,
            I => \N__47794\
        );

    \I__9779\ : Span4Mux_v
    port map (
            O => \N__47804\,
            I => \N__47794\
        );

    \I__9778\ : InMux
    port map (
            O => \N__47803\,
            I => \N__47789\
        );

    \I__9777\ : InMux
    port map (
            O => \N__47802\,
            I => \N__47789\
        );

    \I__9776\ : Odrv4
    port map (
            O => \N__47799\,
            I => data_in_frame_16_1
        );

    \I__9775\ : Odrv4
    port map (
            O => \N__47794\,
            I => data_in_frame_16_1
        );

    \I__9774\ : LocalMux
    port map (
            O => \N__47789\,
            I => data_in_frame_16_1
        );

    \I__9773\ : CascadeMux
    port map (
            O => \N__47782\,
            I => \c0.n12056_cascade_\
        );

    \I__9772\ : InMux
    port map (
            O => \N__47779\,
            I => \N__47776\
        );

    \I__9771\ : LocalMux
    port map (
            O => \N__47776\,
            I => \c0.n12_adj_3249\
        );

    \I__9770\ : InMux
    port map (
            O => \N__47773\,
            I => \N__47769\
        );

    \I__9769\ : InMux
    port map (
            O => \N__47772\,
            I => \N__47764\
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__47769\,
            I => \N__47761\
        );

    \I__9767\ : InMux
    port map (
            O => \N__47768\,
            I => \N__47758\
        );

    \I__9766\ : CascadeMux
    port map (
            O => \N__47767\,
            I => \N__47755\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__47764\,
            I => \N__47752\
        );

    \I__9764\ : Span4Mux_v
    port map (
            O => \N__47761\,
            I => \N__47749\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__47758\,
            I => \N__47746\
        );

    \I__9762\ : InMux
    port map (
            O => \N__47755\,
            I => \N__47742\
        );

    \I__9761\ : Span4Mux_v
    port map (
            O => \N__47752\,
            I => \N__47739\
        );

    \I__9760\ : Span4Mux_h
    port map (
            O => \N__47749\,
            I => \N__47734\
        );

    \I__9759\ : Span4Mux_v
    port map (
            O => \N__47746\,
            I => \N__47734\
        );

    \I__9758\ : InMux
    port map (
            O => \N__47745\,
            I => \N__47731\
        );

    \I__9757\ : LocalMux
    port map (
            O => \N__47742\,
            I => \c0.data_in_frame_12_2\
        );

    \I__9756\ : Odrv4
    port map (
            O => \N__47739\,
            I => \c0.data_in_frame_12_2\
        );

    \I__9755\ : Odrv4
    port map (
            O => \N__47734\,
            I => \c0.data_in_frame_12_2\
        );

    \I__9754\ : LocalMux
    port map (
            O => \N__47731\,
            I => \c0.data_in_frame_12_2\
        );

    \I__9753\ : InMux
    port map (
            O => \N__47722\,
            I => \N__47719\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__47719\,
            I => \N__47716\
        );

    \I__9751\ : Span4Mux_v
    port map (
            O => \N__47716\,
            I => \N__47712\
        );

    \I__9750\ : InMux
    port map (
            O => \N__47715\,
            I => \N__47709\
        );

    \I__9749\ : Odrv4
    port map (
            O => \N__47712\,
            I => \c0.n7_adj_3491\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__47709\,
            I => \c0.n7_adj_3491\
        );

    \I__9747\ : InMux
    port map (
            O => \N__47704\,
            I => \N__47701\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__47701\,
            I => \N__47698\
        );

    \I__9745\ : Span4Mux_v
    port map (
            O => \N__47698\,
            I => \N__47695\
        );

    \I__9744\ : Odrv4
    port map (
            O => \N__47695\,
            I => \c0.n30_adj_3531\
        );

    \I__9743\ : InMux
    port map (
            O => \N__47692\,
            I => \N__47689\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__47689\,
            I => \N__47685\
        );

    \I__9741\ : InMux
    port map (
            O => \N__47688\,
            I => \N__47681\
        );

    \I__9740\ : Span4Mux_v
    port map (
            O => \N__47685\,
            I => \N__47678\
        );

    \I__9739\ : InMux
    port map (
            O => \N__47684\,
            I => \N__47675\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__47681\,
            I => \N__47670\
        );

    \I__9737\ : Span4Mux_h
    port map (
            O => \N__47678\,
            I => \N__47670\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__47675\,
            I => \N__47667\
        );

    \I__9735\ : Span4Mux_v
    port map (
            O => \N__47670\,
            I => \N__47664\
        );

    \I__9734\ : Span4Mux_v
    port map (
            O => \N__47667\,
            I => \N__47661\
        );

    \I__9733\ : Odrv4
    port map (
            O => \N__47664\,
            I => \c0.n12_adj_3034\
        );

    \I__9732\ : Odrv4
    port map (
            O => \N__47661\,
            I => \c0.n12_adj_3034\
        );

    \I__9731\ : CascadeMux
    port map (
            O => \N__47656\,
            I => \c0.n32_adj_3077_cascade_\
        );

    \I__9730\ : CascadeMux
    port map (
            O => \N__47653\,
            I => \N__47650\
        );

    \I__9729\ : InMux
    port map (
            O => \N__47650\,
            I => \N__47647\
        );

    \I__9728\ : LocalMux
    port map (
            O => \N__47647\,
            I => \N__47643\
        );

    \I__9727\ : InMux
    port map (
            O => \N__47646\,
            I => \N__47640\
        );

    \I__9726\ : Span4Mux_h
    port map (
            O => \N__47643\,
            I => \N__47635\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__47640\,
            I => \N__47635\
        );

    \I__9724\ : Odrv4
    port map (
            O => \N__47635\,
            I => \c0.n19372\
        );

    \I__9723\ : CascadeMux
    port map (
            O => \N__47632\,
            I => \c0.n21047_cascade_\
        );

    \I__9722\ : InMux
    port map (
            O => \N__47629\,
            I => \N__47626\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__47626\,
            I => \N__47623\
        );

    \I__9720\ : Odrv4
    port map (
            O => \N__47623\,
            I => \c0.n42_adj_3111\
        );

    \I__9719\ : InMux
    port map (
            O => \N__47620\,
            I => \N__47616\
        );

    \I__9718\ : CascadeMux
    port map (
            O => \N__47619\,
            I => \N__47611\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__47616\,
            I => \N__47608\
        );

    \I__9716\ : InMux
    port map (
            O => \N__47615\,
            I => \N__47605\
        );

    \I__9715\ : InMux
    port map (
            O => \N__47614\,
            I => \N__47602\
        );

    \I__9714\ : InMux
    port map (
            O => \N__47611\,
            I => \N__47599\
        );

    \I__9713\ : Span4Mux_v
    port map (
            O => \N__47608\,
            I => \N__47593\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__47605\,
            I => \N__47588\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__47602\,
            I => \N__47588\
        );

    \I__9710\ : LocalMux
    port map (
            O => \N__47599\,
            I => \N__47585\
        );

    \I__9709\ : InMux
    port map (
            O => \N__47598\,
            I => \N__47582\
        );

    \I__9708\ : InMux
    port map (
            O => \N__47597\,
            I => \N__47577\
        );

    \I__9707\ : InMux
    port map (
            O => \N__47596\,
            I => \N__47577\
        );

    \I__9706\ : Span4Mux_h
    port map (
            O => \N__47593\,
            I => \N__47572\
        );

    \I__9705\ : Span4Mux_v
    port map (
            O => \N__47588\,
            I => \N__47572\
        );

    \I__9704\ : Span4Mux_v
    port map (
            O => \N__47585\,
            I => \N__47569\
        );

    \I__9703\ : LocalMux
    port map (
            O => \N__47582\,
            I => \c0.data_in_frame_3_0\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__47577\,
            I => \c0.data_in_frame_3_0\
        );

    \I__9701\ : Odrv4
    port map (
            O => \N__47572\,
            I => \c0.data_in_frame_3_0\
        );

    \I__9700\ : Odrv4
    port map (
            O => \N__47569\,
            I => \c0.data_in_frame_3_0\
        );

    \I__9699\ : InMux
    port map (
            O => \N__47560\,
            I => \N__47556\
        );

    \I__9698\ : CascadeMux
    port map (
            O => \N__47559\,
            I => \N__47552\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__47556\,
            I => \N__47549\
        );

    \I__9696\ : InMux
    port map (
            O => \N__47555\,
            I => \N__47542\
        );

    \I__9695\ : InMux
    port map (
            O => \N__47552\,
            I => \N__47539\
        );

    \I__9694\ : Span4Mux_h
    port map (
            O => \N__47549\,
            I => \N__47536\
        );

    \I__9693\ : InMux
    port map (
            O => \N__47548\,
            I => \N__47531\
        );

    \I__9692\ : InMux
    port map (
            O => \N__47547\,
            I => \N__47531\
        );

    \I__9691\ : InMux
    port map (
            O => \N__47546\,
            I => \N__47526\
        );

    \I__9690\ : InMux
    port map (
            O => \N__47545\,
            I => \N__47526\
        );

    \I__9689\ : LocalMux
    port map (
            O => \N__47542\,
            I => \N__47521\
        );

    \I__9688\ : LocalMux
    port map (
            O => \N__47539\,
            I => \N__47521\
        );

    \I__9687\ : Odrv4
    port map (
            O => \N__47536\,
            I => \c0.data_in_frame_2_6\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__47531\,
            I => \c0.data_in_frame_2_6\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__47526\,
            I => \c0.data_in_frame_2_6\
        );

    \I__9684\ : Odrv12
    port map (
            O => \N__47521\,
            I => \c0.data_in_frame_2_6\
        );

    \I__9683\ : CascadeMux
    port map (
            O => \N__47512\,
            I => \c0.n10_adj_3014_cascade_\
        );

    \I__9682\ : InMux
    port map (
            O => \N__47509\,
            I => \N__47505\
        );

    \I__9681\ : CascadeMux
    port map (
            O => \N__47508\,
            I => \N__47502\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__47505\,
            I => \N__47499\
        );

    \I__9679\ : InMux
    port map (
            O => \N__47502\,
            I => \N__47496\
        );

    \I__9678\ : Span4Mux_h
    port map (
            O => \N__47499\,
            I => \N__47491\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__47496\,
            I => \N__47491\
        );

    \I__9676\ : Span4Mux_v
    port map (
            O => \N__47491\,
            I => \N__47487\
        );

    \I__9675\ : InMux
    port map (
            O => \N__47490\,
            I => \N__47484\
        );

    \I__9674\ : Odrv4
    port map (
            O => \N__47487\,
            I => \c0.n40\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__47484\,
            I => \c0.n40\
        );

    \I__9672\ : CascadeMux
    port map (
            O => \N__47479\,
            I => \c0.n16_adj_3218_cascade_\
        );

    \I__9671\ : InMux
    port map (
            O => \N__47476\,
            I => \N__47473\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__47473\,
            I => \c0.n10_adj_3538\
        );

    \I__9669\ : InMux
    port map (
            O => \N__47470\,
            I => \N__47467\
        );

    \I__9668\ : LocalMux
    port map (
            O => \N__47467\,
            I => \N__47464\
        );

    \I__9667\ : Odrv12
    port map (
            O => \N__47464\,
            I => \c0.n85\
        );

    \I__9666\ : InMux
    port map (
            O => \N__47461\,
            I => \N__47458\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__47458\,
            I => \N__47455\
        );

    \I__9664\ : Span4Mux_h
    port map (
            O => \N__47455\,
            I => \N__47451\
        );

    \I__9663\ : InMux
    port map (
            O => \N__47454\,
            I => \N__47448\
        );

    \I__9662\ : Odrv4
    port map (
            O => \N__47451\,
            I => \c0.n37\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__47448\,
            I => \c0.n37\
        );

    \I__9660\ : CascadeMux
    port map (
            O => \N__47443\,
            I => \c0.n67_cascade_\
        );

    \I__9659\ : InMux
    port map (
            O => \N__47440\,
            I => \N__47437\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__47437\,
            I => \c0.n96\
        );

    \I__9657\ : InMux
    port map (
            O => \N__47434\,
            I => \N__47431\
        );

    \I__9656\ : LocalMux
    port map (
            O => \N__47431\,
            I => \c0.n83\
        );

    \I__9655\ : InMux
    port map (
            O => \N__47428\,
            I => \N__47425\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__47425\,
            I => \N__47421\
        );

    \I__9653\ : InMux
    port map (
            O => \N__47424\,
            I => \N__47418\
        );

    \I__9652\ : Span4Mux_v
    port map (
            O => \N__47421\,
            I => \N__47413\
        );

    \I__9651\ : LocalMux
    port map (
            O => \N__47418\,
            I => \N__47413\
        );

    \I__9650\ : Span4Mux_h
    port map (
            O => \N__47413\,
            I => \N__47410\
        );

    \I__9649\ : Odrv4
    port map (
            O => \N__47410\,
            I => \c0.n40_adj_3032\
        );

    \I__9648\ : CascadeMux
    port map (
            O => \N__47407\,
            I => \c0.n100_cascade_\
        );

    \I__9647\ : CascadeMux
    port map (
            O => \N__47404\,
            I => \N__47401\
        );

    \I__9646\ : InMux
    port map (
            O => \N__47401\,
            I => \N__47398\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__47398\,
            I => \c0.n102\
        );

    \I__9644\ : InMux
    port map (
            O => \N__47395\,
            I => \N__47392\
        );

    \I__9643\ : LocalMux
    port map (
            O => \N__47392\,
            I => \N__47388\
        );

    \I__9642\ : InMux
    port map (
            O => \N__47391\,
            I => \N__47385\
        );

    \I__9641\ : Span4Mux_h
    port map (
            O => \N__47388\,
            I => \N__47382\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__47385\,
            I => \N__47379\
        );

    \I__9639\ : Odrv4
    port map (
            O => \N__47382\,
            I => \c0.n4_adj_3009\
        );

    \I__9638\ : Odrv12
    port map (
            O => \N__47379\,
            I => \c0.n4_adj_3009\
        );

    \I__9637\ : InMux
    port map (
            O => \N__47374\,
            I => \N__47371\
        );

    \I__9636\ : LocalMux
    port map (
            O => \N__47371\,
            I => \N__47366\
        );

    \I__9635\ : InMux
    port map (
            O => \N__47370\,
            I => \N__47361\
        );

    \I__9634\ : InMux
    port map (
            O => \N__47369\,
            I => \N__47361\
        );

    \I__9633\ : Odrv4
    port map (
            O => \N__47366\,
            I => \c0.n21_adj_3010\
        );

    \I__9632\ : LocalMux
    port map (
            O => \N__47361\,
            I => \c0.n21_adj_3010\
        );

    \I__9631\ : InMux
    port map (
            O => \N__47356\,
            I => \N__47353\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__47353\,
            I => \c0.n28_adj_3023\
        );

    \I__9629\ : InMux
    port map (
            O => \N__47350\,
            I => \N__47347\
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__47347\,
            I => \c0.n17_adj_3508\
        );

    \I__9627\ : CascadeMux
    port map (
            O => \N__47344\,
            I => \N__47341\
        );

    \I__9626\ : InMux
    port map (
            O => \N__47341\,
            I => \N__47337\
        );

    \I__9625\ : InMux
    port map (
            O => \N__47340\,
            I => \N__47333\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__47337\,
            I => \N__47330\
        );

    \I__9623\ : InMux
    port map (
            O => \N__47336\,
            I => \N__47327\
        );

    \I__9622\ : LocalMux
    port map (
            O => \N__47333\,
            I => \N__47322\
        );

    \I__9621\ : Span4Mux_h
    port map (
            O => \N__47330\,
            I => \N__47322\
        );

    \I__9620\ : LocalMux
    port map (
            O => \N__47327\,
            I => \c0.n19966\
        );

    \I__9619\ : Odrv4
    port map (
            O => \N__47322\,
            I => \c0.n19966\
        );

    \I__9618\ : InMux
    port map (
            O => \N__47317\,
            I => \N__47314\
        );

    \I__9617\ : LocalMux
    port map (
            O => \N__47314\,
            I => \c0.n30_adj_3075\
        );

    \I__9616\ : InMux
    port map (
            O => \N__47311\,
            I => \N__47308\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__47308\,
            I => \N__47305\
        );

    \I__9614\ : Span4Mux_v
    port map (
            O => \N__47305\,
            I => \N__47302\
        );

    \I__9613\ : Odrv4
    port map (
            O => \N__47302\,
            I => \c0.n21277\
        );

    \I__9612\ : InMux
    port map (
            O => \N__47299\,
            I => \N__47289\
        );

    \I__9611\ : InMux
    port map (
            O => \N__47298\,
            I => \N__47289\
        );

    \I__9610\ : InMux
    port map (
            O => \N__47297\,
            I => \N__47289\
        );

    \I__9609\ : InMux
    port map (
            O => \N__47296\,
            I => \N__47286\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__47289\,
            I => \c0.n4_adj_3406\
        );

    \I__9607\ : LocalMux
    port map (
            O => \N__47286\,
            I => \c0.n4_adj_3406\
        );

    \I__9606\ : CascadeMux
    port map (
            O => \N__47281\,
            I => \c0.n14_adj_3476_cascade_\
        );

    \I__9605\ : CascadeMux
    port map (
            O => \N__47278\,
            I => \N__47275\
        );

    \I__9604\ : InMux
    port map (
            O => \N__47275\,
            I => \N__47271\
        );

    \I__9603\ : InMux
    port map (
            O => \N__47274\,
            I => \N__47266\
        );

    \I__9602\ : LocalMux
    port map (
            O => \N__47271\,
            I => \N__47263\
        );

    \I__9601\ : InMux
    port map (
            O => \N__47270\,
            I => \N__47260\
        );

    \I__9600\ : CascadeMux
    port map (
            O => \N__47269\,
            I => \N__47256\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__47266\,
            I => \N__47252\
        );

    \I__9598\ : Span4Mux_v
    port map (
            O => \N__47263\,
            I => \N__47247\
        );

    \I__9597\ : LocalMux
    port map (
            O => \N__47260\,
            I => \N__47247\
        );

    \I__9596\ : InMux
    port map (
            O => \N__47259\,
            I => \N__47244\
        );

    \I__9595\ : InMux
    port map (
            O => \N__47256\,
            I => \N__47239\
        );

    \I__9594\ : InMux
    port map (
            O => \N__47255\,
            I => \N__47239\
        );

    \I__9593\ : Span4Mux_v
    port map (
            O => \N__47252\,
            I => \N__47236\
        );

    \I__9592\ : Odrv4
    port map (
            O => \N__47247\,
            I => \c0.data_in_frame_7_3\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__47244\,
            I => \c0.data_in_frame_7_3\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__47239\,
            I => \c0.data_in_frame_7_3\
        );

    \I__9589\ : Odrv4
    port map (
            O => \N__47236\,
            I => \c0.data_in_frame_7_3\
        );

    \I__9588\ : InMux
    port map (
            O => \N__47227\,
            I => \N__47224\
        );

    \I__9587\ : LocalMux
    port map (
            O => \N__47224\,
            I => \c0.n19508\
        );

    \I__9586\ : InMux
    port map (
            O => \N__47221\,
            I => \N__47218\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__47218\,
            I => \N__47213\
        );

    \I__9584\ : InMux
    port map (
            O => \N__47217\,
            I => \N__47210\
        );

    \I__9583\ : CascadeMux
    port map (
            O => \N__47216\,
            I => \N__47207\
        );

    \I__9582\ : Span4Mux_h
    port map (
            O => \N__47213\,
            I => \N__47200\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__47210\,
            I => \N__47200\
        );

    \I__9580\ : InMux
    port map (
            O => \N__47207\,
            I => \N__47197\
        );

    \I__9579\ : InMux
    port map (
            O => \N__47206\,
            I => \N__47192\
        );

    \I__9578\ : InMux
    port map (
            O => \N__47205\,
            I => \N__47192\
        );

    \I__9577\ : Span4Mux_v
    port map (
            O => \N__47200\,
            I => \N__47189\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__47197\,
            I => \c0.data_in_frame_2_0\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__47192\,
            I => \c0.data_in_frame_2_0\
        );

    \I__9574\ : Odrv4
    port map (
            O => \N__47189\,
            I => \c0.data_in_frame_2_0\
        );

    \I__9573\ : CascadeMux
    port map (
            O => \N__47182\,
            I => \N__47179\
        );

    \I__9572\ : InMux
    port map (
            O => \N__47179\,
            I => \N__47176\
        );

    \I__9571\ : LocalMux
    port map (
            O => \N__47176\,
            I => \c0.n8_adj_3397\
        );

    \I__9570\ : CascadeMux
    port map (
            O => \N__47173\,
            I => \c0.n11833_cascade_\
        );

    \I__9569\ : CascadeMux
    port map (
            O => \N__47170\,
            I => \c0.n92_cascade_\
        );

    \I__9568\ : InMux
    port map (
            O => \N__47167\,
            I => \N__47164\
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__47164\,
            I => \c0.n80\
        );

    \I__9566\ : InMux
    port map (
            O => \N__47161\,
            I => \N__47158\
        );

    \I__9565\ : LocalMux
    port map (
            O => \N__47158\,
            I => \c0.n19196\
        );

    \I__9564\ : CascadeMux
    port map (
            O => \N__47155\,
            I => \N__47149\
        );

    \I__9563\ : CascadeMux
    port map (
            O => \N__47154\,
            I => \N__47146\
        );

    \I__9562\ : CascadeMux
    port map (
            O => \N__47153\,
            I => \N__47142\
        );

    \I__9561\ : CascadeMux
    port map (
            O => \N__47152\,
            I => \N__47139\
        );

    \I__9560\ : InMux
    port map (
            O => \N__47149\,
            I => \N__47136\
        );

    \I__9559\ : InMux
    port map (
            O => \N__47146\,
            I => \N__47131\
        );

    \I__9558\ : InMux
    port map (
            O => \N__47145\,
            I => \N__47131\
        );

    \I__9557\ : InMux
    port map (
            O => \N__47142\,
            I => \N__47128\
        );

    \I__9556\ : InMux
    port map (
            O => \N__47139\,
            I => \N__47125\
        );

    \I__9555\ : LocalMux
    port map (
            O => \N__47136\,
            I => \c0.data_in_frame_4_5\
        );

    \I__9554\ : LocalMux
    port map (
            O => \N__47131\,
            I => \c0.data_in_frame_4_5\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__47128\,
            I => \c0.data_in_frame_4_5\
        );

    \I__9552\ : LocalMux
    port map (
            O => \N__47125\,
            I => \c0.data_in_frame_4_5\
        );

    \I__9551\ : InMux
    port map (
            O => \N__47116\,
            I => \N__47113\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__47113\,
            I => \c0.n54\
        );

    \I__9549\ : InMux
    port map (
            O => \N__47110\,
            I => \N__47107\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__47107\,
            I => \c0.n90\
        );

    \I__9547\ : InMux
    port map (
            O => \N__47104\,
            I => \N__47101\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__47101\,
            I => \c0.n98\
        );

    \I__9545\ : InMux
    port map (
            O => \N__47098\,
            I => \N__47095\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__47095\,
            I => \N__47092\
        );

    \I__9543\ : Span4Mux_v
    port map (
            O => \N__47092\,
            I => \N__47089\
        );

    \I__9542\ : Odrv4
    port map (
            O => \N__47089\,
            I => \c0.n12085\
        );

    \I__9541\ : InMux
    port map (
            O => \N__47086\,
            I => \N__47083\
        );

    \I__9540\ : LocalMux
    port map (
            O => \N__47083\,
            I => \N__47079\
        );

    \I__9539\ : InMux
    port map (
            O => \N__47082\,
            I => \N__47076\
        );

    \I__9538\ : Odrv4
    port map (
            O => \N__47079\,
            I => \c0.n11865\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__47076\,
            I => \c0.n11865\
        );

    \I__9536\ : CascadeMux
    port map (
            O => \N__47071\,
            I => \c0.n12085_cascade_\
        );

    \I__9535\ : CascadeMux
    port map (
            O => \N__47068\,
            I => \N__47065\
        );

    \I__9534\ : InMux
    port map (
            O => \N__47065\,
            I => \N__47062\
        );

    \I__9533\ : LocalMux
    port map (
            O => \N__47062\,
            I => \N__47059\
        );

    \I__9532\ : Span4Mux_h
    port map (
            O => \N__47059\,
            I => \N__47056\
        );

    \I__9531\ : Span4Mux_v
    port map (
            O => \N__47056\,
            I => \N__47053\
        );

    \I__9530\ : Span4Mux_h
    port map (
            O => \N__47053\,
            I => \N__47049\
        );

    \I__9529\ : InMux
    port map (
            O => \N__47052\,
            I => \N__47046\
        );

    \I__9528\ : Odrv4
    port map (
            O => \N__47049\,
            I => \c0.n6495\
        );

    \I__9527\ : LocalMux
    port map (
            O => \N__47046\,
            I => \c0.n6495\
        );

    \I__9526\ : InMux
    port map (
            O => \N__47041\,
            I => \N__47038\
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__47038\,
            I => \N__47035\
        );

    \I__9524\ : Span4Mux_h
    port map (
            O => \N__47035\,
            I => \N__47029\
        );

    \I__9523\ : InMux
    port map (
            O => \N__47034\,
            I => \N__47026\
        );

    \I__9522\ : InMux
    port map (
            O => \N__47033\,
            I => \N__47021\
        );

    \I__9521\ : InMux
    port map (
            O => \N__47032\,
            I => \N__47021\
        );

    \I__9520\ : Odrv4
    port map (
            O => \N__47029\,
            I => data_in_2_4
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__47026\,
            I => data_in_2_4
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__47021\,
            I => data_in_2_4
        );

    \I__9517\ : CascadeMux
    port map (
            O => \N__47014\,
            I => \N__47010\
        );

    \I__9516\ : CascadeMux
    port map (
            O => \N__47013\,
            I => \N__47007\
        );

    \I__9515\ : InMux
    port map (
            O => \N__47010\,
            I => \N__47003\
        );

    \I__9514\ : InMux
    port map (
            O => \N__47007\,
            I => \N__47000\
        );

    \I__9513\ : InMux
    port map (
            O => \N__47006\,
            I => \N__46997\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__47003\,
            I => \N__46994\
        );

    \I__9511\ : LocalMux
    port map (
            O => \N__47000\,
            I => \N__46987\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__46997\,
            I => \N__46987\
        );

    \I__9509\ : Span4Mux_h
    port map (
            O => \N__46994\,
            I => \N__46984\
        );

    \I__9508\ : InMux
    port map (
            O => \N__46993\,
            I => \N__46981\
        );

    \I__9507\ : InMux
    port map (
            O => \N__46992\,
            I => \N__46978\
        );

    \I__9506\ : Span4Mux_h
    port map (
            O => \N__46987\,
            I => \N__46975\
        );

    \I__9505\ : Span4Mux_v
    port map (
            O => \N__46984\,
            I => \N__46972\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__46981\,
            I => data_in_1_4
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__46978\,
            I => data_in_1_4
        );

    \I__9502\ : Odrv4
    port map (
            O => \N__46975\,
            I => data_in_1_4
        );

    \I__9501\ : Odrv4
    port map (
            O => \N__46972\,
            I => data_in_1_4
        );

    \I__9500\ : InMux
    port map (
            O => \N__46963\,
            I => \N__46960\
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__46960\,
            I => \N__46957\
        );

    \I__9498\ : Span4Mux_v
    port map (
            O => \N__46957\,
            I => \N__46954\
        );

    \I__9497\ : Odrv4
    port map (
            O => \N__46954\,
            I => \c0.n6_adj_3343\
        );

    \I__9496\ : InMux
    port map (
            O => \N__46951\,
            I => \N__46948\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__46948\,
            I => \N__46945\
        );

    \I__9494\ : Span12Mux_v
    port map (
            O => \N__46945\,
            I => \N__46942\
        );

    \I__9493\ : Odrv12
    port map (
            O => \N__46942\,
            I => \c0.data_out_frame_28_7\
        );

    \I__9492\ : InMux
    port map (
            O => \N__46939\,
            I => \N__46924\
        );

    \I__9491\ : InMux
    port map (
            O => \N__46938\,
            I => \N__46924\
        );

    \I__9490\ : SRMux
    port map (
            O => \N__46937\,
            I => \N__46911\
        );

    \I__9489\ : CEMux
    port map (
            O => \N__46936\,
            I => \N__46908\
        );

    \I__9488\ : InMux
    port map (
            O => \N__46935\,
            I => \N__46890\
        );

    \I__9487\ : InMux
    port map (
            O => \N__46934\,
            I => \N__46890\
        );

    \I__9486\ : InMux
    port map (
            O => \N__46933\,
            I => \N__46890\
        );

    \I__9485\ : InMux
    port map (
            O => \N__46932\,
            I => \N__46890\
        );

    \I__9484\ : InMux
    port map (
            O => \N__46931\,
            I => \N__46890\
        );

    \I__9483\ : InMux
    port map (
            O => \N__46930\,
            I => \N__46881\
        );

    \I__9482\ : InMux
    port map (
            O => \N__46929\,
            I => \N__46881\
        );

    \I__9481\ : LocalMux
    port map (
            O => \N__46924\,
            I => \N__46878\
        );

    \I__9480\ : InMux
    port map (
            O => \N__46923\,
            I => \N__46867\
        );

    \I__9479\ : InMux
    port map (
            O => \N__46922\,
            I => \N__46867\
        );

    \I__9478\ : InMux
    port map (
            O => \N__46921\,
            I => \N__46867\
        );

    \I__9477\ : InMux
    port map (
            O => \N__46920\,
            I => \N__46867\
        );

    \I__9476\ : InMux
    port map (
            O => \N__46919\,
            I => \N__46867\
        );

    \I__9475\ : InMux
    port map (
            O => \N__46918\,
            I => \N__46861\
        );

    \I__9474\ : CascadeMux
    port map (
            O => \N__46917\,
            I => \N__46852\
        );

    \I__9473\ : CascadeMux
    port map (
            O => \N__46916\,
            I => \N__46849\
        );

    \I__9472\ : InMux
    port map (
            O => \N__46915\,
            I => \N__46843\
        );

    \I__9471\ : InMux
    port map (
            O => \N__46914\,
            I => \N__46843\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__46911\,
            I => \N__46840\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__46908\,
            I => \N__46837\
        );

    \I__9468\ : InMux
    port map (
            O => \N__46907\,
            I => \N__46830\
        );

    \I__9467\ : InMux
    port map (
            O => \N__46906\,
            I => \N__46830\
        );

    \I__9466\ : InMux
    port map (
            O => \N__46905\,
            I => \N__46830\
        );

    \I__9465\ : CascadeMux
    port map (
            O => \N__46904\,
            I => \N__46827\
        );

    \I__9464\ : InMux
    port map (
            O => \N__46903\,
            I => \N__46821\
        );

    \I__9463\ : InMux
    port map (
            O => \N__46902\,
            I => \N__46816\
        );

    \I__9462\ : InMux
    port map (
            O => \N__46901\,
            I => \N__46816\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__46890\,
            I => \N__46813\
        );

    \I__9460\ : InMux
    port map (
            O => \N__46889\,
            I => \N__46810\
        );

    \I__9459\ : InMux
    port map (
            O => \N__46888\,
            I => \N__46807\
        );

    \I__9458\ : InMux
    port map (
            O => \N__46887\,
            I => \N__46804\
        );

    \I__9457\ : InMux
    port map (
            O => \N__46886\,
            I => \N__46800\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__46881\,
            I => \N__46788\
        );

    \I__9455\ : Span4Mux_v
    port map (
            O => \N__46878\,
            I => \N__46788\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__46867\,
            I => \N__46788\
        );

    \I__9453\ : InMux
    port map (
            O => \N__46866\,
            I => \N__46781\
        );

    \I__9452\ : InMux
    port map (
            O => \N__46865\,
            I => \N__46781\
        );

    \I__9451\ : InMux
    port map (
            O => \N__46864\,
            I => \N__46781\
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__46861\,
            I => \N__46776\
        );

    \I__9449\ : InMux
    port map (
            O => \N__46860\,
            I => \N__46773\
        );

    \I__9448\ : InMux
    port map (
            O => \N__46859\,
            I => \N__46770\
        );

    \I__9447\ : CEMux
    port map (
            O => \N__46858\,
            I => \N__46767\
        );

    \I__9446\ : CascadeMux
    port map (
            O => \N__46857\,
            I => \N__46761\
        );

    \I__9445\ : InMux
    port map (
            O => \N__46856\,
            I => \N__46756\
        );

    \I__9444\ : InMux
    port map (
            O => \N__46855\,
            I => \N__46756\
        );

    \I__9443\ : InMux
    port map (
            O => \N__46852\,
            I => \N__46749\
        );

    \I__9442\ : InMux
    port map (
            O => \N__46849\,
            I => \N__46749\
        );

    \I__9441\ : InMux
    port map (
            O => \N__46848\,
            I => \N__46749\
        );

    \I__9440\ : LocalMux
    port map (
            O => \N__46843\,
            I => \N__46744\
        );

    \I__9439\ : Span4Mux_v
    port map (
            O => \N__46840\,
            I => \N__46744\
        );

    \I__9438\ : Span4Mux_v
    port map (
            O => \N__46837\,
            I => \N__46739\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__46830\,
            I => \N__46739\
        );

    \I__9436\ : InMux
    port map (
            O => \N__46827\,
            I => \N__46714\
        );

    \I__9435\ : InMux
    port map (
            O => \N__46826\,
            I => \N__46714\
        );

    \I__9434\ : InMux
    port map (
            O => \N__46825\,
            I => \N__46714\
        );

    \I__9433\ : InMux
    port map (
            O => \N__46824\,
            I => \N__46714\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__46821\,
            I => \N__46709\
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__46816\,
            I => \N__46709\
        );

    \I__9430\ : Span4Mux_h
    port map (
            O => \N__46813\,
            I => \N__46704\
        );

    \I__9429\ : LocalMux
    port map (
            O => \N__46810\,
            I => \N__46704\
        );

    \I__9428\ : LocalMux
    port map (
            O => \N__46807\,
            I => \N__46699\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__46804\,
            I => \N__46699\
        );

    \I__9426\ : SRMux
    port map (
            O => \N__46803\,
            I => \N__46696\
        );

    \I__9425\ : LocalMux
    port map (
            O => \N__46800\,
            I => \N__46693\
        );

    \I__9424\ : InMux
    port map (
            O => \N__46799\,
            I => \N__46688\
        );

    \I__9423\ : InMux
    port map (
            O => \N__46798\,
            I => \N__46683\
        );

    \I__9422\ : InMux
    port map (
            O => \N__46797\,
            I => \N__46683\
        );

    \I__9421\ : InMux
    port map (
            O => \N__46796\,
            I => \N__46678\
        );

    \I__9420\ : InMux
    port map (
            O => \N__46795\,
            I => \N__46678\
        );

    \I__9419\ : Span4Mux_h
    port map (
            O => \N__46788\,
            I => \N__46673\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__46781\,
            I => \N__46673\
        );

    \I__9417\ : InMux
    port map (
            O => \N__46780\,
            I => \N__46668\
        );

    \I__9416\ : InMux
    port map (
            O => \N__46779\,
            I => \N__46668\
        );

    \I__9415\ : Span4Mux_h
    port map (
            O => \N__46776\,
            I => \N__46665\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__46773\,
            I => \N__46658\
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__46770\,
            I => \N__46658\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__46767\,
            I => \N__46658\
        );

    \I__9411\ : CascadeMux
    port map (
            O => \N__46766\,
            I => \N__46655\
        );

    \I__9410\ : CascadeMux
    port map (
            O => \N__46765\,
            I => \N__46652\
        );

    \I__9409\ : InMux
    port map (
            O => \N__46764\,
            I => \N__46639\
        );

    \I__9408\ : InMux
    port map (
            O => \N__46761\,
            I => \N__46636\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__46756\,
            I => \N__46627\
        );

    \I__9406\ : LocalMux
    port map (
            O => \N__46749\,
            I => \N__46627\
        );

    \I__9405\ : Span4Mux_h
    port map (
            O => \N__46744\,
            I => \N__46627\
        );

    \I__9404\ : Span4Mux_h
    port map (
            O => \N__46739\,
            I => \N__46627\
        );

    \I__9403\ : SRMux
    port map (
            O => \N__46738\,
            I => \N__46624\
        );

    \I__9402\ : InMux
    port map (
            O => \N__46737\,
            I => \N__46619\
        );

    \I__9401\ : InMux
    port map (
            O => \N__46736\,
            I => \N__46610\
        );

    \I__9400\ : InMux
    port map (
            O => \N__46735\,
            I => \N__46610\
        );

    \I__9399\ : InMux
    port map (
            O => \N__46734\,
            I => \N__46610\
        );

    \I__9398\ : InMux
    port map (
            O => \N__46733\,
            I => \N__46610\
        );

    \I__9397\ : InMux
    port map (
            O => \N__46732\,
            I => \N__46603\
        );

    \I__9396\ : InMux
    port map (
            O => \N__46731\,
            I => \N__46603\
        );

    \I__9395\ : InMux
    port map (
            O => \N__46730\,
            I => \N__46603\
        );

    \I__9394\ : SRMux
    port map (
            O => \N__46729\,
            I => \N__46600\
        );

    \I__9393\ : InMux
    port map (
            O => \N__46728\,
            I => \N__46593\
        );

    \I__9392\ : InMux
    port map (
            O => \N__46727\,
            I => \N__46593\
        );

    \I__9391\ : InMux
    port map (
            O => \N__46726\,
            I => \N__46593\
        );

    \I__9390\ : InMux
    port map (
            O => \N__46725\,
            I => \N__46588\
        );

    \I__9389\ : InMux
    port map (
            O => \N__46724\,
            I => \N__46588\
        );

    \I__9388\ : InMux
    port map (
            O => \N__46723\,
            I => \N__46585\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__46714\,
            I => \N__46582\
        );

    \I__9386\ : Span4Mux_v
    port map (
            O => \N__46709\,
            I => \N__46577\
        );

    \I__9385\ : Span4Mux_v
    port map (
            O => \N__46704\,
            I => \N__46577\
        );

    \I__9384\ : Span4Mux_v
    port map (
            O => \N__46699\,
            I => \N__46572\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__46696\,
            I => \N__46572\
        );

    \I__9382\ : Span4Mux_v
    port map (
            O => \N__46693\,
            I => \N__46569\
        );

    \I__9381\ : InMux
    port map (
            O => \N__46692\,
            I => \N__46564\
        );

    \I__9380\ : InMux
    port map (
            O => \N__46691\,
            I => \N__46564\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__46688\,
            I => \N__46549\
        );

    \I__9378\ : LocalMux
    port map (
            O => \N__46683\,
            I => \N__46549\
        );

    \I__9377\ : LocalMux
    port map (
            O => \N__46678\,
            I => \N__46549\
        );

    \I__9376\ : Span4Mux_h
    port map (
            O => \N__46673\,
            I => \N__46549\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__46668\,
            I => \N__46549\
        );

    \I__9374\ : Span4Mux_h
    port map (
            O => \N__46665\,
            I => \N__46549\
        );

    \I__9373\ : Span4Mux_h
    port map (
            O => \N__46658\,
            I => \N__46549\
        );

    \I__9372\ : InMux
    port map (
            O => \N__46655\,
            I => \N__46542\
        );

    \I__9371\ : InMux
    port map (
            O => \N__46652\,
            I => \N__46542\
        );

    \I__9370\ : InMux
    port map (
            O => \N__46651\,
            I => \N__46542\
        );

    \I__9369\ : InMux
    port map (
            O => \N__46650\,
            I => \N__46531\
        );

    \I__9368\ : InMux
    port map (
            O => \N__46649\,
            I => \N__46531\
        );

    \I__9367\ : InMux
    port map (
            O => \N__46648\,
            I => \N__46531\
        );

    \I__9366\ : InMux
    port map (
            O => \N__46647\,
            I => \N__46531\
        );

    \I__9365\ : InMux
    port map (
            O => \N__46646\,
            I => \N__46531\
        );

    \I__9364\ : InMux
    port map (
            O => \N__46645\,
            I => \N__46526\
        );

    \I__9363\ : InMux
    port map (
            O => \N__46644\,
            I => \N__46526\
        );

    \I__9362\ : InMux
    port map (
            O => \N__46643\,
            I => \N__46523\
        );

    \I__9361\ : InMux
    port map (
            O => \N__46642\,
            I => \N__46520\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__46639\,
            I => \N__46513\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__46636\,
            I => \N__46513\
        );

    \I__9358\ : Span4Mux_v
    port map (
            O => \N__46627\,
            I => \N__46513\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__46624\,
            I => \N__46510\
        );

    \I__9356\ : InMux
    port map (
            O => \N__46623\,
            I => \N__46505\
        );

    \I__9355\ : InMux
    port map (
            O => \N__46622\,
            I => \N__46505\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__46619\,
            I => \N__46498\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__46610\,
            I => \N__46498\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__46603\,
            I => \N__46498\
        );

    \I__9351\ : LocalMux
    port map (
            O => \N__46600\,
            I => \N__46495\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__46593\,
            I => \N__46490\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__46588\,
            I => \N__46490\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__46585\,
            I => \N__46485\
        );

    \I__9347\ : Span4Mux_v
    port map (
            O => \N__46582\,
            I => \N__46485\
        );

    \I__9346\ : Span4Mux_v
    port map (
            O => \N__46577\,
            I => \N__46478\
        );

    \I__9345\ : Span4Mux_v
    port map (
            O => \N__46572\,
            I => \N__46478\
        );

    \I__9344\ : Span4Mux_h
    port map (
            O => \N__46569\,
            I => \N__46478\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__46564\,
            I => \N__46473\
        );

    \I__9342\ : Sp12to4
    port map (
            O => \N__46549\,
            I => \N__46473\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__46542\,
            I => \N__46468\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__46531\,
            I => \N__46468\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__46526\,
            I => \N__46463\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__46523\,
            I => \N__46463\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__46520\,
            I => \N__46458\
        );

    \I__9336\ : Span4Mux_v
    port map (
            O => \N__46513\,
            I => \N__46458\
        );

    \I__9335\ : Span4Mux_v
    port map (
            O => \N__46510\,
            I => \N__46455\
        );

    \I__9334\ : LocalMux
    port map (
            O => \N__46505\,
            I => \N__46450\
        );

    \I__9333\ : Span4Mux_v
    port map (
            O => \N__46498\,
            I => \N__46450\
        );

    \I__9332\ : Span4Mux_h
    port map (
            O => \N__46495\,
            I => \N__46443\
        );

    \I__9331\ : Span4Mux_v
    port map (
            O => \N__46490\,
            I => \N__46443\
        );

    \I__9330\ : Span4Mux_h
    port map (
            O => \N__46485\,
            I => \N__46443\
        );

    \I__9329\ : Sp12to4
    port map (
            O => \N__46478\,
            I => \N__46438\
        );

    \I__9328\ : Span12Mux_v
    port map (
            O => \N__46473\,
            I => \N__46438\
        );

    \I__9327\ : Span4Mux_v
    port map (
            O => \N__46468\,
            I => \N__46431\
        );

    \I__9326\ : Span4Mux_h
    port map (
            O => \N__46463\,
            I => \N__46431\
        );

    \I__9325\ : Span4Mux_h
    port map (
            O => \N__46458\,
            I => \N__46431\
        );

    \I__9324\ : Odrv4
    port map (
            O => \N__46455\,
            I => n8112
        );

    \I__9323\ : Odrv4
    port map (
            O => \N__46450\,
            I => n8112
        );

    \I__9322\ : Odrv4
    port map (
            O => \N__46443\,
            I => n8112
        );

    \I__9321\ : Odrv12
    port map (
            O => \N__46438\,
            I => n8112
        );

    \I__9320\ : Odrv4
    port map (
            O => \N__46431\,
            I => n8112
        );

    \I__9319\ : CascadeMux
    port map (
            O => \N__46420\,
            I => \N__46417\
        );

    \I__9318\ : InMux
    port map (
            O => \N__46417\,
            I => \N__46411\
        );

    \I__9317\ : InMux
    port map (
            O => \N__46416\,
            I => \N__46408\
        );

    \I__9316\ : InMux
    port map (
            O => \N__46415\,
            I => \N__46405\
        );

    \I__9315\ : InMux
    port map (
            O => \N__46414\,
            I => \N__46402\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__46411\,
            I => \c0.data_in_frame_4_3\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__46408\,
            I => \c0.data_in_frame_4_3\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__46405\,
            I => \c0.data_in_frame_4_3\
        );

    \I__9311\ : LocalMux
    port map (
            O => \N__46402\,
            I => \c0.data_in_frame_4_3\
        );

    \I__9310\ : InMux
    port map (
            O => \N__46393\,
            I => \N__46387\
        );

    \I__9309\ : InMux
    port map (
            O => \N__46392\,
            I => \N__46384\
        );

    \I__9308\ : InMux
    port map (
            O => \N__46391\,
            I => \N__46381\
        );

    \I__9307\ : InMux
    port map (
            O => \N__46390\,
            I => \N__46378\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__46387\,
            I => \c0.data_in_frame_4_2\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__46384\,
            I => \c0.data_in_frame_4_2\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__46381\,
            I => \c0.data_in_frame_4_2\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__46378\,
            I => \c0.data_in_frame_4_2\
        );

    \I__9302\ : CascadeMux
    port map (
            O => \N__46369\,
            I => \N__46365\
        );

    \I__9301\ : CascadeMux
    port map (
            O => \N__46368\,
            I => \N__46362\
        );

    \I__9300\ : InMux
    port map (
            O => \N__46365\,
            I => \N__46359\
        );

    \I__9299\ : InMux
    port map (
            O => \N__46362\,
            I => \N__46356\
        );

    \I__9298\ : LocalMux
    port map (
            O => \N__46359\,
            I => \N__46351\
        );

    \I__9297\ : LocalMux
    port map (
            O => \N__46356\,
            I => \N__46351\
        );

    \I__9296\ : Odrv12
    port map (
            O => \N__46351\,
            I => \c0.data_in_frame_6_4\
        );

    \I__9295\ : CascadeMux
    port map (
            O => \N__46348\,
            I => \c0.n13_adj_3496_cascade_\
        );

    \I__9294\ : CascadeMux
    port map (
            O => \N__46345\,
            I => \N__46342\
        );

    \I__9293\ : InMux
    port map (
            O => \N__46342\,
            I => \N__46338\
        );

    \I__9292\ : InMux
    port map (
            O => \N__46341\,
            I => \N__46335\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__46338\,
            I => \N__46330\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__46335\,
            I => \N__46327\
        );

    \I__9289\ : InMux
    port map (
            O => \N__46334\,
            I => \N__46324\
        );

    \I__9288\ : InMux
    port map (
            O => \N__46333\,
            I => \N__46321\
        );

    \I__9287\ : Span4Mux_h
    port map (
            O => \N__46330\,
            I => \N__46318\
        );

    \I__9286\ : Span4Mux_h
    port map (
            O => \N__46327\,
            I => \N__46315\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__46324\,
            I => \N__46312\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__46321\,
            I => \c0.data_in_frame_2_2\
        );

    \I__9283\ : Odrv4
    port map (
            O => \N__46318\,
            I => \c0.data_in_frame_2_2\
        );

    \I__9282\ : Odrv4
    port map (
            O => \N__46315\,
            I => \c0.data_in_frame_2_2\
        );

    \I__9281\ : Odrv12
    port map (
            O => \N__46312\,
            I => \c0.data_in_frame_2_2\
        );

    \I__9280\ : InMux
    port map (
            O => \N__46303\,
            I => \N__46297\
        );

    \I__9279\ : InMux
    port map (
            O => \N__46302\,
            I => \N__46294\
        );

    \I__9278\ : InMux
    port map (
            O => \N__46301\,
            I => \N__46289\
        );

    \I__9277\ : CascadeMux
    port map (
            O => \N__46300\,
            I => \N__46284\
        );

    \I__9276\ : LocalMux
    port map (
            O => \N__46297\,
            I => \N__46280\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__46294\,
            I => \N__46277\
        );

    \I__9274\ : CascadeMux
    port map (
            O => \N__46293\,
            I => \N__46274\
        );

    \I__9273\ : CascadeMux
    port map (
            O => \N__46292\,
            I => \N__46270\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__46289\,
            I => \N__46266\
        );

    \I__9271\ : CascadeMux
    port map (
            O => \N__46288\,
            I => \N__46262\
        );

    \I__9270\ : InMux
    port map (
            O => \N__46287\,
            I => \N__46257\
        );

    \I__9269\ : InMux
    port map (
            O => \N__46284\,
            I => \N__46257\
        );

    \I__9268\ : InMux
    port map (
            O => \N__46283\,
            I => \N__46254\
        );

    \I__9267\ : Span4Mux_v
    port map (
            O => \N__46280\,
            I => \N__46251\
        );

    \I__9266\ : Span4Mux_h
    port map (
            O => \N__46277\,
            I => \N__46248\
        );

    \I__9265\ : InMux
    port map (
            O => \N__46274\,
            I => \N__46241\
        );

    \I__9264\ : InMux
    port map (
            O => \N__46273\,
            I => \N__46241\
        );

    \I__9263\ : InMux
    port map (
            O => \N__46270\,
            I => \N__46241\
        );

    \I__9262\ : InMux
    port map (
            O => \N__46269\,
            I => \N__46238\
        );

    \I__9261\ : Span4Mux_h
    port map (
            O => \N__46266\,
            I => \N__46235\
        );

    \I__9260\ : InMux
    port map (
            O => \N__46265\,
            I => \N__46230\
        );

    \I__9259\ : InMux
    port map (
            O => \N__46262\,
            I => \N__46230\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__46257\,
            I => data_in_frame_0_0
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__46254\,
            I => data_in_frame_0_0
        );

    \I__9256\ : Odrv4
    port map (
            O => \N__46251\,
            I => data_in_frame_0_0
        );

    \I__9255\ : Odrv4
    port map (
            O => \N__46248\,
            I => data_in_frame_0_0
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__46241\,
            I => data_in_frame_0_0
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__46238\,
            I => data_in_frame_0_0
        );

    \I__9252\ : Odrv4
    port map (
            O => \N__46235\,
            I => data_in_frame_0_0
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__46230\,
            I => data_in_frame_0_0
        );

    \I__9250\ : InMux
    port map (
            O => \N__46213\,
            I => \N__46210\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__46210\,
            I => \c0.n19277\
        );

    \I__9248\ : InMux
    port map (
            O => \N__46207\,
            I => \N__46203\
        );

    \I__9247\ : CascadeMux
    port map (
            O => \N__46206\,
            I => \N__46200\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__46203\,
            I => \N__46197\
        );

    \I__9245\ : InMux
    port map (
            O => \N__46200\,
            I => \N__46194\
        );

    \I__9244\ : Odrv4
    port map (
            O => \N__46197\,
            I => \c0.n7_adj_3078\
        );

    \I__9243\ : LocalMux
    port map (
            O => \N__46194\,
            I => \c0.n7_adj_3078\
        );

    \I__9242\ : InMux
    port map (
            O => \N__46189\,
            I => \N__46186\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__46186\,
            I => \N__46183\
        );

    \I__9240\ : Span4Mux_v
    port map (
            O => \N__46183\,
            I => \N__46180\
        );

    \I__9239\ : Odrv4
    port map (
            O => \N__46180\,
            I => \c0.n17880\
        );

    \I__9238\ : InMux
    port map (
            O => \N__46177\,
            I => \N__46174\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__46174\,
            I => \N__46171\
        );

    \I__9236\ : Odrv4
    port map (
            O => \N__46171\,
            I => \c0.n26_adj_3523\
        );

    \I__9235\ : CascadeMux
    port map (
            O => \N__46168\,
            I => \N__46164\
        );

    \I__9234\ : InMux
    port map (
            O => \N__46167\,
            I => \N__46161\
        );

    \I__9233\ : InMux
    port map (
            O => \N__46164\,
            I => \N__46158\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__46161\,
            I => data_in_0_4
        );

    \I__9231\ : LocalMux
    port map (
            O => \N__46158\,
            I => data_in_0_4
        );

    \I__9230\ : InMux
    port map (
            O => \N__46153\,
            I => \N__46149\
        );

    \I__9229\ : InMux
    port map (
            O => \N__46152\,
            I => \N__46146\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__46149\,
            I => \N__46143\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__46146\,
            I => \N__46140\
        );

    \I__9226\ : Span4Mux_h
    port map (
            O => \N__46143\,
            I => \N__46131\
        );

    \I__9225\ : Span4Mux_v
    port map (
            O => \N__46140\,
            I => \N__46128\
        );

    \I__9224\ : InMux
    port map (
            O => \N__46139\,
            I => \N__46125\
        );

    \I__9223\ : InMux
    port map (
            O => \N__46138\,
            I => \N__46116\
        );

    \I__9222\ : InMux
    port map (
            O => \N__46137\,
            I => \N__46116\
        );

    \I__9221\ : InMux
    port map (
            O => \N__46136\,
            I => \N__46116\
        );

    \I__9220\ : InMux
    port map (
            O => \N__46135\,
            I => \N__46116\
        );

    \I__9219\ : InMux
    port map (
            O => \N__46134\,
            I => \N__46113\
        );

    \I__9218\ : Odrv4
    port map (
            O => \N__46131\,
            I => n20896
        );

    \I__9217\ : Odrv4
    port map (
            O => \N__46128\,
            I => n20896
        );

    \I__9216\ : LocalMux
    port map (
            O => \N__46125\,
            I => n20896
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__46116\,
            I => n20896
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__46113\,
            I => n20896
        );

    \I__9213\ : InMux
    port map (
            O => \N__46102\,
            I => \N__46099\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__46099\,
            I => \c0.n18457\
        );

    \I__9211\ : InMux
    port map (
            O => \N__46096\,
            I => \N__46090\
        );

    \I__9210\ : InMux
    port map (
            O => \N__46095\,
            I => \N__46087\
        );

    \I__9209\ : InMux
    port map (
            O => \N__46094\,
            I => \N__46084\
        );

    \I__9208\ : InMux
    port map (
            O => \N__46093\,
            I => \N__46081\
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__46090\,
            I => \N__46078\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__46087\,
            I => \N__46075\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__46084\,
            I => \c0.n21076\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__46081\,
            I => \c0.n21076\
        );

    \I__9203\ : Odrv4
    port map (
            O => \N__46078\,
            I => \c0.n21076\
        );

    \I__9202\ : Odrv4
    port map (
            O => \N__46075\,
            I => \c0.n21076\
        );

    \I__9201\ : InMux
    port map (
            O => \N__46066\,
            I => \N__46063\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__46063\,
            I => \N__46060\
        );

    \I__9199\ : Odrv12
    port map (
            O => \N__46060\,
            I => \c0.n33_adj_3308\
        );

    \I__9198\ : CascadeMux
    port map (
            O => \N__46057\,
            I => \N__46054\
        );

    \I__9197\ : InMux
    port map (
            O => \N__46054\,
            I => \N__46048\
        );

    \I__9196\ : InMux
    port map (
            O => \N__46053\,
            I => \N__46048\
        );

    \I__9195\ : LocalMux
    port map (
            O => \N__46048\,
            I => \c0.n18417\
        );

    \I__9194\ : CascadeMux
    port map (
            O => \N__46045\,
            I => \c0.n18417_cascade_\
        );

    \I__9193\ : InMux
    port map (
            O => \N__46042\,
            I => \N__46039\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__46039\,
            I => \c0.n19_adj_3292\
        );

    \I__9191\ : InMux
    port map (
            O => \N__46036\,
            I => \N__46030\
        );

    \I__9190\ : InMux
    port map (
            O => \N__46035\,
            I => \N__46030\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__46030\,
            I => \c0.data_in_frame_29_4\
        );

    \I__9188\ : InMux
    port map (
            O => \N__46027\,
            I => \N__46024\
        );

    \I__9187\ : LocalMux
    port map (
            O => \N__46024\,
            I => \N__46020\
        );

    \I__9186\ : CascadeMux
    port map (
            O => \N__46023\,
            I => \N__46017\
        );

    \I__9185\ : Span4Mux_h
    port map (
            O => \N__46020\,
            I => \N__46014\
        );

    \I__9184\ : InMux
    port map (
            O => \N__46017\,
            I => \N__46011\
        );

    \I__9183\ : Span4Mux_v
    port map (
            O => \N__46014\,
            I => \N__46008\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__46011\,
            I => \c0.data_in_frame_29_2\
        );

    \I__9181\ : Odrv4
    port map (
            O => \N__46008\,
            I => \c0.data_in_frame_29_2\
        );

    \I__9180\ : InMux
    port map (
            O => \N__46003\,
            I => \N__46000\
        );

    \I__9179\ : LocalMux
    port map (
            O => \N__46000\,
            I => \N__45996\
        );

    \I__9178\ : InMux
    port map (
            O => \N__45999\,
            I => \N__45993\
        );

    \I__9177\ : Span4Mux_h
    port map (
            O => \N__45996\,
            I => \N__45990\
        );

    \I__9176\ : LocalMux
    port map (
            O => \N__45993\,
            I => \c0.data_in_frame_29_1\
        );

    \I__9175\ : Odrv4
    port map (
            O => \N__45990\,
            I => \c0.data_in_frame_29_1\
        );

    \I__9174\ : CascadeMux
    port map (
            O => \N__45985\,
            I => \N__45982\
        );

    \I__9173\ : InMux
    port map (
            O => \N__45982\,
            I => \N__45979\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__45979\,
            I => \N__45976\
        );

    \I__9171\ : Span4Mux_v
    port map (
            O => \N__45976\,
            I => \N__45972\
        );

    \I__9170\ : InMux
    port map (
            O => \N__45975\,
            I => \N__45969\
        );

    \I__9169\ : Span4Mux_v
    port map (
            O => \N__45972\,
            I => \N__45966\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__45969\,
            I => \N__45963\
        );

    \I__9167\ : Span4Mux_h
    port map (
            O => \N__45966\,
            I => \N__45960\
        );

    \I__9166\ : Odrv4
    port map (
            O => \N__45963\,
            I => \c0.data_in_frame_28_1\
        );

    \I__9165\ : Odrv4
    port map (
            O => \N__45960\,
            I => \c0.data_in_frame_28_1\
        );

    \I__9164\ : CascadeMux
    port map (
            O => \N__45955\,
            I => \N__45951\
        );

    \I__9163\ : CascadeMux
    port map (
            O => \N__45954\,
            I => \N__45948\
        );

    \I__9162\ : InMux
    port map (
            O => \N__45951\,
            I => \N__45945\
        );

    \I__9161\ : InMux
    port map (
            O => \N__45948\,
            I => \N__45942\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__45945\,
            I => \c0.data_in_frame_28_0\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__45942\,
            I => \c0.data_in_frame_28_0\
        );

    \I__9158\ : InMux
    port map (
            O => \N__45937\,
            I => \N__45932\
        );

    \I__9157\ : InMux
    port map (
            O => \N__45936\,
            I => \N__45926\
        );

    \I__9156\ : InMux
    port map (
            O => \N__45935\,
            I => \N__45923\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__45932\,
            I => \N__45920\
        );

    \I__9154\ : CascadeMux
    port map (
            O => \N__45931\,
            I => \N__45917\
        );

    \I__9153\ : InMux
    port map (
            O => \N__45930\,
            I => \N__45912\
        );

    \I__9152\ : InMux
    port map (
            O => \N__45929\,
            I => \N__45912\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__45926\,
            I => \N__45909\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__45923\,
            I => \N__45906\
        );

    \I__9149\ : Span4Mux_h
    port map (
            O => \N__45920\,
            I => \N__45903\
        );

    \I__9148\ : InMux
    port map (
            O => \N__45917\,
            I => \N__45900\
        );

    \I__9147\ : LocalMux
    port map (
            O => \N__45912\,
            I => \c0.n20324\
        );

    \I__9146\ : Odrv4
    port map (
            O => \N__45909\,
            I => \c0.n20324\
        );

    \I__9145\ : Odrv12
    port map (
            O => \N__45906\,
            I => \c0.n20324\
        );

    \I__9144\ : Odrv4
    port map (
            O => \N__45903\,
            I => \c0.n20324\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__45900\,
            I => \c0.n20324\
        );

    \I__9142\ : InMux
    port map (
            O => \N__45889\,
            I => \N__45886\
        );

    \I__9141\ : LocalMux
    port map (
            O => \N__45886\,
            I => \N__45883\
        );

    \I__9140\ : Odrv4
    port map (
            O => \N__45883\,
            I => \c0.n14_adj_3349\
        );

    \I__9139\ : CascadeMux
    port map (
            O => \N__45880\,
            I => \c0.n21044_cascade_\
        );

    \I__9138\ : InMux
    port map (
            O => \N__45877\,
            I => \N__45871\
        );

    \I__9137\ : InMux
    port map (
            O => \N__45876\,
            I => \N__45871\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__45871\,
            I => \N__45865\
        );

    \I__9135\ : CascadeMux
    port map (
            O => \N__45870\,
            I => \N__45862\
        );

    \I__9134\ : InMux
    port map (
            O => \N__45869\,
            I => \N__45859\
        );

    \I__9133\ : CascadeMux
    port map (
            O => \N__45868\,
            I => \N__45856\
        );

    \I__9132\ : Span4Mux_v
    port map (
            O => \N__45865\,
            I => \N__45853\
        );

    \I__9131\ : InMux
    port map (
            O => \N__45862\,
            I => \N__45850\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__45859\,
            I => \N__45847\
        );

    \I__9129\ : InMux
    port map (
            O => \N__45856\,
            I => \N__45844\
        );

    \I__9128\ : Span4Mux_h
    port map (
            O => \N__45853\,
            I => \N__45841\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__45850\,
            I => \N__45836\
        );

    \I__9126\ : Span4Mux_h
    port map (
            O => \N__45847\,
            I => \N__45836\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__45844\,
            I => \c0.data_in_frame_26_7\
        );

    \I__9124\ : Odrv4
    port map (
            O => \N__45841\,
            I => \c0.data_in_frame_26_7\
        );

    \I__9123\ : Odrv4
    port map (
            O => \N__45836\,
            I => \c0.data_in_frame_26_7\
        );

    \I__9122\ : CascadeMux
    port map (
            O => \N__45829\,
            I => \c0.n16_adj_3109_cascade_\
        );

    \I__9121\ : InMux
    port map (
            O => \N__45826\,
            I => \N__45822\
        );

    \I__9120\ : InMux
    port map (
            O => \N__45825\,
            I => \N__45819\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__45822\,
            I => \c0.n21071\
        );

    \I__9118\ : LocalMux
    port map (
            O => \N__45819\,
            I => \c0.n21071\
        );

    \I__9117\ : CascadeMux
    port map (
            O => \N__45814\,
            I => \N__45811\
        );

    \I__9116\ : InMux
    port map (
            O => \N__45811\,
            I => \N__45805\
        );

    \I__9115\ : InMux
    port map (
            O => \N__45810\,
            I => \N__45805\
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__45805\,
            I => \N__45801\
        );

    \I__9113\ : InMux
    port map (
            O => \N__45804\,
            I => \N__45798\
        );

    \I__9112\ : Span4Mux_v
    port map (
            O => \N__45801\,
            I => \N__45793\
        );

    \I__9111\ : LocalMux
    port map (
            O => \N__45798\,
            I => \N__45793\
        );

    \I__9110\ : Odrv4
    port map (
            O => \N__45793\,
            I => \c0.n20479\
        );

    \I__9109\ : InMux
    port map (
            O => \N__45790\,
            I => \N__45787\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__45787\,
            I => \c0.n77\
        );

    \I__9107\ : InMux
    port map (
            O => \N__45784\,
            I => \N__45781\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__45781\,
            I => \N__45777\
        );

    \I__9105\ : InMux
    port map (
            O => \N__45780\,
            I => \N__45774\
        );

    \I__9104\ : Span4Mux_h
    port map (
            O => \N__45777\,
            I => \N__45771\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__45774\,
            I => \c0.n34_adj_3096\
        );

    \I__9102\ : Odrv4
    port map (
            O => \N__45771\,
            I => \c0.n34_adj_3096\
        );

    \I__9101\ : InMux
    port map (
            O => \N__45766\,
            I => \N__45762\
        );

    \I__9100\ : InMux
    port map (
            O => \N__45765\,
            I => \N__45759\
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__45762\,
            I => \N__45756\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__45759\,
            I => \N__45753\
        );

    \I__9097\ : Odrv12
    port map (
            O => \N__45756\,
            I => \c0.n32_adj_3095\
        );

    \I__9096\ : Odrv4
    port map (
            O => \N__45753\,
            I => \c0.n32_adj_3095\
        );

    \I__9095\ : CascadeMux
    port map (
            O => \N__45748\,
            I => \c0.n18457_cascade_\
        );

    \I__9094\ : InMux
    port map (
            O => \N__45745\,
            I => \N__45741\
        );

    \I__9093\ : InMux
    port map (
            O => \N__45744\,
            I => \N__45738\
        );

    \I__9092\ : LocalMux
    port map (
            O => \N__45741\,
            I => \c0.n23_adj_3222\
        );

    \I__9091\ : LocalMux
    port map (
            O => \N__45738\,
            I => \c0.n23_adj_3222\
        );

    \I__9090\ : CascadeMux
    port map (
            O => \N__45733\,
            I => \c0.n43_adj_3280_cascade_\
        );

    \I__9089\ : InMux
    port map (
            O => \N__45730\,
            I => \N__45727\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__45727\,
            I => \c0.n41_adj_3281\
        );

    \I__9087\ : InMux
    port map (
            O => \N__45724\,
            I => \N__45721\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__45721\,
            I => \c0.n50_adj_3283\
        );

    \I__9085\ : CascadeMux
    port map (
            O => \N__45718\,
            I => \c0.n19511_cascade_\
        );

    \I__9084\ : InMux
    port map (
            O => \N__45715\,
            I => \N__45710\
        );

    \I__9083\ : InMux
    port map (
            O => \N__45714\,
            I => \N__45705\
        );

    \I__9082\ : InMux
    port map (
            O => \N__45713\,
            I => \N__45705\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__45710\,
            I => \N__45699\
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__45705\,
            I => \N__45696\
        );

    \I__9079\ : InMux
    port map (
            O => \N__45704\,
            I => \N__45691\
        );

    \I__9078\ : InMux
    port map (
            O => \N__45703\,
            I => \N__45691\
        );

    \I__9077\ : InMux
    port map (
            O => \N__45702\,
            I => \N__45688\
        );

    \I__9076\ : Span4Mux_v
    port map (
            O => \N__45699\,
            I => \N__45685\
        );

    \I__9075\ : Sp12to4
    port map (
            O => \N__45696\,
            I => \N__45680\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__45691\,
            I => \N__45680\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__45688\,
            I => \c0.n21110\
        );

    \I__9072\ : Odrv4
    port map (
            O => \N__45685\,
            I => \c0.n21110\
        );

    \I__9071\ : Odrv12
    port map (
            O => \N__45680\,
            I => \c0.n21110\
        );

    \I__9070\ : InMux
    port map (
            O => \N__45673\,
            I => \N__45670\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__45670\,
            I => \N__45667\
        );

    \I__9068\ : Span12Mux_v
    port map (
            O => \N__45667\,
            I => \N__45664\
        );

    \I__9067\ : Odrv12
    port map (
            O => \N__45664\,
            I => \c0.n20_adj_3448\
        );

    \I__9066\ : InMux
    port map (
            O => \N__45661\,
            I => \N__45657\
        );

    \I__9065\ : InMux
    port map (
            O => \N__45660\,
            I => \N__45654\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__45657\,
            I => \c0.n20431\
        );

    \I__9063\ : LocalMux
    port map (
            O => \N__45654\,
            I => \c0.n20431\
        );

    \I__9062\ : InMux
    port map (
            O => \N__45649\,
            I => \N__45646\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__45646\,
            I => \N__45643\
        );

    \I__9060\ : Odrv12
    port map (
            O => \N__45643\,
            I => \c0.n64_adj_3512\
        );

    \I__9059\ : InMux
    port map (
            O => \N__45640\,
            I => \N__45634\
        );

    \I__9058\ : CascadeMux
    port map (
            O => \N__45639\,
            I => \N__45630\
        );

    \I__9057\ : InMux
    port map (
            O => \N__45638\,
            I => \N__45626\
        );

    \I__9056\ : InMux
    port map (
            O => \N__45637\,
            I => \N__45623\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__45634\,
            I => \N__45620\
        );

    \I__9054\ : InMux
    port map (
            O => \N__45633\,
            I => \N__45613\
        );

    \I__9053\ : InMux
    port map (
            O => \N__45630\,
            I => \N__45613\
        );

    \I__9052\ : InMux
    port map (
            O => \N__45629\,
            I => \N__45613\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__45626\,
            I => \N__45609\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__45623\,
            I => \N__45606\
        );

    \I__9049\ : Span4Mux_v
    port map (
            O => \N__45620\,
            I => \N__45603\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__45613\,
            I => \N__45600\
        );

    \I__9047\ : InMux
    port map (
            O => \N__45612\,
            I => \N__45597\
        );

    \I__9046\ : Span4Mux_h
    port map (
            O => \N__45609\,
            I => \N__45594\
        );

    \I__9045\ : Span12Mux_h
    port map (
            O => \N__45606\,
            I => \N__45591\
        );

    \I__9044\ : Span4Mux_v
    port map (
            O => \N__45603\,
            I => \N__45586\
        );

    \I__9043\ : Span4Mux_h
    port map (
            O => \N__45600\,
            I => \N__45586\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__45597\,
            I => data_in_frame_16_4
        );

    \I__9041\ : Odrv4
    port map (
            O => \N__45594\,
            I => data_in_frame_16_4
        );

    \I__9040\ : Odrv12
    port map (
            O => \N__45591\,
            I => data_in_frame_16_4
        );

    \I__9039\ : Odrv4
    port map (
            O => \N__45586\,
            I => data_in_frame_16_4
        );

    \I__9038\ : InMux
    port map (
            O => \N__45577\,
            I => \N__45574\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__45574\,
            I => \N__45571\
        );

    \I__9036\ : Span4Mux_v
    port map (
            O => \N__45571\,
            I => \N__45568\
        );

    \I__9035\ : Odrv4
    port map (
            O => \N__45568\,
            I => \c0.n7_adj_3440\
        );

    \I__9034\ : InMux
    port map (
            O => \N__45565\,
            I => \N__45561\
        );

    \I__9033\ : InMux
    port map (
            O => \N__45564\,
            I => \N__45557\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__45561\,
            I => \N__45554\
        );

    \I__9031\ : InMux
    port map (
            O => \N__45560\,
            I => \N__45551\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__45557\,
            I => \N__45546\
        );

    \I__9029\ : Span4Mux_v
    port map (
            O => \N__45554\,
            I => \N__45546\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__45551\,
            I => \c0.data_in_frame_13_0\
        );

    \I__9027\ : Odrv4
    port map (
            O => \N__45546\,
            I => \c0.data_in_frame_13_0\
        );

    \I__9026\ : CascadeMux
    port map (
            O => \N__45541\,
            I => \N__45538\
        );

    \I__9025\ : InMux
    port map (
            O => \N__45538\,
            I => \N__45535\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__45535\,
            I => \N__45532\
        );

    \I__9023\ : Span4Mux_h
    port map (
            O => \N__45532\,
            I => \N__45529\
        );

    \I__9022\ : Span4Mux_v
    port map (
            O => \N__45529\,
            I => \N__45526\
        );

    \I__9021\ : Odrv4
    port map (
            O => \N__45526\,
            I => \c0.n11_adj_3219\
        );

    \I__9020\ : InMux
    port map (
            O => \N__45523\,
            I => \N__45520\
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__45520\,
            I => \N__45517\
        );

    \I__9018\ : Odrv12
    port map (
            O => \N__45517\,
            I => \c0.n13_adj_3221\
        );

    \I__9017\ : InMux
    port map (
            O => \N__45514\,
            I => \N__45511\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__45511\,
            I => \N__45506\
        );

    \I__9015\ : InMux
    port map (
            O => \N__45510\,
            I => \N__45501\
        );

    \I__9014\ : InMux
    port map (
            O => \N__45509\,
            I => \N__45501\
        );

    \I__9013\ : Odrv4
    port map (
            O => \N__45506\,
            I => data_in_frame_23_3
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__45501\,
            I => data_in_frame_23_3
        );

    \I__9011\ : InMux
    port map (
            O => \N__45496\,
            I => \N__45493\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__45493\,
            I => \c0.n25_adj_3524\
        );

    \I__9009\ : InMux
    port map (
            O => \N__45490\,
            I => \N__45487\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__45487\,
            I => \c0.n19384\
        );

    \I__9007\ : InMux
    port map (
            O => \N__45484\,
            I => \N__45481\
        );

    \I__9006\ : LocalMux
    port map (
            O => \N__45481\,
            I => \N__45478\
        );

    \I__9005\ : Odrv4
    port map (
            O => \N__45478\,
            I => \c0.n13_adj_3463\
        );

    \I__9004\ : InMux
    port map (
            O => \N__45475\,
            I => \N__45472\
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__45472\,
            I => \N__45469\
        );

    \I__9002\ : Span4Mux_v
    port map (
            O => \N__45469\,
            I => \N__45466\
        );

    \I__9001\ : Odrv4
    port map (
            O => \N__45466\,
            I => \c0.n10\
        );

    \I__9000\ : CascadeMux
    port map (
            O => \N__45463\,
            I => \c0.n19384_cascade_\
        );

    \I__8999\ : InMux
    port map (
            O => \N__45460\,
            I => \N__45453\
        );

    \I__8998\ : InMux
    port map (
            O => \N__45459\,
            I => \N__45453\
        );

    \I__8997\ : CascadeMux
    port map (
            O => \N__45458\,
            I => \N__45449\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__45453\,
            I => \N__45446\
        );

    \I__8995\ : CascadeMux
    port map (
            O => \N__45452\,
            I => \N__45443\
        );

    \I__8994\ : InMux
    port map (
            O => \N__45449\,
            I => \N__45440\
        );

    \I__8993\ : Span4Mux_v
    port map (
            O => \N__45446\,
            I => \N__45437\
        );

    \I__8992\ : InMux
    port map (
            O => \N__45443\,
            I => \N__45434\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__45440\,
            I => \N__45430\
        );

    \I__8990\ : Span4Mux_v
    port map (
            O => \N__45437\,
            I => \N__45425\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__45434\,
            I => \N__45425\
        );

    \I__8988\ : InMux
    port map (
            O => \N__45433\,
            I => \N__45422\
        );

    \I__8987\ : Span4Mux_h
    port map (
            O => \N__45430\,
            I => \N__45417\
        );

    \I__8986\ : Span4Mux_h
    port map (
            O => \N__45425\,
            I => \N__45417\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__45422\,
            I => data_in_frame_16_5
        );

    \I__8984\ : Odrv4
    port map (
            O => \N__45417\,
            I => data_in_frame_16_5
        );

    \I__8983\ : InMux
    port map (
            O => \N__45412\,
            I => \N__45409\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__45409\,
            I => \N__45405\
        );

    \I__8981\ : InMux
    port map (
            O => \N__45408\,
            I => \N__45402\
        );

    \I__8980\ : Span4Mux_v
    port map (
            O => \N__45405\,
            I => \N__45399\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__45402\,
            I => data_in_frame_19_0
        );

    \I__8978\ : Odrv4
    port map (
            O => \N__45399\,
            I => data_in_frame_19_0
        );

    \I__8977\ : CascadeMux
    port map (
            O => \N__45394\,
            I => \c0.n9_adj_3430_cascade_\
        );

    \I__8976\ : InMux
    port map (
            O => \N__45391\,
            I => \N__45385\
        );

    \I__8975\ : InMux
    port map (
            O => \N__45390\,
            I => \N__45385\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__45385\,
            I => \N__45382\
        );

    \I__8973\ : Span4Mux_v
    port map (
            O => \N__45382\,
            I => \N__45379\
        );

    \I__8972\ : Odrv4
    port map (
            O => \N__45379\,
            I => \c0.n10_adj_3445\
        );

    \I__8971\ : InMux
    port map (
            O => \N__45376\,
            I => \N__45373\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__45373\,
            I => \c0.n9_adj_3430\
        );

    \I__8969\ : CascadeMux
    port map (
            O => \N__45370\,
            I => \N__45367\
        );

    \I__8968\ : InMux
    port map (
            O => \N__45367\,
            I => \N__45361\
        );

    \I__8967\ : InMux
    port map (
            O => \N__45366\,
            I => \N__45361\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__45361\,
            I => \c0.n14_adj_3421\
        );

    \I__8965\ : CascadeMux
    port map (
            O => \N__45358\,
            I => \c0.n18433_cascade_\
        );

    \I__8964\ : InMux
    port map (
            O => \N__45355\,
            I => \N__45352\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__45352\,
            I => \N__45349\
        );

    \I__8962\ : Odrv4
    port map (
            O => \N__45349\,
            I => \c0.n19511\
        );

    \I__8961\ : InMux
    port map (
            O => \N__45346\,
            I => \N__45340\
        );

    \I__8960\ : InMux
    port map (
            O => \N__45345\,
            I => \N__45340\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__45340\,
            I => \N__45335\
        );

    \I__8958\ : InMux
    port map (
            O => \N__45339\,
            I => \N__45329\
        );

    \I__8957\ : InMux
    port map (
            O => \N__45338\,
            I => \N__45329\
        );

    \I__8956\ : Span4Mux_h
    port map (
            O => \N__45335\,
            I => \N__45326\
        );

    \I__8955\ : InMux
    port map (
            O => \N__45334\,
            I => \N__45323\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__45329\,
            I => \c0.n49\
        );

    \I__8953\ : Odrv4
    port map (
            O => \N__45326\,
            I => \c0.n49\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__45323\,
            I => \c0.n49\
        );

    \I__8951\ : InMux
    port map (
            O => \N__45316\,
            I => \N__45310\
        );

    \I__8950\ : InMux
    port map (
            O => \N__45315\,
            I => \N__45310\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__45310\,
            I => \N__45307\
        );

    \I__8948\ : Span4Mux_h
    port map (
            O => \N__45307\,
            I => \N__45303\
        );

    \I__8947\ : InMux
    port map (
            O => \N__45306\,
            I => \N__45300\
        );

    \I__8946\ : Span4Mux_h
    port map (
            O => \N__45303\,
            I => \N__45297\
        );

    \I__8945\ : LocalMux
    port map (
            O => \N__45300\,
            I => \N__45294\
        );

    \I__8944\ : Span4Mux_h
    port map (
            O => \N__45297\,
            I => \N__45291\
        );

    \I__8943\ : Span4Mux_h
    port map (
            O => \N__45294\,
            I => \N__45287\
        );

    \I__8942\ : Sp12to4
    port map (
            O => \N__45291\,
            I => \N__45284\
        );

    \I__8941\ : InMux
    port map (
            O => \N__45290\,
            I => \N__45281\
        );

    \I__8940\ : Odrv4
    port map (
            O => \N__45287\,
            I => \c0.n48_adj_3409\
        );

    \I__8939\ : Odrv12
    port map (
            O => \N__45284\,
            I => \c0.n48_adj_3409\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__45281\,
            I => \c0.n48_adj_3409\
        );

    \I__8937\ : CascadeMux
    port map (
            O => \N__45274\,
            I => \c0.n22_adj_3287_cascade_\
        );

    \I__8936\ : InMux
    port map (
            O => \N__45271\,
            I => \N__45267\
        );

    \I__8935\ : InMux
    port map (
            O => \N__45270\,
            I => \N__45264\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__45267\,
            I => \N__45259\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__45264\,
            I => \N__45259\
        );

    \I__8932\ : Span4Mux_v
    port map (
            O => \N__45259\,
            I => \N__45256\
        );

    \I__8931\ : Odrv4
    port map (
            O => \N__45256\,
            I => \c0.n39_adj_3050\
        );

    \I__8930\ : CascadeMux
    port map (
            O => \N__45253\,
            I => \c0.n20451_cascade_\
        );

    \I__8929\ : InMux
    port map (
            O => \N__45250\,
            I => \N__45247\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__45247\,
            I => \N__45244\
        );

    \I__8927\ : Span4Mux_h
    port map (
            O => \N__45244\,
            I => \N__45241\
        );

    \I__8926\ : Odrv4
    port map (
            O => \N__45241\,
            I => \c0.n5_adj_3220\
        );

    \I__8925\ : InMux
    port map (
            O => \N__45238\,
            I => \N__45235\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__45235\,
            I => \N__45231\
        );

    \I__8923\ : InMux
    port map (
            O => \N__45234\,
            I => \N__45228\
        );

    \I__8922\ : Span4Mux_v
    port map (
            O => \N__45231\,
            I => \N__45225\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__45228\,
            I => data_in_frame_18_1
        );

    \I__8920\ : Odrv4
    port map (
            O => \N__45225\,
            I => data_in_frame_18_1
        );

    \I__8919\ : CascadeMux
    port map (
            O => \N__45220\,
            I => \c0.n27_adj_3529_cascade_\
        );

    \I__8918\ : CascadeMux
    port map (
            O => \N__45217\,
            I => \c0.n32_adj_3530_cascade_\
        );

    \I__8917\ : CascadeMux
    port map (
            O => \N__45214\,
            I => \c0.n19244_cascade_\
        );

    \I__8916\ : InMux
    port map (
            O => \N__45211\,
            I => \N__45208\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__45208\,
            I => \N__45205\
        );

    \I__8914\ : Span4Mux_h
    port map (
            O => \N__45205\,
            I => \N__45202\
        );

    \I__8913\ : Odrv4
    port map (
            O => \N__45202\,
            I => \c0.n85_adj_3074\
        );

    \I__8912\ : CascadeMux
    port map (
            O => \N__45199\,
            I => \c0.n85_adj_3074_cascade_\
        );

    \I__8911\ : InMux
    port map (
            O => \N__45196\,
            I => \N__45193\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__45193\,
            I => \c0.n10_adj_3474\
        );

    \I__8909\ : InMux
    port map (
            O => \N__45190\,
            I => \N__45183\
        );

    \I__8908\ : InMux
    port map (
            O => \N__45189\,
            I => \N__45183\
        );

    \I__8907\ : InMux
    port map (
            O => \N__45188\,
            I => \N__45176\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__45183\,
            I => \N__45173\
        );

    \I__8905\ : InMux
    port map (
            O => \N__45182\,
            I => \N__45170\
        );

    \I__8904\ : InMux
    port map (
            O => \N__45181\,
            I => \N__45163\
        );

    \I__8903\ : InMux
    port map (
            O => \N__45180\,
            I => \N__45163\
        );

    \I__8902\ : InMux
    port map (
            O => \N__45179\,
            I => \N__45163\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__45176\,
            I => \c0.n20801\
        );

    \I__8900\ : Odrv4
    port map (
            O => \N__45173\,
            I => \c0.n20801\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__45170\,
            I => \c0.n20801\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__45163\,
            I => \c0.n20801\
        );

    \I__8897\ : InMux
    port map (
            O => \N__45154\,
            I => \N__45151\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__45151\,
            I => \N__45148\
        );

    \I__8895\ : Span4Mux_v
    port map (
            O => \N__45148\,
            I => \N__45145\
        );

    \I__8894\ : Odrv4
    port map (
            O => \N__45145\,
            I => \c0.n12_adj_3477\
        );

    \I__8893\ : InMux
    port map (
            O => \N__45142\,
            I => \N__45138\
        );

    \I__8892\ : InMux
    port map (
            O => \N__45141\,
            I => \N__45134\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__45138\,
            I => \N__45131\
        );

    \I__8890\ : InMux
    port map (
            O => \N__45137\,
            I => \N__45128\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__45134\,
            I => \N__45124\
        );

    \I__8888\ : Span4Mux_v
    port map (
            O => \N__45131\,
            I => \N__45121\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__45128\,
            I => \N__45118\
        );

    \I__8886\ : InMux
    port map (
            O => \N__45127\,
            I => \N__45115\
        );

    \I__8885\ : Span12Mux_v
    port map (
            O => \N__45124\,
            I => \N__45112\
        );

    \I__8884\ : Span4Mux_h
    port map (
            O => \N__45121\,
            I => \N__45107\
        );

    \I__8883\ : Span4Mux_v
    port map (
            O => \N__45118\,
            I => \N__45107\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__45115\,
            I => \c0.data_in_frame_14_4\
        );

    \I__8881\ : Odrv12
    port map (
            O => \N__45112\,
            I => \c0.data_in_frame_14_4\
        );

    \I__8880\ : Odrv4
    port map (
            O => \N__45107\,
            I => \c0.data_in_frame_14_4\
        );

    \I__8879\ : CascadeMux
    port map (
            O => \N__45100\,
            I => \c0.n21110_cascade_\
        );

    \I__8878\ : InMux
    port map (
            O => \N__45097\,
            I => \N__45094\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__45094\,
            I => \N__45090\
        );

    \I__8876\ : InMux
    port map (
            O => \N__45093\,
            I => \N__45087\
        );

    \I__8875\ : Span4Mux_v
    port map (
            O => \N__45090\,
            I => \N__45084\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__45087\,
            I => \N__45081\
        );

    \I__8873\ : Span4Mux_v
    port map (
            O => \N__45084\,
            I => \N__45078\
        );

    \I__8872\ : Span4Mux_v
    port map (
            O => \N__45081\,
            I => \N__45075\
        );

    \I__8871\ : Odrv4
    port map (
            O => \N__45078\,
            I => \c0.n20246\
        );

    \I__8870\ : Odrv4
    port map (
            O => \N__45075\,
            I => \c0.n20246\
        );

    \I__8869\ : CascadeMux
    port map (
            O => \N__45070\,
            I => \N__45066\
        );

    \I__8868\ : CascadeMux
    port map (
            O => \N__45069\,
            I => \N__45063\
        );

    \I__8867\ : InMux
    port map (
            O => \N__45066\,
            I => \N__45060\
        );

    \I__8866\ : InMux
    port map (
            O => \N__45063\,
            I => \N__45057\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__45060\,
            I => \c0.data_in_frame_14_3\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__45057\,
            I => \c0.data_in_frame_14_3\
        );

    \I__8863\ : InMux
    port map (
            O => \N__45052\,
            I => \N__45048\
        );

    \I__8862\ : CascadeMux
    port map (
            O => \N__45051\,
            I => \N__45045\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__45048\,
            I => \N__45042\
        );

    \I__8860\ : InMux
    port map (
            O => \N__45045\,
            I => \N__45039\
        );

    \I__8859\ : Span4Mux_h
    port map (
            O => \N__45042\,
            I => \N__45035\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__45039\,
            I => \N__45032\
        );

    \I__8857\ : InMux
    port map (
            O => \N__45038\,
            I => \N__45029\
        );

    \I__8856\ : Odrv4
    port map (
            O => \N__45035\,
            I => \c0.n67_adj_3063\
        );

    \I__8855\ : Odrv12
    port map (
            O => \N__45032\,
            I => \c0.n67_adj_3063\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__45029\,
            I => \c0.n67_adj_3063\
        );

    \I__8853\ : CascadeMux
    port map (
            O => \N__45022\,
            I => \N__45017\
        );

    \I__8852\ : InMux
    port map (
            O => \N__45021\,
            I => \N__45009\
        );

    \I__8851\ : InMux
    port map (
            O => \N__45020\,
            I => \N__45009\
        );

    \I__8850\ : InMux
    port map (
            O => \N__45017\,
            I => \N__45006\
        );

    \I__8849\ : InMux
    port map (
            O => \N__45016\,
            I => \N__44999\
        );

    \I__8848\ : InMux
    port map (
            O => \N__45015\,
            I => \N__44999\
        );

    \I__8847\ : InMux
    port map (
            O => \N__45014\,
            I => \N__44999\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__45009\,
            I => \N__44996\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__45006\,
            I => \N__44991\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__44999\,
            I => \N__44991\
        );

    \I__8843\ : Odrv12
    port map (
            O => \N__44996\,
            I => \c0.n20490\
        );

    \I__8842\ : Odrv4
    port map (
            O => \N__44991\,
            I => \c0.n20490\
        );

    \I__8841\ : InMux
    port map (
            O => \N__44986\,
            I => \N__44980\
        );

    \I__8840\ : InMux
    port map (
            O => \N__44985\,
            I => \N__44980\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__44980\,
            I => \N__44976\
        );

    \I__8838\ : InMux
    port map (
            O => \N__44979\,
            I => \N__44973\
        );

    \I__8837\ : Span4Mux_v
    port map (
            O => \N__44976\,
            I => \N__44964\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__44973\,
            I => \N__44964\
        );

    \I__8835\ : InMux
    port map (
            O => \N__44972\,
            I => \N__44957\
        );

    \I__8834\ : InMux
    port map (
            O => \N__44971\,
            I => \N__44957\
        );

    \I__8833\ : InMux
    port map (
            O => \N__44970\,
            I => \N__44957\
        );

    \I__8832\ : InMux
    port map (
            O => \N__44969\,
            I => \N__44954\
        );

    \I__8831\ : Odrv4
    port map (
            O => \N__44964\,
            I => \c0.n19433\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__44957\,
            I => \c0.n19433\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__44954\,
            I => \c0.n19433\
        );

    \I__8828\ : CascadeMux
    port map (
            O => \N__44947\,
            I => \N__44941\
        );

    \I__8827\ : InMux
    port map (
            O => \N__44946\,
            I => \N__44938\
        );

    \I__8826\ : InMux
    port map (
            O => \N__44945\,
            I => \N__44935\
        );

    \I__8825\ : InMux
    port map (
            O => \N__44944\,
            I => \N__44932\
        );

    \I__8824\ : InMux
    port map (
            O => \N__44941\,
            I => \N__44929\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__44938\,
            I => \c0.n42_adj_3064\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__44935\,
            I => \c0.n42_adj_3064\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__44932\,
            I => \c0.n42_adj_3064\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__44929\,
            I => \c0.n42_adj_3064\
        );

    \I__8819\ : InMux
    port map (
            O => \N__44920\,
            I => \N__44917\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__44917\,
            I => \N__44914\
        );

    \I__8817\ : Span4Mux_v
    port map (
            O => \N__44914\,
            I => \N__44911\
        );

    \I__8816\ : Odrv4
    port map (
            O => \N__44911\,
            I => \c0.n12_adj_3518\
        );

    \I__8815\ : CascadeMux
    port map (
            O => \N__44908\,
            I => \c0.n12_adj_3517_cascade_\
        );

    \I__8814\ : CascadeMux
    port map (
            O => \N__44905\,
            I => \N__44901\
        );

    \I__8813\ : CascadeMux
    port map (
            O => \N__44904\,
            I => \N__44898\
        );

    \I__8812\ : InMux
    port map (
            O => \N__44901\,
            I => \N__44894\
        );

    \I__8811\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44889\
        );

    \I__8810\ : InMux
    port map (
            O => \N__44897\,
            I => \N__44886\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__44894\,
            I => \N__44883\
        );

    \I__8808\ : InMux
    port map (
            O => \N__44893\,
            I => \N__44880\
        );

    \I__8807\ : InMux
    port map (
            O => \N__44892\,
            I => \N__44877\
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__44889\,
            I => \N__44874\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__44886\,
            I => \N__44871\
        );

    \I__8804\ : Span4Mux_v
    port map (
            O => \N__44883\,
            I => \N__44868\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__44880\,
            I => \N__44865\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__44877\,
            I => \N__44860\
        );

    \I__8801\ : Span4Mux_v
    port map (
            O => \N__44874\,
            I => \N__44860\
        );

    \I__8800\ : Span4Mux_v
    port map (
            O => \N__44871\,
            I => \N__44855\
        );

    \I__8799\ : Span4Mux_h
    port map (
            O => \N__44868\,
            I => \N__44855\
        );

    \I__8798\ : Odrv4
    port map (
            O => \N__44865\,
            I => data_in_frame_18_5
        );

    \I__8797\ : Odrv4
    port map (
            O => \N__44860\,
            I => data_in_frame_18_5
        );

    \I__8796\ : Odrv4
    port map (
            O => \N__44855\,
            I => data_in_frame_18_5
        );

    \I__8795\ : InMux
    port map (
            O => \N__44848\,
            I => \N__44845\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__44845\,
            I => \N__44842\
        );

    \I__8793\ : Odrv4
    port map (
            O => \N__44842\,
            I => \c0.n21_adj_3337\
        );

    \I__8792\ : CascadeMux
    port map (
            O => \N__44839\,
            I => \N__44836\
        );

    \I__8791\ : InMux
    port map (
            O => \N__44836\,
            I => \N__44833\
        );

    \I__8790\ : LocalMux
    port map (
            O => \N__44833\,
            I => \N__44830\
        );

    \I__8789\ : Odrv12
    port map (
            O => \N__44830\,
            I => \c0.n20_adj_3487\
        );

    \I__8788\ : InMux
    port map (
            O => \N__44827\,
            I => \N__44824\
        );

    \I__8787\ : LocalMux
    port map (
            O => \N__44824\,
            I => \N__44821\
        );

    \I__8786\ : Odrv4
    port map (
            O => \N__44821\,
            I => \c0.n18_adj_3369\
        );

    \I__8785\ : CascadeMux
    port map (
            O => \N__44818\,
            I => \c0.n19477_cascade_\
        );

    \I__8784\ : CascadeMux
    port map (
            O => \N__44815\,
            I => \c0.n12_adj_3348_cascade_\
        );

    \I__8783\ : CascadeMux
    port map (
            O => \N__44812\,
            I => \c0.n21045_cascade_\
        );

    \I__8782\ : InMux
    port map (
            O => \N__44809\,
            I => \N__44806\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__44806\,
            I => \N__44801\
        );

    \I__8780\ : InMux
    port map (
            O => \N__44805\,
            I => \N__44798\
        );

    \I__8779\ : InMux
    port map (
            O => \N__44804\,
            I => \N__44795\
        );

    \I__8778\ : Odrv4
    port map (
            O => \N__44801\,
            I => \c0.n27_adj_3118\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__44798\,
            I => \c0.n27_adj_3118\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__44795\,
            I => \c0.n27_adj_3118\
        );

    \I__8775\ : InMux
    port map (
            O => \N__44788\,
            I => \N__44785\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__44785\,
            I => \N__44782\
        );

    \I__8773\ : Span4Mux_v
    port map (
            O => \N__44782\,
            I => \N__44779\
        );

    \I__8772\ : Span4Mux_h
    port map (
            O => \N__44779\,
            I => \N__44776\
        );

    \I__8771\ : Span4Mux_v
    port map (
            O => \N__44776\,
            I => \N__44772\
        );

    \I__8770\ : InMux
    port map (
            O => \N__44775\,
            I => \N__44769\
        );

    \I__8769\ : Odrv4
    port map (
            O => \N__44772\,
            I => \c0.n19_adj_3303\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__44769\,
            I => \c0.n19_adj_3303\
        );

    \I__8767\ : InMux
    port map (
            O => \N__44764\,
            I => \N__44761\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__44761\,
            I => \N__44758\
        );

    \I__8765\ : Span12Mux_v
    port map (
            O => \N__44758\,
            I => \N__44755\
        );

    \I__8764\ : Odrv12
    port map (
            O => \N__44755\,
            I => \c0.n12\
        );

    \I__8763\ : InMux
    port map (
            O => \N__44752\,
            I => \N__44749\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__44749\,
            I => \N__44746\
        );

    \I__8761\ : Odrv4
    port map (
            O => \N__44746\,
            I => \c0.n44_adj_3117\
        );

    \I__8760\ : InMux
    port map (
            O => \N__44743\,
            I => \N__44740\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__44740\,
            I => \c0.n43_adj_3116\
        );

    \I__8758\ : CascadeMux
    port map (
            O => \N__44737\,
            I => \c0.n27_adj_3118_cascade_\
        );

    \I__8757\ : InMux
    port map (
            O => \N__44734\,
            I => \N__44731\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__44731\,
            I => \N__44727\
        );

    \I__8755\ : InMux
    port map (
            O => \N__44730\,
            I => \N__44724\
        );

    \I__8754\ : Odrv4
    port map (
            O => \N__44727\,
            I => \c0.n20052\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__44724\,
            I => \c0.n20052\
        );

    \I__8752\ : InMux
    port map (
            O => \N__44719\,
            I => \N__44713\
        );

    \I__8751\ : InMux
    port map (
            O => \N__44718\,
            I => \N__44707\
        );

    \I__8750\ : InMux
    port map (
            O => \N__44717\,
            I => \N__44707\
        );

    \I__8749\ : InMux
    port map (
            O => \N__44716\,
            I => \N__44704\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__44713\,
            I => \N__44701\
        );

    \I__8747\ : CascadeMux
    port map (
            O => \N__44712\,
            I => \N__44698\
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__44707\,
            I => \N__44693\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__44704\,
            I => \N__44693\
        );

    \I__8744\ : Span4Mux_v
    port map (
            O => \N__44701\,
            I => \N__44690\
        );

    \I__8743\ : InMux
    port map (
            O => \N__44698\,
            I => \N__44687\
        );

    \I__8742\ : Span4Mux_v
    port map (
            O => \N__44693\,
            I => \N__44684\
        );

    \I__8741\ : Span4Mux_v
    port map (
            O => \N__44690\,
            I => \N__44681\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__44687\,
            I => \N__44676\
        );

    \I__8739\ : Span4Mux_v
    port map (
            O => \N__44684\,
            I => \N__44676\
        );

    \I__8738\ : Odrv4
    port map (
            O => \N__44681\,
            I => \c0.data_in_frame_14_5\
        );

    \I__8737\ : Odrv4
    port map (
            O => \N__44676\,
            I => \c0.data_in_frame_14_5\
        );

    \I__8736\ : InMux
    port map (
            O => \N__44671\,
            I => \N__44668\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__44668\,
            I => \N__44665\
        );

    \I__8734\ : Odrv12
    port map (
            O => \N__44665\,
            I => \c0.n11_adj_3340\
        );

    \I__8733\ : CascadeMux
    port map (
            O => \N__44662\,
            I => \c0.n19916_cascade_\
        );

    \I__8732\ : CascadeMux
    port map (
            O => \N__44659\,
            I => \N__44655\
        );

    \I__8731\ : InMux
    port map (
            O => \N__44658\,
            I => \N__44651\
        );

    \I__8730\ : InMux
    port map (
            O => \N__44655\,
            I => \N__44646\
        );

    \I__8729\ : InMux
    port map (
            O => \N__44654\,
            I => \N__44646\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__44651\,
            I => \c0.n22_adj_3356\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__44646\,
            I => \c0.n22_adj_3356\
        );

    \I__8726\ : InMux
    port map (
            O => \N__44641\,
            I => \N__44638\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__44638\,
            I => \c0.n22_adj_3022\
        );

    \I__8724\ : CascadeMux
    port map (
            O => \N__44635\,
            I => \N__44628\
        );

    \I__8723\ : CascadeMux
    port map (
            O => \N__44634\,
            I => \N__44625\
        );

    \I__8722\ : InMux
    port map (
            O => \N__44633\,
            I => \N__44619\
        );

    \I__8721\ : InMux
    port map (
            O => \N__44632\,
            I => \N__44619\
        );

    \I__8720\ : InMux
    port map (
            O => \N__44631\,
            I => \N__44616\
        );

    \I__8719\ : InMux
    port map (
            O => \N__44628\,
            I => \N__44613\
        );

    \I__8718\ : InMux
    port map (
            O => \N__44625\,
            I => \N__44610\
        );

    \I__8717\ : CascadeMux
    port map (
            O => \N__44624\,
            I => \N__44607\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__44619\,
            I => \N__44602\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__44616\,
            I => \N__44602\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__44613\,
            I => \N__44597\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__44610\,
            I => \N__44597\
        );

    \I__8712\ : InMux
    port map (
            O => \N__44607\,
            I => \N__44594\
        );

    \I__8711\ : Span4Mux_v
    port map (
            O => \N__44602\,
            I => \N__44589\
        );

    \I__8710\ : Span4Mux_h
    port map (
            O => \N__44597\,
            I => \N__44589\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__44594\,
            I => \c0.data_in_frame_12_4\
        );

    \I__8708\ : Odrv4
    port map (
            O => \N__44589\,
            I => \c0.data_in_frame_12_4\
        );

    \I__8707\ : InMux
    port map (
            O => \N__44584\,
            I => \N__44581\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__44581\,
            I => \N__44578\
        );

    \I__8705\ : Span4Mux_v
    port map (
            O => \N__44578\,
            I => \N__44575\
        );

    \I__8704\ : Odrv4
    port map (
            O => \N__44575\,
            I => \c0.n18_adj_3372\
        );

    \I__8703\ : InMux
    port map (
            O => \N__44572\,
            I => \N__44568\
        );

    \I__8702\ : CascadeMux
    port map (
            O => \N__44571\,
            I => \N__44565\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__44568\,
            I => \N__44562\
        );

    \I__8700\ : InMux
    port map (
            O => \N__44565\,
            I => \N__44559\
        );

    \I__8699\ : Odrv4
    port map (
            O => \N__44562\,
            I => \c0.n88\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__44559\,
            I => \c0.n88\
        );

    \I__8697\ : CascadeMux
    port map (
            O => \N__44554\,
            I => \N__44551\
        );

    \I__8696\ : InMux
    port map (
            O => \N__44551\,
            I => \N__44548\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__44548\,
            I => \c0.n33\
        );

    \I__8694\ : InMux
    port map (
            O => \N__44545\,
            I => \N__44542\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__44542\,
            I => \N__44539\
        );

    \I__8692\ : Span4Mux_h
    port map (
            O => \N__44539\,
            I => \N__44535\
        );

    \I__8691\ : InMux
    port map (
            O => \N__44538\,
            I => \N__44532\
        );

    \I__8690\ : Odrv4
    port map (
            O => \N__44535\,
            I => \c0.n20029\
        );

    \I__8689\ : LocalMux
    port map (
            O => \N__44532\,
            I => \c0.n20029\
        );

    \I__8688\ : InMux
    port map (
            O => \N__44527\,
            I => \N__44524\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__44524\,
            I => \c0.n26_adj_3114\
        );

    \I__8686\ : CascadeMux
    port map (
            O => \N__44521\,
            I => \N__44518\
        );

    \I__8685\ : InMux
    port map (
            O => \N__44518\,
            I => \N__44514\
        );

    \I__8684\ : InMux
    port map (
            O => \N__44517\,
            I => \N__44511\
        );

    \I__8683\ : LocalMux
    port map (
            O => \N__44514\,
            I => \c0.n30\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__44511\,
            I => \c0.n30\
        );

    \I__8681\ : InMux
    port map (
            O => \N__44506\,
            I => \N__44503\
        );

    \I__8680\ : LocalMux
    port map (
            O => \N__44503\,
            I => \N__44500\
        );

    \I__8679\ : Span4Mux_h
    port map (
            O => \N__44500\,
            I => \N__44496\
        );

    \I__8678\ : InMux
    port map (
            O => \N__44499\,
            I => \N__44493\
        );

    \I__8677\ : Odrv4
    port map (
            O => \N__44496\,
            I => \c0.n18422\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__44493\,
            I => \c0.n18422\
        );

    \I__8675\ : CascadeMux
    port map (
            O => \N__44488\,
            I => \c0.n18422_cascade_\
        );

    \I__8674\ : CascadeMux
    port map (
            O => \N__44485\,
            I => \c0.n19433_cascade_\
        );

    \I__8673\ : CascadeMux
    port map (
            O => \N__44482\,
            I => \N__44476\
        );

    \I__8672\ : CascadeMux
    port map (
            O => \N__44481\,
            I => \N__44473\
        );

    \I__8671\ : CascadeMux
    port map (
            O => \N__44480\,
            I => \N__44469\
        );

    \I__8670\ : InMux
    port map (
            O => \N__44479\,
            I => \N__44466\
        );

    \I__8669\ : InMux
    port map (
            O => \N__44476\,
            I => \N__44462\
        );

    \I__8668\ : InMux
    port map (
            O => \N__44473\,
            I => \N__44459\
        );

    \I__8667\ : InMux
    port map (
            O => \N__44472\,
            I => \N__44454\
        );

    \I__8666\ : InMux
    port map (
            O => \N__44469\,
            I => \N__44454\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__44466\,
            I => \N__44451\
        );

    \I__8664\ : InMux
    port map (
            O => \N__44465\,
            I => \N__44448\
        );

    \I__8663\ : LocalMux
    port map (
            O => \N__44462\,
            I => \N__44445\
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__44459\,
            I => \c0.data_in_frame_10_3\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__44454\,
            I => \c0.data_in_frame_10_3\
        );

    \I__8660\ : Odrv4
    port map (
            O => \N__44451\,
            I => \c0.data_in_frame_10_3\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__44448\,
            I => \c0.data_in_frame_10_3\
        );

    \I__8658\ : Odrv4
    port map (
            O => \N__44445\,
            I => \c0.data_in_frame_10_3\
        );

    \I__8657\ : CascadeMux
    port map (
            O => \N__44434\,
            I => \c0.n11891_cascade_\
        );

    \I__8656\ : InMux
    port map (
            O => \N__44431\,
            I => \N__44428\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__44428\,
            I => \c0.n14_adj_3371\
        );

    \I__8654\ : InMux
    port map (
            O => \N__44425\,
            I => \N__44420\
        );

    \I__8653\ : CascadeMux
    port map (
            O => \N__44424\,
            I => \N__44417\
        );

    \I__8652\ : CascadeMux
    port map (
            O => \N__44423\,
            I => \N__44414\
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__44420\,
            I => \N__44410\
        );

    \I__8650\ : InMux
    port map (
            O => \N__44417\,
            I => \N__44403\
        );

    \I__8649\ : InMux
    port map (
            O => \N__44414\,
            I => \N__44403\
        );

    \I__8648\ : InMux
    port map (
            O => \N__44413\,
            I => \N__44403\
        );

    \I__8647\ : Odrv4
    port map (
            O => \N__44410\,
            I => \c0.data_in_frame_3_6\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__44403\,
            I => \c0.data_in_frame_3_6\
        );

    \I__8645\ : CascadeMux
    port map (
            O => \N__44398\,
            I => \c0.n10_adj_3538_cascade_\
        );

    \I__8644\ : CascadeMux
    port map (
            O => \N__44395\,
            I => \N__44390\
        );

    \I__8643\ : InMux
    port map (
            O => \N__44394\,
            I => \N__44387\
        );

    \I__8642\ : CascadeMux
    port map (
            O => \N__44393\,
            I => \N__44384\
        );

    \I__8641\ : InMux
    port map (
            O => \N__44390\,
            I => \N__44379\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__44387\,
            I => \N__44376\
        );

    \I__8639\ : InMux
    port map (
            O => \N__44384\,
            I => \N__44373\
        );

    \I__8638\ : InMux
    port map (
            O => \N__44383\,
            I => \N__44368\
        );

    \I__8637\ : InMux
    port map (
            O => \N__44382\,
            I => \N__44368\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__44379\,
            I => \c0.data_in_frame_2_5\
        );

    \I__8635\ : Odrv12
    port map (
            O => \N__44376\,
            I => \c0.data_in_frame_2_5\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__44373\,
            I => \c0.data_in_frame_2_5\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__44368\,
            I => \c0.data_in_frame_2_5\
        );

    \I__8632\ : CascadeMux
    port map (
            O => \N__44359\,
            I => \c0.n22_adj_3356_cascade_\
        );

    \I__8631\ : InMux
    port map (
            O => \N__44356\,
            I => \N__44352\
        );

    \I__8630\ : InMux
    port map (
            O => \N__44355\,
            I => \N__44349\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__44352\,
            I => \c0.n13_adj_3513\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__44349\,
            I => \c0.n13_adj_3513\
        );

    \I__8627\ : CascadeMux
    port map (
            O => \N__44344\,
            I => \N__44341\
        );

    \I__8626\ : InMux
    port map (
            O => \N__44341\,
            I => \N__44338\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__44338\,
            I => \c0.n23_adj_3021\
        );

    \I__8624\ : CascadeMux
    port map (
            O => \N__44335\,
            I => \c0.n23_adj_3021_cascade_\
        );

    \I__8623\ : CascadeMux
    port map (
            O => \N__44332\,
            I => \c0.n26_adj_3114_cascade_\
        );

    \I__8622\ : InMux
    port map (
            O => \N__44329\,
            I => \N__44323\
        );

    \I__8621\ : InMux
    port map (
            O => \N__44328\,
            I => \N__44323\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__44323\,
            I => \c0.n24_adj_3011\
        );

    \I__8619\ : InMux
    port map (
            O => \N__44320\,
            I => \N__44317\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__44317\,
            I => \N__44314\
        );

    \I__8617\ : Odrv4
    port map (
            O => \N__44314\,
            I => \c0.n22\
        );

    \I__8616\ : InMux
    port map (
            O => \N__44311\,
            I => \N__44305\
        );

    \I__8615\ : InMux
    port map (
            O => \N__44310\,
            I => \N__44305\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__44305\,
            I => \N__44301\
        );

    \I__8613\ : InMux
    port map (
            O => \N__44304\,
            I => \N__44298\
        );

    \I__8612\ : Odrv12
    port map (
            O => \N__44301\,
            I => \c0.n12131\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__44298\,
            I => \c0.n12131\
        );

    \I__8610\ : InMux
    port map (
            O => \N__44293\,
            I => \N__44287\
        );

    \I__8609\ : InMux
    port map (
            O => \N__44292\,
            I => \N__44287\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__44287\,
            I => \c0.n19415\
        );

    \I__8607\ : CascadeMux
    port map (
            O => \N__44284\,
            I => \c0.n19415_cascade_\
        );

    \I__8606\ : InMux
    port map (
            O => \N__44281\,
            I => \N__44275\
        );

    \I__8605\ : InMux
    port map (
            O => \N__44280\,
            I => \N__44275\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__44275\,
            I => \c0.n54_adj_3502\
        );

    \I__8603\ : InMux
    port map (
            O => \N__44272\,
            I => \N__44268\
        );

    \I__8602\ : InMux
    port map (
            O => \N__44271\,
            I => \N__44265\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__44268\,
            I => \c0.n39_adj_3398\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__44265\,
            I => \c0.n39_adj_3398\
        );

    \I__8599\ : InMux
    port map (
            O => \N__44260\,
            I => \N__44257\
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__44257\,
            I => \N__44254\
        );

    \I__8597\ : Span4Mux_h
    port map (
            O => \N__44254\,
            I => \N__44249\
        );

    \I__8596\ : CascadeMux
    port map (
            O => \N__44253\,
            I => \N__44244\
        );

    \I__8595\ : InMux
    port map (
            O => \N__44252\,
            I => \N__44241\
        );

    \I__8594\ : Span4Mux_v
    port map (
            O => \N__44249\,
            I => \N__44237\
        );

    \I__8593\ : InMux
    port map (
            O => \N__44248\,
            I => \N__44234\
        );

    \I__8592\ : InMux
    port map (
            O => \N__44247\,
            I => \N__44230\
        );

    \I__8591\ : InMux
    port map (
            O => \N__44244\,
            I => \N__44227\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__44241\,
            I => \N__44224\
        );

    \I__8589\ : InMux
    port map (
            O => \N__44240\,
            I => \N__44221\
        );

    \I__8588\ : Span4Mux_v
    port map (
            O => \N__44237\,
            I => \N__44217\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__44234\,
            I => \N__44212\
        );

    \I__8586\ : InMux
    port map (
            O => \N__44233\,
            I => \N__44209\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__44230\,
            I => \N__44206\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__44227\,
            I => \N__44199\
        );

    \I__8583\ : Span4Mux_h
    port map (
            O => \N__44224\,
            I => \N__44199\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__44221\,
            I => \N__44199\
        );

    \I__8581\ : InMux
    port map (
            O => \N__44220\,
            I => \N__44196\
        );

    \I__8580\ : Span4Mux_v
    port map (
            O => \N__44217\,
            I => \N__44193\
        );

    \I__8579\ : InMux
    port map (
            O => \N__44216\,
            I => \N__44188\
        );

    \I__8578\ : InMux
    port map (
            O => \N__44215\,
            I => \N__44188\
        );

    \I__8577\ : Span12Mux_h
    port map (
            O => \N__44212\,
            I => \N__44185\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__44209\,
            I => \N__44180\
        );

    \I__8575\ : Span4Mux_v
    port map (
            O => \N__44206\,
            I => \N__44180\
        );

    \I__8574\ : Span4Mux_v
    port map (
            O => \N__44199\,
            I => \N__44177\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__44196\,
            I => \N__44174\
        );

    \I__8572\ : Span4Mux_h
    port map (
            O => \N__44193\,
            I => \N__44171\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__44188\,
            I => \c0.n9_adj_3025\
        );

    \I__8570\ : Odrv12
    port map (
            O => \N__44185\,
            I => \c0.n9_adj_3025\
        );

    \I__8569\ : Odrv4
    port map (
            O => \N__44180\,
            I => \c0.n9_adj_3025\
        );

    \I__8568\ : Odrv4
    port map (
            O => \N__44177\,
            I => \c0.n9_adj_3025\
        );

    \I__8567\ : Odrv12
    port map (
            O => \N__44174\,
            I => \c0.n9_adj_3025\
        );

    \I__8566\ : Odrv4
    port map (
            O => \N__44171\,
            I => \c0.n9_adj_3025\
        );

    \I__8565\ : InMux
    port map (
            O => \N__44158\,
            I => \N__44152\
        );

    \I__8564\ : InMux
    port map (
            O => \N__44157\,
            I => \N__44148\
        );

    \I__8563\ : InMux
    port map (
            O => \N__44156\,
            I => \N__44143\
        );

    \I__8562\ : InMux
    port map (
            O => \N__44155\,
            I => \N__44143\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__44152\,
            I => \N__44140\
        );

    \I__8560\ : InMux
    port map (
            O => \N__44151\,
            I => \N__44137\
        );

    \I__8559\ : LocalMux
    port map (
            O => \N__44148\,
            I => \c0.data_in_frame_2_7\
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__44143\,
            I => \c0.data_in_frame_2_7\
        );

    \I__8557\ : Odrv12
    port map (
            O => \N__44140\,
            I => \c0.data_in_frame_2_7\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__44137\,
            I => \c0.data_in_frame_2_7\
        );

    \I__8555\ : CascadeMux
    port map (
            O => \N__44128\,
            I => \N__44121\
        );

    \I__8554\ : InMux
    port map (
            O => \N__44127\,
            I => \N__44114\
        );

    \I__8553\ : InMux
    port map (
            O => \N__44126\,
            I => \N__44109\
        );

    \I__8552\ : InMux
    port map (
            O => \N__44125\,
            I => \N__44109\
        );

    \I__8551\ : InMux
    port map (
            O => \N__44124\,
            I => \N__44102\
        );

    \I__8550\ : InMux
    port map (
            O => \N__44121\,
            I => \N__44102\
        );

    \I__8549\ : InMux
    port map (
            O => \N__44120\,
            I => \N__44102\
        );

    \I__8548\ : InMux
    port map (
            O => \N__44119\,
            I => \N__44099\
        );

    \I__8547\ : InMux
    port map (
            O => \N__44118\,
            I => \N__44094\
        );

    \I__8546\ : InMux
    port map (
            O => \N__44117\,
            I => \N__44094\
        );

    \I__8545\ : LocalMux
    port map (
            O => \N__44114\,
            I => \N__44091\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__44109\,
            I => \N__44088\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__44102\,
            I => \N__44083\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__44099\,
            I => \N__44083\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__44094\,
            I => \N__44080\
        );

    \I__8540\ : Span4Mux_v
    port map (
            O => \N__44091\,
            I => \N__44077\
        );

    \I__8539\ : Span4Mux_v
    port map (
            O => \N__44088\,
            I => \N__44072\
        );

    \I__8538\ : Span4Mux_v
    port map (
            O => \N__44083\,
            I => \N__44072\
        );

    \I__8537\ : Span4Mux_h
    port map (
            O => \N__44080\,
            I => \N__44069\
        );

    \I__8536\ : Span4Mux_h
    port map (
            O => \N__44077\,
            I => \N__44066\
        );

    \I__8535\ : Span4Mux_h
    port map (
            O => \N__44072\,
            I => \N__44063\
        );

    \I__8534\ : Span4Mux_h
    port map (
            O => \N__44069\,
            I => \N__44058\
        );

    \I__8533\ : Span4Mux_v
    port map (
            O => \N__44066\,
            I => \N__44058\
        );

    \I__8532\ : Odrv4
    port map (
            O => \N__44063\,
            I => \c0.n9_adj_3351\
        );

    \I__8531\ : Odrv4
    port map (
            O => \N__44058\,
            I => \c0.n9_adj_3351\
        );

    \I__8530\ : CascadeMux
    port map (
            O => \N__44053\,
            I => \N__44050\
        );

    \I__8529\ : InMux
    port map (
            O => \N__44050\,
            I => \N__44042\
        );

    \I__8528\ : InMux
    port map (
            O => \N__44049\,
            I => \N__44042\
        );

    \I__8527\ : InMux
    port map (
            O => \N__44048\,
            I => \N__44039\
        );

    \I__8526\ : CascadeMux
    port map (
            O => \N__44047\,
            I => \N__44036\
        );

    \I__8525\ : LocalMux
    port map (
            O => \N__44042\,
            I => \N__44031\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__44039\,
            I => \N__44031\
        );

    \I__8523\ : InMux
    port map (
            O => \N__44036\,
            I => \N__44025\
        );

    \I__8522\ : Span4Mux_h
    port map (
            O => \N__44031\,
            I => \N__44022\
        );

    \I__8521\ : InMux
    port map (
            O => \N__44030\,
            I => \N__44019\
        );

    \I__8520\ : InMux
    port map (
            O => \N__44029\,
            I => \N__44014\
        );

    \I__8519\ : InMux
    port map (
            O => \N__44028\,
            I => \N__44014\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__44025\,
            I => \c0.data_in_frame_4_6\
        );

    \I__8517\ : Odrv4
    port map (
            O => \N__44022\,
            I => \c0.data_in_frame_4_6\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__44019\,
            I => \c0.data_in_frame_4_6\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__44014\,
            I => \c0.data_in_frame_4_6\
        );

    \I__8514\ : InMux
    port map (
            O => \N__44005\,
            I => \N__44002\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__44002\,
            I => \N__43999\
        );

    \I__8512\ : Span4Mux_h
    port map (
            O => \N__43999\,
            I => \N__43996\
        );

    \I__8511\ : Odrv4
    port map (
            O => \N__43996\,
            I => \c0.n11_adj_3507\
        );

    \I__8510\ : CascadeMux
    port map (
            O => \N__43993\,
            I => \N__43990\
        );

    \I__8509\ : InMux
    port map (
            O => \N__43990\,
            I => \N__43987\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__43987\,
            I => \c0.n13_adj_3504\
        );

    \I__8507\ : CascadeMux
    port map (
            O => \N__43984\,
            I => \c0.n12131_cascade_\
        );

    \I__8506\ : InMux
    port map (
            O => \N__43981\,
            I => \N__43978\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__43978\,
            I => \N__43975\
        );

    \I__8504\ : Span4Mux_h
    port map (
            O => \N__43975\,
            I => \N__43969\
        );

    \I__8503\ : InMux
    port map (
            O => \N__43974\,
            I => \N__43966\
        );

    \I__8502\ : InMux
    port map (
            O => \N__43973\,
            I => \N__43961\
        );

    \I__8501\ : InMux
    port map (
            O => \N__43972\,
            I => \N__43961\
        );

    \I__8500\ : Odrv4
    port map (
            O => \N__43969\,
            I => data_in_3_4
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__43966\,
            I => data_in_3_4
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__43961\,
            I => data_in_3_4
        );

    \I__8497\ : InMux
    port map (
            O => \N__43954\,
            I => \N__43950\
        );

    \I__8496\ : InMux
    port map (
            O => \N__43953\,
            I => \N__43947\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__43950\,
            I => data_in_0_0
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__43947\,
            I => data_in_0_0
        );

    \I__8493\ : InMux
    port map (
            O => \N__43942\,
            I => \N__43937\
        );

    \I__8492\ : InMux
    port map (
            O => \N__43941\,
            I => \N__43934\
        );

    \I__8491\ : InMux
    port map (
            O => \N__43940\,
            I => \N__43931\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__43937\,
            I => data_in_1_7
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__43934\,
            I => data_in_1_7
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__43931\,
            I => data_in_1_7
        );

    \I__8487\ : InMux
    port map (
            O => \N__43924\,
            I => \N__43918\
        );

    \I__8486\ : InMux
    port map (
            O => \N__43923\,
            I => \N__43918\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__43918\,
            I => \c0.n10_adj_3231\
        );

    \I__8484\ : InMux
    port map (
            O => \N__43915\,
            I => \N__43912\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__43912\,
            I => \N__43909\
        );

    \I__8482\ : Span4Mux_v
    port map (
            O => \N__43909\,
            I => \N__43903\
        );

    \I__8481\ : InMux
    port map (
            O => \N__43908\,
            I => \N__43898\
        );

    \I__8480\ : InMux
    port map (
            O => \N__43907\,
            I => \N__43898\
        );

    \I__8479\ : InMux
    port map (
            O => \N__43906\,
            I => \N__43895\
        );

    \I__8478\ : Odrv4
    port map (
            O => \N__43903\,
            I => data_in_2_1
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__43898\,
            I => data_in_2_1
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__43895\,
            I => data_in_2_1
        );

    \I__8475\ : InMux
    port map (
            O => \N__43888\,
            I => \N__43883\
        );

    \I__8474\ : InMux
    port map (
            O => \N__43887\,
            I => \N__43880\
        );

    \I__8473\ : InMux
    port map (
            O => \N__43886\,
            I => \N__43877\
        );

    \I__8472\ : LocalMux
    port map (
            O => \N__43883\,
            I => data_in_1_1
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__43880\,
            I => data_in_1_1
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__43877\,
            I => data_in_1_1
        );

    \I__8469\ : InMux
    port map (
            O => \N__43870\,
            I => \N__43866\
        );

    \I__8468\ : InMux
    port map (
            O => \N__43869\,
            I => \N__43863\
        );

    \I__8467\ : LocalMux
    port map (
            O => \N__43866\,
            I => \N__43860\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__43863\,
            I => \N__43856\
        );

    \I__8465\ : Span4Mux_v
    port map (
            O => \N__43860\,
            I => \N__43853\
        );

    \I__8464\ : InMux
    port map (
            O => \N__43859\,
            I => \N__43850\
        );

    \I__8463\ : Span4Mux_h
    port map (
            O => \N__43856\,
            I => \N__43846\
        );

    \I__8462\ : Sp12to4
    port map (
            O => \N__43853\,
            I => \N__43841\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__43850\,
            I => \N__43841\
        );

    \I__8460\ : InMux
    port map (
            O => \N__43849\,
            I => \N__43836\
        );

    \I__8459\ : Sp12to4
    port map (
            O => \N__43846\,
            I => \N__43831\
        );

    \I__8458\ : Span12Mux_h
    port map (
            O => \N__43841\,
            I => \N__43831\
        );

    \I__8457\ : InMux
    port map (
            O => \N__43840\,
            I => \N__43826\
        );

    \I__8456\ : InMux
    port map (
            O => \N__43839\,
            I => \N__43826\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__43836\,
            I => \r_Bit_Index_2\
        );

    \I__8454\ : Odrv12
    port map (
            O => \N__43831\,
            I => \r_Bit_Index_2\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__43826\,
            I => \r_Bit_Index_2\
        );

    \I__8452\ : InMux
    port map (
            O => \N__43819\,
            I => \N__43814\
        );

    \I__8451\ : InMux
    port map (
            O => \N__43818\,
            I => \N__43811\
        );

    \I__8450\ : InMux
    port map (
            O => \N__43817\,
            I => \N__43808\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__43814\,
            I => \N__43805\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__43811\,
            I => \N__43802\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__43808\,
            I => \N__43794\
        );

    \I__8446\ : Span4Mux_h
    port map (
            O => \N__43805\,
            I => \N__43794\
        );

    \I__8445\ : Sp12to4
    port map (
            O => \N__43802\,
            I => \N__43791\
        );

    \I__8444\ : InMux
    port map (
            O => \N__43801\,
            I => \N__43783\
        );

    \I__8443\ : InMux
    port map (
            O => \N__43800\,
            I => \N__43783\
        );

    \I__8442\ : InMux
    port map (
            O => \N__43799\,
            I => \N__43783\
        );

    \I__8441\ : Sp12to4
    port map (
            O => \N__43794\,
            I => \N__43778\
        );

    \I__8440\ : Span12Mux_s7_v
    port map (
            O => \N__43791\,
            I => \N__43778\
        );

    \I__8439\ : InMux
    port map (
            O => \N__43790\,
            I => \N__43775\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__43783\,
            I => \N__43772\
        );

    \I__8437\ : Span12Mux_v
    port map (
            O => \N__43778\,
            I => \N__43769\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__43775\,
            I => \r_Bit_Index_1\
        );

    \I__8435\ : Odrv12
    port map (
            O => \N__43772\,
            I => \r_Bit_Index_1\
        );

    \I__8434\ : Odrv12
    port map (
            O => \N__43769\,
            I => \r_Bit_Index_1\
        );

    \I__8433\ : InMux
    port map (
            O => \N__43762\,
            I => \N__43759\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__43759\,
            I => \N__43756\
        );

    \I__8431\ : Span4Mux_h
    port map (
            O => \N__43756\,
            I => \N__43752\
        );

    \I__8430\ : InMux
    port map (
            O => \N__43755\,
            I => \N__43749\
        );

    \I__8429\ : Odrv4
    port map (
            O => \N__43752\,
            I => n4
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__43749\,
            I => n4
        );

    \I__8427\ : InMux
    port map (
            O => \N__43744\,
            I => \N__43738\
        );

    \I__8426\ : InMux
    port map (
            O => \N__43743\,
            I => \N__43738\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__43738\,
            I => \N__43735\
        );

    \I__8424\ : Span4Mux_h
    port map (
            O => \N__43735\,
            I => \N__43732\
        );

    \I__8423\ : Odrv4
    port map (
            O => \N__43732\,
            I => n4_adj_3579
        );

    \I__8422\ : CascadeMux
    port map (
            O => \N__43729\,
            I => \c0.n15_adj_3297_cascade_\
        );

    \I__8421\ : InMux
    port map (
            O => \N__43726\,
            I => \N__43723\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__43723\,
            I => \c0.n21003\
        );

    \I__8419\ : CascadeMux
    port map (
            O => \N__43720\,
            I => \c0.n21_adj_3300_cascade_\
        );

    \I__8418\ : InMux
    port map (
            O => \N__43717\,
            I => \N__43714\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__43714\,
            I => \c0.n23_adj_3304\
        );

    \I__8416\ : CascadeMux
    port map (
            O => \N__43711\,
            I => \c0.n21247_cascade_\
        );

    \I__8415\ : InMux
    port map (
            O => \N__43708\,
            I => \N__43705\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__43705\,
            I => \c0.n24_adj_3298\
        );

    \I__8413\ : InMux
    port map (
            O => \N__43702\,
            I => \N__43699\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__43699\,
            I => \c0.n14_adj_3354\
        );

    \I__8411\ : InMux
    port map (
            O => \N__43696\,
            I => \N__43690\
        );

    \I__8410\ : InMux
    port map (
            O => \N__43695\,
            I => \N__43690\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__43690\,
            I => \c0.n34\
        );

    \I__8408\ : CascadeMux
    port map (
            O => \N__43687\,
            I => \N__43684\
        );

    \I__8407\ : InMux
    port map (
            O => \N__43684\,
            I => \N__43681\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__43681\,
            I => \c0.n19403\
        );

    \I__8405\ : CascadeMux
    port map (
            O => \N__43678\,
            I => \N__43674\
        );

    \I__8404\ : InMux
    port map (
            O => \N__43677\,
            I => \N__43669\
        );

    \I__8403\ : InMux
    port map (
            O => \N__43674\,
            I => \N__43669\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__43669\,
            I => \N__43665\
        );

    \I__8401\ : InMux
    port map (
            O => \N__43668\,
            I => \N__43662\
        );

    \I__8400\ : Span4Mux_v
    port map (
            O => \N__43665\,
            I => \N__43659\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__43662\,
            I => \c0.data_in_frame_26_6\
        );

    \I__8398\ : Odrv4
    port map (
            O => \N__43659\,
            I => \c0.data_in_frame_26_6\
        );

    \I__8397\ : CascadeMux
    port map (
            O => \N__43654\,
            I => \N__43651\
        );

    \I__8396\ : InMux
    port map (
            O => \N__43651\,
            I => \N__43648\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__43648\,
            I => \c0.n38_adj_3051\
        );

    \I__8394\ : CascadeMux
    port map (
            O => \N__43645\,
            I => \c0.n38_adj_3051_cascade_\
        );

    \I__8393\ : InMux
    port map (
            O => \N__43642\,
            I => \N__43638\
        );

    \I__8392\ : InMux
    port map (
            O => \N__43641\,
            I => \N__43635\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__43638\,
            I => \N__43632\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__43635\,
            I => \c0.n19496\
        );

    \I__8389\ : Odrv4
    port map (
            O => \N__43632\,
            I => \c0.n19496\
        );

    \I__8388\ : InMux
    port map (
            O => \N__43627\,
            I => \N__43624\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__43624\,
            I => \N__43621\
        );

    \I__8386\ : Odrv4
    port map (
            O => \N__43621\,
            I => \c0.n17947\
        );

    \I__8385\ : InMux
    port map (
            O => \N__43618\,
            I => \N__43614\
        );

    \I__8384\ : InMux
    port map (
            O => \N__43617\,
            I => \N__43611\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__43614\,
            I => \N__43606\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__43611\,
            I => \N__43606\
        );

    \I__8381\ : Span4Mux_v
    port map (
            O => \N__43606\,
            I => \N__43603\
        );

    \I__8380\ : Odrv4
    port map (
            O => \N__43603\,
            I => \c0.n60_adj_3065\
        );

    \I__8379\ : InMux
    port map (
            O => \N__43600\,
            I => \N__43597\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__43597\,
            I => \N__43594\
        );

    \I__8377\ : Span4Mux_v
    port map (
            O => \N__43594\,
            I => \N__43591\
        );

    \I__8376\ : Odrv4
    port map (
            O => \N__43591\,
            I => \c0.n64\
        );

    \I__8375\ : CascadeMux
    port map (
            O => \N__43588\,
            I => \c0.n51_cascade_\
        );

    \I__8374\ : InMux
    port map (
            O => \N__43585\,
            I => \N__43579\
        );

    \I__8373\ : InMux
    port map (
            O => \N__43584\,
            I => \N__43579\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__43579\,
            I => \c0.n32_adj_3052\
        );

    \I__8371\ : InMux
    port map (
            O => \N__43576\,
            I => \N__43573\
        );

    \I__8370\ : LocalMux
    port map (
            O => \N__43573\,
            I => \c0.n45_adj_3284\
        );

    \I__8369\ : CascadeMux
    port map (
            O => \N__43570\,
            I => \N__43567\
        );

    \I__8368\ : InMux
    port map (
            O => \N__43567\,
            I => \N__43564\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__43564\,
            I => \c0.n40_adj_3282\
        );

    \I__8366\ : InMux
    port map (
            O => \N__43561\,
            I => \N__43558\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__43558\,
            I => \c0.n20930\
        );

    \I__8364\ : InMux
    port map (
            O => \N__43555\,
            I => \N__43551\
        );

    \I__8363\ : InMux
    port map (
            O => \N__43554\,
            I => \N__43548\
        );

    \I__8362\ : LocalMux
    port map (
            O => \N__43551\,
            I => \N__43544\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__43548\,
            I => \N__43541\
        );

    \I__8360\ : InMux
    port map (
            O => \N__43547\,
            I => \N__43538\
        );

    \I__8359\ : Odrv4
    port map (
            O => \N__43544\,
            I => \c0.n19342\
        );

    \I__8358\ : Odrv12
    port map (
            O => \N__43541\,
            I => \c0.n19342\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__43538\,
            I => \c0.n19342\
        );

    \I__8356\ : CascadeMux
    port map (
            O => \N__43531\,
            I => \c0.n36_adj_3307_cascade_\
        );

    \I__8355\ : InMux
    port map (
            O => \N__43528\,
            I => \N__43525\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__43525\,
            I => \c0.n39_adj_3312\
        );

    \I__8353\ : InMux
    port map (
            O => \N__43522\,
            I => \N__43517\
        );

    \I__8352\ : InMux
    port map (
            O => \N__43521\,
            I => \N__43514\
        );

    \I__8351\ : InMux
    port map (
            O => \N__43520\,
            I => \N__43511\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__43517\,
            I => \N__43506\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__43514\,
            I => \N__43506\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__43511\,
            I => \N__43503\
        );

    \I__8347\ : Span4Mux_v
    port map (
            O => \N__43506\,
            I => \N__43498\
        );

    \I__8346\ : Span4Mux_v
    port map (
            O => \N__43503\,
            I => \N__43498\
        );

    \I__8345\ : Odrv4
    port map (
            O => \N__43498\,
            I => \c0.n29_adj_3148\
        );

    \I__8344\ : InMux
    port map (
            O => \N__43495\,
            I => \N__43492\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__43492\,
            I => \c0.n78_adj_3357\
        );

    \I__8342\ : CascadeMux
    port map (
            O => \N__43489\,
            I => \c0.n75_cascade_\
        );

    \I__8341\ : CascadeMux
    port map (
            O => \N__43486\,
            I => \c0.n93_adj_3373_cascade_\
        );

    \I__8340\ : InMux
    port map (
            O => \N__43483\,
            I => \N__43480\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__43480\,
            I => \N__43477\
        );

    \I__8338\ : Odrv4
    port map (
            O => \N__43477\,
            I => \c0.n96_adj_3419\
        );

    \I__8337\ : CascadeMux
    port map (
            O => \N__43474\,
            I => \c0.n23_adj_3222_cascade_\
        );

    \I__8336\ : InMux
    port map (
            O => \N__43471\,
            I => \N__43468\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__43468\,
            I => \c0.n76\
        );

    \I__8334\ : CascadeMux
    port map (
            O => \N__43465\,
            I => \N__43462\
        );

    \I__8333\ : InMux
    port map (
            O => \N__43462\,
            I => \N__43459\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__43459\,
            I => \N__43456\
        );

    \I__8331\ : Span12Mux_v
    port map (
            O => \N__43456\,
            I => \N__43451\
        );

    \I__8330\ : InMux
    port map (
            O => \N__43455\,
            I => \N__43446\
        );

    \I__8329\ : InMux
    port map (
            O => \N__43454\,
            I => \N__43446\
        );

    \I__8328\ : Odrv12
    port map (
            O => \N__43451\,
            I => encoder0_position_31
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__43446\,
            I => encoder0_position_31
        );

    \I__8326\ : InMux
    port map (
            O => \N__43441\,
            I => \N__43438\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__43438\,
            I => \N__43435\
        );

    \I__8324\ : Span4Mux_h
    port map (
            O => \N__43435\,
            I => \N__43431\
        );

    \I__8323\ : InMux
    port map (
            O => \N__43434\,
            I => \N__43428\
        );

    \I__8322\ : Span4Mux_v
    port map (
            O => \N__43431\,
            I => \N__43425\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__43428\,
            I => data_out_frame_6_7
        );

    \I__8320\ : Odrv4
    port map (
            O => \N__43425\,
            I => data_out_frame_6_7
        );

    \I__8319\ : CascadeMux
    port map (
            O => \N__43420\,
            I => \N__43416\
        );

    \I__8318\ : InMux
    port map (
            O => \N__43419\,
            I => \N__43411\
        );

    \I__8317\ : InMux
    port map (
            O => \N__43416\,
            I => \N__43411\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__43411\,
            I => \N__43407\
        );

    \I__8315\ : InMux
    port map (
            O => \N__43410\,
            I => \N__43404\
        );

    \I__8314\ : Span4Mux_v
    port map (
            O => \N__43407\,
            I => \N__43401\
        );

    \I__8313\ : LocalMux
    port map (
            O => \N__43404\,
            I => data_in_frame_23_2
        );

    \I__8312\ : Odrv4
    port map (
            O => \N__43401\,
            I => data_in_frame_23_2
        );

    \I__8311\ : CascadeMux
    port map (
            O => \N__43396\,
            I => \c0.n13_adj_3405_cascade_\
        );

    \I__8310\ : CascadeMux
    port map (
            O => \N__43393\,
            I => \N__43390\
        );

    \I__8309\ : InMux
    port map (
            O => \N__43390\,
            I => \N__43386\
        );

    \I__8308\ : InMux
    port map (
            O => \N__43389\,
            I => \N__43382\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__43386\,
            I => \N__43379\
        );

    \I__8306\ : InMux
    port map (
            O => \N__43385\,
            I => \N__43376\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__43382\,
            I => \N__43373\
        );

    \I__8304\ : Span4Mux_v
    port map (
            O => \N__43379\,
            I => \N__43370\
        );

    \I__8303\ : LocalMux
    port map (
            O => \N__43376\,
            I => \c0.data_in_frame_27_0\
        );

    \I__8302\ : Odrv4
    port map (
            O => \N__43373\,
            I => \c0.data_in_frame_27_0\
        );

    \I__8301\ : Odrv4
    port map (
            O => \N__43370\,
            I => \c0.data_in_frame_27_0\
        );

    \I__8300\ : CascadeMux
    port map (
            O => \N__43363\,
            I => \c0.n17880_cascade_\
        );

    \I__8299\ : CascadeMux
    port map (
            O => \N__43360\,
            I => \c0.n19342_cascade_\
        );

    \I__8298\ : InMux
    port map (
            O => \N__43357\,
            I => \N__43354\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__43354\,
            I => \c0.n12035\
        );

    \I__8296\ : CascadeMux
    port map (
            O => \N__43351\,
            I => \c0.n19496_cascade_\
        );

    \I__8295\ : InMux
    port map (
            O => \N__43348\,
            I => \N__43345\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__43345\,
            I => \N__43342\
        );

    \I__8293\ : Span4Mux_h
    port map (
            O => \N__43342\,
            I => \N__43339\
        );

    \I__8292\ : Odrv4
    port map (
            O => \N__43339\,
            I => \c0.n15_adj_3395\
        );

    \I__8291\ : CascadeMux
    port map (
            O => \N__43336\,
            I => \c0.n15489_cascade_\
        );

    \I__8290\ : InMux
    port map (
            O => \N__43333\,
            I => \N__43329\
        );

    \I__8289\ : InMux
    port map (
            O => \N__43332\,
            I => \N__43326\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__43329\,
            I => \c0.data_in_frame_15_2\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__43326\,
            I => \c0.data_in_frame_15_2\
        );

    \I__8286\ : CascadeMux
    port map (
            O => \N__43321\,
            I => \c0.n20801_cascade_\
        );

    \I__8285\ : CascadeMux
    port map (
            O => \N__43318\,
            I => \c0.n96_adj_3401_cascade_\
        );

    \I__8284\ : InMux
    port map (
            O => \N__43315\,
            I => \N__43312\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__43312\,
            I => \N__43309\
        );

    \I__8282\ : Span4Mux_v
    port map (
            O => \N__43309\,
            I => \N__43306\
        );

    \I__8281\ : Odrv4
    port map (
            O => \N__43306\,
            I => \c0.n99\
        );

    \I__8280\ : InMux
    port map (
            O => \N__43303\,
            I => \N__43300\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__43300\,
            I => \N__43296\
        );

    \I__8278\ : InMux
    port map (
            O => \N__43299\,
            I => \N__43293\
        );

    \I__8277\ : Span4Mux_v
    port map (
            O => \N__43296\,
            I => \N__43290\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__43293\,
            I => \N__43287\
        );

    \I__8275\ : Odrv4
    port map (
            O => \N__43290\,
            I => \c0.n47_adj_3408\
        );

    \I__8274\ : Odrv4
    port map (
            O => \N__43287\,
            I => \c0.n47_adj_3408\
        );

    \I__8273\ : InMux
    port map (
            O => \N__43282\,
            I => \N__43279\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__43279\,
            I => \N__43270\
        );

    \I__8271\ : InMux
    port map (
            O => \N__43278\,
            I => \N__43267\
        );

    \I__8270\ : InMux
    port map (
            O => \N__43277\,
            I => \N__43262\
        );

    \I__8269\ : InMux
    port map (
            O => \N__43276\,
            I => \N__43262\
        );

    \I__8268\ : InMux
    port map (
            O => \N__43275\,
            I => \N__43257\
        );

    \I__8267\ : InMux
    port map (
            O => \N__43274\,
            I => \N__43257\
        );

    \I__8266\ : InMux
    port map (
            O => \N__43273\,
            I => \N__43254\
        );

    \I__8265\ : Span4Mux_v
    port map (
            O => \N__43270\,
            I => \N__43247\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__43267\,
            I => \N__43247\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__43262\,
            I => \N__43247\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__43257\,
            I => \c0.n18435\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__43254\,
            I => \c0.n18435\
        );

    \I__8260\ : Odrv4
    port map (
            O => \N__43247\,
            I => \c0.n18435\
        );

    \I__8259\ : CascadeMux
    port map (
            O => \N__43240\,
            I => \c0.n42_adj_3064_cascade_\
        );

    \I__8258\ : InMux
    port map (
            O => \N__43237\,
            I => \N__43234\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__43234\,
            I => \N__43231\
        );

    \I__8256\ : Span4Mux_v
    port map (
            O => \N__43231\,
            I => \N__43227\
        );

    \I__8255\ : InMux
    port map (
            O => \N__43230\,
            I => \N__43224\
        );

    \I__8254\ : Span4Mux_v
    port map (
            O => \N__43227\,
            I => \N__43221\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__43224\,
            I => \N__43218\
        );

    \I__8252\ : Odrv4
    port map (
            O => \N__43221\,
            I => \c0.n5_adj_3040\
        );

    \I__8251\ : Odrv4
    port map (
            O => \N__43218\,
            I => \c0.n5_adj_3040\
        );

    \I__8250\ : InMux
    port map (
            O => \N__43213\,
            I => \N__43210\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__43210\,
            I => \N__43207\
        );

    \I__8248\ : Span4Mux_v
    port map (
            O => \N__43207\,
            I => \N__43204\
        );

    \I__8247\ : Span4Mux_v
    port map (
            O => \N__43204\,
            I => \N__43201\
        );

    \I__8246\ : Odrv4
    port map (
            O => \N__43201\,
            I => \c0.n42_adj_3560\
        );

    \I__8245\ : CascadeMux
    port map (
            O => \N__43198\,
            I => \c0.n35_adj_3342_cascade_\
        );

    \I__8244\ : InMux
    port map (
            O => \N__43195\,
            I => \N__43192\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__43192\,
            I => \N__43189\
        );

    \I__8242\ : Span4Mux_h
    port map (
            O => \N__43189\,
            I => \N__43186\
        );

    \I__8241\ : Span4Mux_v
    port map (
            O => \N__43186\,
            I => \N__43183\
        );

    \I__8240\ : Odrv4
    port map (
            O => \N__43183\,
            I => \c0.n39_adj_3339\
        );

    \I__8239\ : InMux
    port map (
            O => \N__43180\,
            I => \N__43176\
        );

    \I__8238\ : CascadeMux
    port map (
            O => \N__43179\,
            I => \N__43173\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__43176\,
            I => \N__43170\
        );

    \I__8236\ : InMux
    port map (
            O => \N__43173\,
            I => \N__43167\
        );

    \I__8235\ : Span4Mux_v
    port map (
            O => \N__43170\,
            I => \N__43164\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__43167\,
            I => \N__43161\
        );

    \I__8233\ : Odrv4
    port map (
            O => \N__43164\,
            I => \c0.n12_adj_3015\
        );

    \I__8232\ : Odrv4
    port map (
            O => \N__43161\,
            I => \c0.n12_adj_3015\
        );

    \I__8231\ : CascadeMux
    port map (
            O => \N__43156\,
            I => \c0.n44_adj_3561_cascade_\
        );

    \I__8230\ : InMux
    port map (
            O => \N__43153\,
            I => \N__43150\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__43150\,
            I => \N__43146\
        );

    \I__8228\ : InMux
    port map (
            O => \N__43149\,
            I => \N__43143\
        );

    \I__8227\ : Span4Mux_h
    port map (
            O => \N__43146\,
            I => \N__43140\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__43143\,
            I => \N__43137\
        );

    \I__8225\ : Span4Mux_v
    port map (
            O => \N__43140\,
            I => \N__43132\
        );

    \I__8224\ : Span4Mux_h
    port map (
            O => \N__43137\,
            I => \N__43132\
        );

    \I__8223\ : Span4Mux_h
    port map (
            O => \N__43132\,
            I => \N__43129\
        );

    \I__8222\ : Odrv4
    port map (
            O => \N__43129\,
            I => \c0.n13_adj_3017\
        );

    \I__8221\ : InMux
    port map (
            O => \N__43126\,
            I => \N__43123\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__43123\,
            I => \c0.n21118\
        );

    \I__8219\ : InMux
    port map (
            O => \N__43120\,
            I => \N__43117\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__43117\,
            I => \N__43113\
        );

    \I__8217\ : InMux
    port map (
            O => \N__43116\,
            I => \N__43110\
        );

    \I__8216\ : Span4Mux_h
    port map (
            O => \N__43113\,
            I => \N__43107\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__43110\,
            I => data_in_frame_18_2
        );

    \I__8214\ : Odrv4
    port map (
            O => \N__43107\,
            I => data_in_frame_18_2
        );

    \I__8213\ : CascadeMux
    port map (
            O => \N__43102\,
            I => \c0.n21118_cascade_\
        );

    \I__8212\ : InMux
    port map (
            O => \N__43099\,
            I => \N__43096\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__43096\,
            I => \c0.n13_adj_3139\
        );

    \I__8210\ : InMux
    port map (
            O => \N__43093\,
            I => \N__43090\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__43090\,
            I => \N__43084\
        );

    \I__8208\ : InMux
    port map (
            O => \N__43089\,
            I => \N__43081\
        );

    \I__8207\ : InMux
    port map (
            O => \N__43088\,
            I => \N__43078\
        );

    \I__8206\ : InMux
    port map (
            O => \N__43087\,
            I => \N__43075\
        );

    \I__8205\ : Sp12to4
    port map (
            O => \N__43084\,
            I => \N__43070\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__43081\,
            I => \N__43070\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__43078\,
            I => \c0.n36_adj_3267\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__43075\,
            I => \c0.n36_adj_3267\
        );

    \I__8201\ : Odrv12
    port map (
            O => \N__43070\,
            I => \c0.n36_adj_3267\
        );

    \I__8200\ : CascadeMux
    port map (
            O => \N__43063\,
            I => \c0.n96_adj_3418_cascade_\
        );

    \I__8199\ : InMux
    port map (
            O => \N__43060\,
            I => \N__43057\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__43057\,
            I => \N__43054\
        );

    \I__8197\ : Span4Mux_v
    port map (
            O => \N__43054\,
            I => \N__43051\
        );

    \I__8196\ : Odrv4
    port map (
            O => \N__43051\,
            I => \c0.n99_adj_3424\
        );

    \I__8195\ : InMux
    port map (
            O => \N__43048\,
            I => \N__43045\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__43045\,
            I => \c0.n77_adj_3415\
        );

    \I__8193\ : CascadeMux
    port map (
            O => \N__43042\,
            I => \N__43038\
        );

    \I__8192\ : CascadeMux
    port map (
            O => \N__43041\,
            I => \N__43035\
        );

    \I__8191\ : InMux
    port map (
            O => \N__43038\,
            I => \N__43027\
        );

    \I__8190\ : InMux
    port map (
            O => \N__43035\,
            I => \N__43027\
        );

    \I__8189\ : InMux
    port map (
            O => \N__43034\,
            I => \N__43027\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__43027\,
            I => \c0.data_in_frame_10_2\
        );

    \I__8187\ : InMux
    port map (
            O => \N__43024\,
            I => \N__43018\
        );

    \I__8186\ : InMux
    port map (
            O => \N__43023\,
            I => \N__43018\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__43018\,
            I => \N__43015\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__43015\,
            I => \c0.n14_adj_3007\
        );

    \I__8183\ : InMux
    port map (
            O => \N__43012\,
            I => \N__43009\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__43009\,
            I => \N__43006\
        );

    \I__8181\ : Span12Mux_v
    port map (
            O => \N__43006\,
            I => \N__43003\
        );

    \I__8180\ : Odrv12
    port map (
            O => \N__43003\,
            I => \c0.n31_adj_3121\
        );

    \I__8179\ : InMux
    port map (
            O => \N__43000\,
            I => \N__42997\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__42997\,
            I => \N__42994\
        );

    \I__8177\ : Odrv12
    port map (
            O => \N__42994\,
            I => \c0.n27\
        );

    \I__8176\ : CascadeMux
    port map (
            O => \N__42991\,
            I => \c0.n28_adj_3120_cascade_\
        );

    \I__8175\ : InMux
    port map (
            O => \N__42988\,
            I => \N__42985\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__42985\,
            I => \N__42982\
        );

    \I__8173\ : Odrv4
    port map (
            O => \N__42982\,
            I => \c0.n33_adj_3122\
        );

    \I__8172\ : CascadeMux
    port map (
            O => \N__42979\,
            I => \c0.n20052_cascade_\
        );

    \I__8171\ : CascadeMux
    port map (
            O => \N__42976\,
            I => \c0.n10_adj_3129_cascade_\
        );

    \I__8170\ : CascadeMux
    port map (
            O => \N__42973\,
            I => \c0.n18400_cascade_\
        );

    \I__8169\ : InMux
    port map (
            O => \N__42970\,
            I => \N__42965\
        );

    \I__8168\ : InMux
    port map (
            O => \N__42969\,
            I => \N__42962\
        );

    \I__8167\ : CascadeMux
    port map (
            O => \N__42968\,
            I => \N__42959\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__42965\,
            I => \N__42956\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__42962\,
            I => \N__42953\
        );

    \I__8164\ : InMux
    port map (
            O => \N__42959\,
            I => \N__42950\
        );

    \I__8163\ : Odrv4
    port map (
            O => \N__42956\,
            I => \c0.n20088\
        );

    \I__8162\ : Odrv4
    port map (
            O => \N__42953\,
            I => \c0.n20088\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__42950\,
            I => \c0.n20088\
        );

    \I__8160\ : CascadeMux
    port map (
            O => \N__42943\,
            I => \c0.n20055_cascade_\
        );

    \I__8159\ : CascadeMux
    port map (
            O => \N__42940\,
            I => \N__42937\
        );

    \I__8158\ : InMux
    port map (
            O => \N__42937\,
            I => \N__42934\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__42934\,
            I => \N__42930\
        );

    \I__8156\ : InMux
    port map (
            O => \N__42933\,
            I => \N__42927\
        );

    \I__8155\ : Span4Mux_h
    port map (
            O => \N__42930\,
            I => \N__42923\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__42927\,
            I => \N__42920\
        );

    \I__8153\ : InMux
    port map (
            O => \N__42926\,
            I => \N__42917\
        );

    \I__8152\ : Span4Mux_v
    port map (
            O => \N__42923\,
            I => \N__42914\
        );

    \I__8151\ : Sp12to4
    port map (
            O => \N__42920\,
            I => \N__42909\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__42917\,
            I => \N__42909\
        );

    \I__8149\ : Odrv4
    port map (
            O => \N__42914\,
            I => \c0.n5_adj_3099\
        );

    \I__8148\ : Odrv12
    port map (
            O => \N__42909\,
            I => \c0.n5_adj_3099\
        );

    \I__8147\ : CascadeMux
    port map (
            O => \N__42904\,
            I => \c0.n37_adj_3110_cascade_\
        );

    \I__8146\ : InMux
    port map (
            O => \N__42901\,
            I => \N__42897\
        );

    \I__8145\ : InMux
    port map (
            O => \N__42900\,
            I => \N__42894\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__42897\,
            I => \c0.n22_adj_3115\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__42894\,
            I => \c0.n22_adj_3115\
        );

    \I__8142\ : CascadeMux
    port map (
            O => \N__42889\,
            I => \c0.n6_adj_3024_cascade_\
        );

    \I__8141\ : CascadeMux
    port map (
            O => \N__42886\,
            I => \c0.n18435_cascade_\
        );

    \I__8140\ : InMux
    port map (
            O => \N__42883\,
            I => \N__42880\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__42880\,
            I => \c0.n28_adj_3519\
        );

    \I__8138\ : CascadeMux
    port map (
            O => \N__42877\,
            I => \c0.n16_adj_3416_cascade_\
        );

    \I__8137\ : InMux
    port map (
            O => \N__42874\,
            I => \N__42871\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__42871\,
            I => \c0.n16_adj_3542\
        );

    \I__8135\ : CascadeMux
    port map (
            O => \N__42868\,
            I => \N__42865\
        );

    \I__8134\ : InMux
    port map (
            O => \N__42865\,
            I => \N__42862\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__42862\,
            I => \N__42858\
        );

    \I__8132\ : InMux
    port map (
            O => \N__42861\,
            I => \N__42855\
        );

    \I__8131\ : Odrv4
    port map (
            O => \N__42858\,
            I => \c0.n5_adj_3528\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__42855\,
            I => \c0.n5_adj_3528\
        );

    \I__8129\ : CascadeMux
    port map (
            O => \N__42850\,
            I => \c0.n78_cascade_\
        );

    \I__8128\ : CascadeMux
    port map (
            O => \N__42847\,
            I => \c0.n30_adj_3119_cascade_\
        );

    \I__8127\ : CascadeMux
    port map (
            O => \N__42844\,
            I => \N__42841\
        );

    \I__8126\ : InMux
    port map (
            O => \N__42841\,
            I => \N__42838\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__42838\,
            I => \N__42835\
        );

    \I__8124\ : Span4Mux_h
    port map (
            O => \N__42835\,
            I => \N__42832\
        );

    \I__8123\ : Span4Mux_v
    port map (
            O => \N__42832\,
            I => \N__42829\
        );

    \I__8122\ : Odrv4
    port map (
            O => \N__42829\,
            I => \c0.n6_adj_3453\
        );

    \I__8121\ : CascadeMux
    port map (
            O => \N__42826\,
            I => \c0.n39_adj_3398_cascade_\
        );

    \I__8120\ : InMux
    port map (
            O => \N__42823\,
            I => \N__42820\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__42820\,
            I => \c0.n13_adj_3526\
        );

    \I__8118\ : InMux
    port map (
            O => \N__42817\,
            I => \N__42813\
        );

    \I__8117\ : InMux
    port map (
            O => \N__42816\,
            I => \N__42810\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__42813\,
            I => \c0.n14_adj_3525\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__42810\,
            I => \c0.n14_adj_3525\
        );

    \I__8114\ : InMux
    port map (
            O => \N__42805\,
            I => \N__42802\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__42802\,
            I => \c0.n15_adj_3543\
        );

    \I__8112\ : CascadeMux
    port map (
            O => \N__42799\,
            I => \c0.n13_adj_3526_cascade_\
        );

    \I__8111\ : CascadeMux
    port map (
            O => \N__42796\,
            I => \N__42793\
        );

    \I__8110\ : InMux
    port map (
            O => \N__42793\,
            I => \N__42787\
        );

    \I__8109\ : InMux
    port map (
            O => \N__42792\,
            I => \N__42787\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__42787\,
            I => \c0.n11_adj_3394\
        );

    \I__8107\ : InMux
    port map (
            O => \N__42784\,
            I => \N__42780\
        );

    \I__8106\ : InMux
    port map (
            O => \N__42783\,
            I => \N__42777\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__42780\,
            I => \c0.n11516\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__42777\,
            I => \c0.n11516\
        );

    \I__8103\ : InMux
    port map (
            O => \N__42772\,
            I => \N__42769\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__42769\,
            I => \c0.n14_adj_3480\
        );

    \I__8101\ : CascadeMux
    port map (
            O => \N__42766\,
            I => \c0.n13_adj_3490_cascade_\
        );

    \I__8100\ : InMux
    port map (
            O => \N__42763\,
            I => \N__42760\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__42760\,
            I => \c0.n13_adj_3546\
        );

    \I__8098\ : InMux
    port map (
            O => \N__42757\,
            I => \N__42753\
        );

    \I__8097\ : CascadeMux
    port map (
            O => \N__42756\,
            I => \N__42750\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__42753\,
            I => \N__42747\
        );

    \I__8095\ : InMux
    port map (
            O => \N__42750\,
            I => \N__42744\
        );

    \I__8094\ : Span4Mux_h
    port map (
            O => \N__42747\,
            I => \N__42741\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__42744\,
            I => \N__42738\
        );

    \I__8092\ : Odrv4
    port map (
            O => \N__42741\,
            I => \c0.n15497\
        );

    \I__8091\ : Odrv4
    port map (
            O => \N__42738\,
            I => \c0.n15497\
        );

    \I__8090\ : InMux
    port map (
            O => \N__42733\,
            I => \N__42730\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__42730\,
            I => \N__42727\
        );

    \I__8088\ : Odrv4
    port map (
            O => \N__42727\,
            I => \c0.n14_adj_3459\
        );

    \I__8087\ : InMux
    port map (
            O => \N__42724\,
            I => \N__42721\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__42721\,
            I => \c0.n10_adj_3068\
        );

    \I__8085\ : CascadeMux
    port map (
            O => \N__42718\,
            I => \N__42714\
        );

    \I__8084\ : InMux
    port map (
            O => \N__42717\,
            I => \N__42709\
        );

    \I__8083\ : InMux
    port map (
            O => \N__42714\,
            I => \N__42709\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__42709\,
            I => \N__42706\
        );

    \I__8081\ : Odrv4
    port map (
            O => \N__42706\,
            I => \c0.n22_adj_3041\
        );

    \I__8080\ : CascadeMux
    port map (
            O => \N__42703\,
            I => \N__42700\
        );

    \I__8079\ : InMux
    port map (
            O => \N__42700\,
            I => \N__42697\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__42697\,
            I => \N__42694\
        );

    \I__8077\ : Odrv4
    port map (
            O => \N__42694\,
            I => \c0.n21079\
        );

    \I__8076\ : InMux
    port map (
            O => \N__42691\,
            I => \N__42687\
        );

    \I__8075\ : InMux
    port map (
            O => \N__42690\,
            I => \N__42684\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__42687\,
            I => \N__42681\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__42684\,
            I => \N__42676\
        );

    \I__8072\ : Span4Mux_h
    port map (
            O => \N__42681\,
            I => \N__42676\
        );

    \I__8071\ : Odrv4
    port map (
            O => \N__42676\,
            I => \c0.n26\
        );

    \I__8070\ : InMux
    port map (
            O => \N__42673\,
            I => \N__42668\
        );

    \I__8069\ : InMux
    port map (
            O => \N__42672\,
            I => \N__42665\
        );

    \I__8068\ : InMux
    port map (
            O => \N__42671\,
            I => \N__42662\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__42668\,
            I => \N__42659\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__42665\,
            I => \N__42654\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__42662\,
            I => \N__42654\
        );

    \I__8064\ : Odrv4
    port map (
            O => \N__42659\,
            I => \c0.n5_adj_3044\
        );

    \I__8063\ : Odrv12
    port map (
            O => \N__42654\,
            I => \c0.n5_adj_3044\
        );

    \I__8062\ : InMux
    port map (
            O => \N__42649\,
            I => \N__42646\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__42646\,
            I => \c0.n25_adj_3045\
        );

    \I__8060\ : CascadeMux
    port map (
            O => \N__42643\,
            I => \c0.n14_adj_3073_cascade_\
        );

    \I__8059\ : InMux
    port map (
            O => \N__42640\,
            I => \N__42637\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__42637\,
            I => \N__42633\
        );

    \I__8057\ : CascadeMux
    port map (
            O => \N__42636\,
            I => \N__42629\
        );

    \I__8056\ : Span4Mux_v
    port map (
            O => \N__42633\,
            I => \N__42625\
        );

    \I__8055\ : InMux
    port map (
            O => \N__42632\,
            I => \N__42622\
        );

    \I__8054\ : InMux
    port map (
            O => \N__42629\,
            I => \N__42619\
        );

    \I__8053\ : InMux
    port map (
            O => \N__42628\,
            I => \N__42616\
        );

    \I__8052\ : Odrv4
    port map (
            O => \N__42625\,
            I => data_in_2_0
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__42622\,
            I => data_in_2_0
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__42619\,
            I => data_in_2_0
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__42616\,
            I => data_in_2_0
        );

    \I__8048\ : InMux
    port map (
            O => \N__42607\,
            I => \N__42599\
        );

    \I__8047\ : InMux
    port map (
            O => \N__42606\,
            I => \N__42599\
        );

    \I__8046\ : InMux
    port map (
            O => \N__42605\,
            I => \N__42594\
        );

    \I__8045\ : InMux
    port map (
            O => \N__42604\,
            I => \N__42594\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__42599\,
            I => data_in_1_0
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__42594\,
            I => data_in_1_0
        );

    \I__8042\ : InMux
    port map (
            O => \N__42589\,
            I => \N__42586\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__42586\,
            I => \N__42583\
        );

    \I__8040\ : Span4Mux_v
    port map (
            O => \N__42583\,
            I => \N__42580\
        );

    \I__8039\ : Odrv4
    port map (
            O => \N__42580\,
            I => \c0.n12_adj_3230\
        );

    \I__8038\ : InMux
    port map (
            O => \N__42577\,
            I => \N__42571\
        );

    \I__8037\ : InMux
    port map (
            O => \N__42576\,
            I => \N__42568\
        );

    \I__8036\ : InMux
    port map (
            O => \N__42575\,
            I => \N__42565\
        );

    \I__8035\ : InMux
    port map (
            O => \N__42574\,
            I => \N__42562\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__42571\,
            I => \N__42555\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__42568\,
            I => \N__42555\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__42565\,
            I => \N__42555\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__42562\,
            I => data_in_2_7
        );

    \I__8030\ : Odrv12
    port map (
            O => \N__42555\,
            I => data_in_2_7
        );

    \I__8029\ : InMux
    port map (
            O => \N__42550\,
            I => \N__42547\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__42547\,
            I => \c0.n11443\
        );

    \I__8027\ : InMux
    port map (
            O => \N__42544\,
            I => \N__42541\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__42541\,
            I => \N__42537\
        );

    \I__8025\ : InMux
    port map (
            O => \N__42540\,
            I => \N__42533\
        );

    \I__8024\ : Span4Mux_h
    port map (
            O => \N__42537\,
            I => \N__42530\
        );

    \I__8023\ : InMux
    port map (
            O => \N__42536\,
            I => \N__42527\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__42533\,
            I => data_in_0_1
        );

    \I__8021\ : Odrv4
    port map (
            O => \N__42530\,
            I => data_in_0_1
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__42527\,
            I => data_in_0_1
        );

    \I__8019\ : CascadeMux
    port map (
            O => \N__42520\,
            I => \N__42513\
        );

    \I__8018\ : CascadeMux
    port map (
            O => \N__42519\,
            I => \N__42509\
        );

    \I__8017\ : InMux
    port map (
            O => \N__42518\,
            I => \N__42501\
        );

    \I__8016\ : InMux
    port map (
            O => \N__42517\,
            I => \N__42498\
        );

    \I__8015\ : InMux
    port map (
            O => \N__42516\,
            I => \N__42488\
        );

    \I__8014\ : InMux
    port map (
            O => \N__42513\,
            I => \N__42488\
        );

    \I__8013\ : InMux
    port map (
            O => \N__42512\,
            I => \N__42488\
        );

    \I__8012\ : InMux
    port map (
            O => \N__42509\,
            I => \N__42483\
        );

    \I__8011\ : InMux
    port map (
            O => \N__42508\,
            I => \N__42483\
        );

    \I__8010\ : CascadeMux
    port map (
            O => \N__42507\,
            I => \N__42480\
        );

    \I__8009\ : InMux
    port map (
            O => \N__42506\,
            I => \N__42476\
        );

    \I__8008\ : InMux
    port map (
            O => \N__42505\,
            I => \N__42473\
        );

    \I__8007\ : InMux
    port map (
            O => \N__42504\,
            I => \N__42470\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__42501\,
            I => \N__42467\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__42498\,
            I => \N__42464\
        );

    \I__8004\ : CascadeMux
    port map (
            O => \N__42497\,
            I => \N__42461\
        );

    \I__8003\ : CascadeMux
    port map (
            O => \N__42496\,
            I => \N__42456\
        );

    \I__8002\ : CascadeMux
    port map (
            O => \N__42495\,
            I => \N__42453\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__42488\,
            I => \N__42448\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__42483\,
            I => \N__42448\
        );

    \I__7999\ : InMux
    port map (
            O => \N__42480\,
            I => \N__42443\
        );

    \I__7998\ : InMux
    port map (
            O => \N__42479\,
            I => \N__42443\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__42476\,
            I => \N__42438\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__42473\,
            I => \N__42438\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__42470\,
            I => \N__42435\
        );

    \I__7994\ : Span4Mux_h
    port map (
            O => \N__42467\,
            I => \N__42430\
        );

    \I__7993\ : Span4Mux_h
    port map (
            O => \N__42464\,
            I => \N__42430\
        );

    \I__7992\ : InMux
    port map (
            O => \N__42461\,
            I => \N__42423\
        );

    \I__7991\ : InMux
    port map (
            O => \N__42460\,
            I => \N__42418\
        );

    \I__7990\ : InMux
    port map (
            O => \N__42459\,
            I => \N__42418\
        );

    \I__7989\ : InMux
    port map (
            O => \N__42456\,
            I => \N__42415\
        );

    \I__7988\ : InMux
    port map (
            O => \N__42453\,
            I => \N__42412\
        );

    \I__7987\ : Span4Mux_v
    port map (
            O => \N__42448\,
            I => \N__42403\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__42443\,
            I => \N__42403\
        );

    \I__7985\ : Span4Mux_v
    port map (
            O => \N__42438\,
            I => \N__42403\
        );

    \I__7984\ : Span4Mux_h
    port map (
            O => \N__42435\,
            I => \N__42403\
        );

    \I__7983\ : Span4Mux_v
    port map (
            O => \N__42430\,
            I => \N__42400\
        );

    \I__7982\ : InMux
    port map (
            O => \N__42429\,
            I => \N__42393\
        );

    \I__7981\ : InMux
    port map (
            O => \N__42428\,
            I => \N__42393\
        );

    \I__7980\ : InMux
    port map (
            O => \N__42427\,
            I => \N__42393\
        );

    \I__7979\ : InMux
    port map (
            O => \N__42426\,
            I => \N__42390\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__42423\,
            I => \N__42385\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__42418\,
            I => \N__42385\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__42415\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__42412\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7974\ : Odrv4
    port map (
            O => \N__42403\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7973\ : Odrv4
    port map (
            O => \N__42400\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__42393\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__42390\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7970\ : Odrv12
    port map (
            O => \N__42385\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7969\ : InMux
    port map (
            O => \N__42370\,
            I => \N__42365\
        );

    \I__7968\ : InMux
    port map (
            O => \N__42369\,
            I => \N__42361\
        );

    \I__7967\ : InMux
    port map (
            O => \N__42368\,
            I => \N__42358\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__42365\,
            I => \N__42355\
        );

    \I__7965\ : InMux
    port map (
            O => \N__42364\,
            I => \N__42352\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__42361\,
            I => \N__42349\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__42358\,
            I => \N__42346\
        );

    \I__7962\ : Span4Mux_v
    port map (
            O => \N__42355\,
            I => \N__42343\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__42352\,
            I => \N__42338\
        );

    \I__7960\ : Span4Mux_h
    port map (
            O => \N__42349\,
            I => \N__42338\
        );

    \I__7959\ : Odrv12
    port map (
            O => \N__42346\,
            I => n4_adj_3596
        );

    \I__7958\ : Odrv4
    port map (
            O => \N__42343\,
            I => n4_adj_3596
        );

    \I__7957\ : Odrv4
    port map (
            O => \N__42338\,
            I => n4_adj_3596
        );

    \I__7956\ : InMux
    port map (
            O => \N__42331\,
            I => \N__42325\
        );

    \I__7955\ : InMux
    port map (
            O => \N__42330\,
            I => \N__42320\
        );

    \I__7954\ : InMux
    port map (
            O => \N__42329\,
            I => \N__42317\
        );

    \I__7953\ : InMux
    port map (
            O => \N__42328\,
            I => \N__42314\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__42325\,
            I => \N__42311\
        );

    \I__7951\ : InMux
    port map (
            O => \N__42324\,
            I => \N__42305\
        );

    \I__7950\ : InMux
    port map (
            O => \N__42323\,
            I => \N__42305\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__42320\,
            I => \N__42302\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__42317\,
            I => \N__42299\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__42314\,
            I => \N__42294\
        );

    \I__7946\ : Span4Mux_h
    port map (
            O => \N__42311\,
            I => \N__42294\
        );

    \I__7945\ : InMux
    port map (
            O => \N__42310\,
            I => \N__42290\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__42305\,
            I => \N__42287\
        );

    \I__7943\ : Span4Mux_h
    port map (
            O => \N__42302\,
            I => \N__42280\
        );

    \I__7942\ : Span4Mux_h
    port map (
            O => \N__42299\,
            I => \N__42280\
        );

    \I__7941\ : Span4Mux_v
    port map (
            O => \N__42294\,
            I => \N__42280\
        );

    \I__7940\ : InMux
    port map (
            O => \N__42293\,
            I => \N__42277\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__42290\,
            I => n11421
        );

    \I__7938\ : Odrv12
    port map (
            O => \N__42287\,
            I => n11421
        );

    \I__7937\ : Odrv4
    port map (
            O => \N__42280\,
            I => n11421
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__42277\,
            I => n11421
        );

    \I__7935\ : InMux
    port map (
            O => \N__42268\,
            I => \N__42262\
        );

    \I__7934\ : InMux
    port map (
            O => \N__42267\,
            I => \N__42259\
        );

    \I__7933\ : InMux
    port map (
            O => \N__42266\,
            I => \N__42256\
        );

    \I__7932\ : InMux
    port map (
            O => \N__42265\,
            I => \N__42253\
        );

    \I__7931\ : LocalMux
    port map (
            O => \N__42262\,
            I => \N__42240\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__42259\,
            I => \N__42240\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__42256\,
            I => \N__42240\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__42253\,
            I => \N__42240\
        );

    \I__7927\ : InMux
    port map (
            O => \N__42252\,
            I => \N__42237\
        );

    \I__7926\ : InMux
    port map (
            O => \N__42251\,
            I => \N__42234\
        );

    \I__7925\ : InMux
    port map (
            O => \N__42250\,
            I => \N__42231\
        );

    \I__7924\ : InMux
    port map (
            O => \N__42249\,
            I => \N__42228\
        );

    \I__7923\ : Span4Mux_v
    port map (
            O => \N__42240\,
            I => \N__42213\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__42237\,
            I => \N__42213\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__42234\,
            I => \N__42213\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__42231\,
            I => \N__42213\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__42228\,
            I => \N__42213\
        );

    \I__7918\ : InMux
    port map (
            O => \N__42227\,
            I => \N__42210\
        );

    \I__7917\ : InMux
    port map (
            O => \N__42226\,
            I => \N__42207\
        );

    \I__7916\ : InMux
    port map (
            O => \N__42225\,
            I => \N__42204\
        );

    \I__7915\ : InMux
    port map (
            O => \N__42224\,
            I => \N__42201\
        );

    \I__7914\ : Span4Mux_v
    port map (
            O => \N__42213\,
            I => \N__42184\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__42210\,
            I => \N__42184\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__42207\,
            I => \N__42184\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__42204\,
            I => \N__42184\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__42201\,
            I => \N__42184\
        );

    \I__7909\ : InMux
    port map (
            O => \N__42200\,
            I => \N__42181\
        );

    \I__7908\ : InMux
    port map (
            O => \N__42199\,
            I => \N__42178\
        );

    \I__7907\ : InMux
    port map (
            O => \N__42198\,
            I => \N__42175\
        );

    \I__7906\ : InMux
    port map (
            O => \N__42197\,
            I => \N__42172\
        );

    \I__7905\ : InMux
    port map (
            O => \N__42196\,
            I => \N__42164\
        );

    \I__7904\ : InMux
    port map (
            O => \N__42195\,
            I => \N__42164\
        );

    \I__7903\ : Span4Mux_v
    port map (
            O => \N__42184\,
            I => \N__42153\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__42181\,
            I => \N__42153\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__42178\,
            I => \N__42153\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__42175\,
            I => \N__42153\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__42172\,
            I => \N__42153\
        );

    \I__7898\ : InMux
    port map (
            O => \N__42171\,
            I => \N__42146\
        );

    \I__7897\ : InMux
    port map (
            O => \N__42170\,
            I => \N__42146\
        );

    \I__7896\ : InMux
    port map (
            O => \N__42169\,
            I => \N__42146\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__42164\,
            I => \N__42133\
        );

    \I__7894\ : Span4Mux_v
    port map (
            O => \N__42153\,
            I => \N__42133\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__42146\,
            I => \N__42133\
        );

    \I__7892\ : InMux
    port map (
            O => \N__42145\,
            I => \N__42128\
        );

    \I__7891\ : InMux
    port map (
            O => \N__42144\,
            I => \N__42122\
        );

    \I__7890\ : InMux
    port map (
            O => \N__42143\,
            I => \N__42118\
        );

    \I__7889\ : InMux
    port map (
            O => \N__42142\,
            I => \N__42115\
        );

    \I__7888\ : InMux
    port map (
            O => \N__42141\,
            I => \N__42112\
        );

    \I__7887\ : InMux
    port map (
            O => \N__42140\,
            I => \N__42109\
        );

    \I__7886\ : Span4Mux_h
    port map (
            O => \N__42133\,
            I => \N__42106\
        );

    \I__7885\ : InMux
    port map (
            O => \N__42132\,
            I => \N__42103\
        );

    \I__7884\ : InMux
    port map (
            O => \N__42131\,
            I => \N__42100\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__42128\,
            I => \N__42097\
        );

    \I__7882\ : InMux
    port map (
            O => \N__42127\,
            I => \N__42094\
        );

    \I__7881\ : InMux
    port map (
            O => \N__42126\,
            I => \N__42091\
        );

    \I__7880\ : InMux
    port map (
            O => \N__42125\,
            I => \N__42088\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__42122\,
            I => \N__42085\
        );

    \I__7878\ : InMux
    port map (
            O => \N__42121\,
            I => \N__42082\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__42118\,
            I => \N__42075\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__42115\,
            I => \N__42075\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__42112\,
            I => \N__42075\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__42109\,
            I => \N__42072\
        );

    \I__7873\ : Sp12to4
    port map (
            O => \N__42106\,
            I => \N__42068\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__42103\,
            I => \N__42065\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__42100\,
            I => \N__42062\
        );

    \I__7870\ : Span4Mux_h
    port map (
            O => \N__42097\,
            I => \N__42057\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__42094\,
            I => \N__42057\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__42091\,
            I => \N__42048\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__42088\,
            I => \N__42048\
        );

    \I__7866\ : Span4Mux_s1_v
    port map (
            O => \N__42085\,
            I => \N__42048\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__42082\,
            I => \N__42048\
        );

    \I__7864\ : Span4Mux_v
    port map (
            O => \N__42075\,
            I => \N__42043\
        );

    \I__7863\ : Span4Mux_v
    port map (
            O => \N__42072\,
            I => \N__42043\
        );

    \I__7862\ : InMux
    port map (
            O => \N__42071\,
            I => \N__42040\
        );

    \I__7861\ : Span12Mux_s7_v
    port map (
            O => \N__42068\,
            I => \N__42037\
        );

    \I__7860\ : Span12Mux_h
    port map (
            O => \N__42065\,
            I => \N__42034\
        );

    \I__7859\ : Span4Mux_h
    port map (
            O => \N__42062\,
            I => \N__42031\
        );

    \I__7858\ : Span4Mux_v
    port map (
            O => \N__42057\,
            I => \N__42026\
        );

    \I__7857\ : Span4Mux_v
    port map (
            O => \N__42048\,
            I => \N__42026\
        );

    \I__7856\ : Span4Mux_h
    port map (
            O => \N__42043\,
            I => \N__42021\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__42040\,
            I => \N__42021\
        );

    \I__7854\ : Span12Mux_v
    port map (
            O => \N__42037\,
            I => \N__42018\
        );

    \I__7853\ : Span12Mux_v
    port map (
            O => \N__42034\,
            I => \N__42015\
        );

    \I__7852\ : Odrv4
    port map (
            O => \N__42031\,
            I => n1295
        );

    \I__7851\ : Odrv4
    port map (
            O => \N__42026\,
            I => n1295
        );

    \I__7850\ : Odrv4
    port map (
            O => \N__42021\,
            I => n1295
        );

    \I__7849\ : Odrv12
    port map (
            O => \N__42018\,
            I => n1295
        );

    \I__7848\ : Odrv12
    port map (
            O => \N__42015\,
            I => n1295
        );

    \I__7847\ : CascadeMux
    port map (
            O => \N__42004\,
            I => \N__41999\
        );

    \I__7846\ : InMux
    port map (
            O => \N__42003\,
            I => \N__41995\
        );

    \I__7845\ : InMux
    port map (
            O => \N__42002\,
            I => \N__41992\
        );

    \I__7844\ : InMux
    port map (
            O => \N__41999\,
            I => \N__41987\
        );

    \I__7843\ : InMux
    port map (
            O => \N__41998\,
            I => \N__41987\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__41995\,
            I => \N__41982\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__41992\,
            I => \N__41982\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__41987\,
            I => \c0.data_in_frame_27_7\
        );

    \I__7839\ : Odrv12
    port map (
            O => \N__41982\,
            I => \c0.data_in_frame_27_7\
        );

    \I__7838\ : InMux
    port map (
            O => \N__41977\,
            I => \N__41974\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__41974\,
            I => \N__41968\
        );

    \I__7836\ : InMux
    port map (
            O => \N__41973\,
            I => \N__41965\
        );

    \I__7835\ : InMux
    port map (
            O => \N__41972\,
            I => \N__41960\
        );

    \I__7834\ : InMux
    port map (
            O => \N__41971\,
            I => \N__41960\
        );

    \I__7833\ : Sp12to4
    port map (
            O => \N__41968\,
            I => \N__41955\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__41965\,
            I => \N__41955\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__41960\,
            I => \c0.data_in_frame_27_6\
        );

    \I__7830\ : Odrv12
    port map (
            O => \N__41955\,
            I => \c0.data_in_frame_27_6\
        );

    \I__7829\ : CascadeMux
    port map (
            O => \N__41950\,
            I => \N__41946\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__41949\,
            I => \N__41943\
        );

    \I__7827\ : InMux
    port map (
            O => \N__41946\,
            I => \N__41939\
        );

    \I__7826\ : InMux
    port map (
            O => \N__41943\,
            I => \N__41934\
        );

    \I__7825\ : InMux
    port map (
            O => \N__41942\,
            I => \N__41934\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__41939\,
            I => \c0.data_in_frame_26_4\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__41934\,
            I => \c0.data_in_frame_26_4\
        );

    \I__7822\ : InMux
    port map (
            O => \N__41929\,
            I => \N__41923\
        );

    \I__7821\ : InMux
    port map (
            O => \N__41928\,
            I => \N__41918\
        );

    \I__7820\ : InMux
    port map (
            O => \N__41927\,
            I => \N__41918\
        );

    \I__7819\ : InMux
    port map (
            O => \N__41926\,
            I => \N__41915\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__41923\,
            I => data_in_2_2
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__41918\,
            I => data_in_2_2
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__41915\,
            I => data_in_2_2
        );

    \I__7815\ : InMux
    port map (
            O => \N__41908\,
            I => \N__41905\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__41905\,
            I => \c0.n10_adj_3238\
        );

    \I__7813\ : InMux
    port map (
            O => \N__41902\,
            I => \N__41899\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__41899\,
            I => \N__41896\
        );

    \I__7811\ : Span4Mux_v
    port map (
            O => \N__41896\,
            I => \N__41892\
        );

    \I__7810\ : InMux
    port map (
            O => \N__41895\,
            I => \N__41889\
        );

    \I__7809\ : Odrv4
    port map (
            O => \N__41892\,
            I => \c0.n110\
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__41889\,
            I => \c0.n110\
        );

    \I__7807\ : InMux
    port map (
            O => \N__41884\,
            I => \N__41881\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__41881\,
            I => \N__41878\
        );

    \I__7805\ : Span4Mux_v
    port map (
            O => \N__41878\,
            I => \N__41872\
        );

    \I__7804\ : InMux
    port map (
            O => \N__41877\,
            I => \N__41869\
        );

    \I__7803\ : InMux
    port map (
            O => \N__41876\,
            I => \N__41866\
        );

    \I__7802\ : InMux
    port map (
            O => \N__41875\,
            I => \N__41863\
        );

    \I__7801\ : Odrv4
    port map (
            O => \N__41872\,
            I => data_in_2_5
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__41869\,
            I => data_in_2_5
        );

    \I__7799\ : LocalMux
    port map (
            O => \N__41866\,
            I => data_in_2_5
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__41863\,
            I => data_in_2_5
        );

    \I__7797\ : InMux
    port map (
            O => \N__41854\,
            I => \N__41848\
        );

    \I__7796\ : InMux
    port map (
            O => \N__41853\,
            I => \N__41845\
        );

    \I__7795\ : InMux
    port map (
            O => \N__41852\,
            I => \N__41840\
        );

    \I__7794\ : InMux
    port map (
            O => \N__41851\,
            I => \N__41840\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__41848\,
            I => data_in_1_5
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__41845\,
            I => data_in_1_5
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__41840\,
            I => data_in_1_5
        );

    \I__7790\ : InMux
    port map (
            O => \N__41833\,
            I => \N__41830\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__41830\,
            I => \N__41826\
        );

    \I__7788\ : CascadeMux
    port map (
            O => \N__41829\,
            I => \N__41823\
        );

    \I__7787\ : Span12Mux_s9_v
    port map (
            O => \N__41826\,
            I => \N__41820\
        );

    \I__7786\ : InMux
    port map (
            O => \N__41823\,
            I => \N__41817\
        );

    \I__7785\ : Span12Mux_h
    port map (
            O => \N__41820\,
            I => \N__41814\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__41817\,
            I => \N__41811\
        );

    \I__7783\ : Span12Mux_v
    port map (
            O => \N__41814\,
            I => \N__41808\
        );

    \I__7782\ : Span4Mux_v
    port map (
            O => \N__41811\,
            I => \N__41805\
        );

    \I__7781\ : Odrv12
    port map (
            O => \N__41808\,
            I => \c0.n160\
        );

    \I__7780\ : Odrv4
    port map (
            O => \N__41805\,
            I => \c0.n160\
        );

    \I__7779\ : InMux
    port map (
            O => \N__41800\,
            I => \N__41794\
        );

    \I__7778\ : InMux
    port map (
            O => \N__41799\,
            I => \N__41794\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__41794\,
            I => \c0.data_in_frame_29_0\
        );

    \I__7776\ : CascadeMux
    port map (
            O => \N__41791\,
            I => \c0.n21117_cascade_\
        );

    \I__7775\ : InMux
    port map (
            O => \N__41788\,
            I => \N__41785\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__41785\,
            I => \c0.n18\
        );

    \I__7773\ : InMux
    port map (
            O => \N__41782\,
            I => \N__41779\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__41779\,
            I => \c0.n5_adj_3142\
        );

    \I__7771\ : CascadeMux
    port map (
            O => \N__41776\,
            I => \c0.n5_adj_3142_cascade_\
        );

    \I__7770\ : CascadeMux
    port map (
            O => \N__41773\,
            I => \c0.n22_adj_3305_cascade_\
        );

    \I__7769\ : CascadeMux
    port map (
            O => \N__41770\,
            I => \c0.n37_adj_3309_cascade_\
        );

    \I__7768\ : CascadeMux
    port map (
            O => \N__41767\,
            I => \c0.n21099_cascade_\
        );

    \I__7767\ : InMux
    port map (
            O => \N__41764\,
            I => \N__41761\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__41761\,
            I => \c0.n18_adj_3314\
        );

    \I__7765\ : CascadeMux
    port map (
            O => \N__41758\,
            I => \c0.n10_adj_3353_cascade_\
        );

    \I__7764\ : InMux
    port map (
            O => \N__41755\,
            I => \N__41752\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__41752\,
            I => \N__41749\
        );

    \I__7762\ : Span12Mux_v
    port map (
            O => \N__41749\,
            I => \N__41746\
        );

    \I__7761\ : Odrv12
    port map (
            O => \N__41746\,
            I => \c0.n21111\
        );

    \I__7760\ : CascadeMux
    port map (
            O => \N__41743\,
            I => \c0.n9_adj_3352_cascade_\
        );

    \I__7759\ : InMux
    port map (
            O => \N__41740\,
            I => \N__41737\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__41737\,
            I => \c0.n21051\
        );

    \I__7757\ : InMux
    port map (
            O => \N__41734\,
            I => \N__41731\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__41731\,
            I => \N__41728\
        );

    \I__7755\ : Span4Mux_v
    port map (
            O => \N__41728\,
            I => \N__41725\
        );

    \I__7754\ : Odrv4
    port map (
            O => \N__41725\,
            I => \c0.n18537\
        );

    \I__7753\ : InMux
    port map (
            O => \N__41722\,
            I => \N__41718\
        );

    \I__7752\ : InMux
    port map (
            O => \N__41721\,
            I => \N__41715\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__41718\,
            I => \c0.n20370\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__41715\,
            I => \c0.n20370\
        );

    \I__7749\ : CascadeMux
    port map (
            O => \N__41710\,
            I => \N__41707\
        );

    \I__7748\ : InMux
    port map (
            O => \N__41707\,
            I => \N__41703\
        );

    \I__7747\ : InMux
    port map (
            O => \N__41706\,
            I => \N__41700\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__41703\,
            I => \c0.data_in_frame_29_7\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__41700\,
            I => \c0.data_in_frame_29_7\
        );

    \I__7744\ : CascadeMux
    port map (
            O => \N__41695\,
            I => \N__41691\
        );

    \I__7743\ : CascadeMux
    port map (
            O => \N__41694\,
            I => \N__41688\
        );

    \I__7742\ : InMux
    port map (
            O => \N__41691\,
            I => \N__41685\
        );

    \I__7741\ : InMux
    port map (
            O => \N__41688\,
            I => \N__41682\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__41685\,
            I => \c0.data_in_frame_29_6\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__41682\,
            I => \c0.data_in_frame_29_6\
        );

    \I__7738\ : CascadeMux
    port map (
            O => \N__41677\,
            I => \c0.n10_adj_3152_cascade_\
        );

    \I__7737\ : InMux
    port map (
            O => \N__41674\,
            I => \N__41671\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__41671\,
            I => \c0.n21117\
        );

    \I__7735\ : CascadeMux
    port map (
            O => \N__41668\,
            I => \c0.n61_cascade_\
        );

    \I__7734\ : InMux
    port map (
            O => \N__41665\,
            I => \N__41662\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__41662\,
            I => \c0.n50\
        );

    \I__7732\ : InMux
    port map (
            O => \N__41659\,
            I => \N__41656\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__41656\,
            I => \c0.n61\
        );

    \I__7730\ : CascadeMux
    port map (
            O => \N__41653\,
            I => \c0.n86_adj_3393_cascade_\
        );

    \I__7729\ : CascadeMux
    port map (
            O => \N__41650\,
            I => \c0.n95_cascade_\
        );

    \I__7728\ : InMux
    port map (
            O => \N__41647\,
            I => \N__41644\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__41644\,
            I => \N__41641\
        );

    \I__7726\ : Span4Mux_v
    port map (
            O => \N__41641\,
            I => \N__41638\
        );

    \I__7725\ : Odrv4
    port map (
            O => \N__41638\,
            I => \c0.n15_adj_3441\
        );

    \I__7724\ : InMux
    port map (
            O => \N__41635\,
            I => \N__41632\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__41632\,
            I => \N__41628\
        );

    \I__7722\ : InMux
    port map (
            O => \N__41631\,
            I => \N__41625\
        );

    \I__7721\ : Span4Mux_v
    port map (
            O => \N__41628\,
            I => \N__41620\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__41625\,
            I => \N__41617\
        );

    \I__7719\ : InMux
    port map (
            O => \N__41624\,
            I => \N__41612\
        );

    \I__7718\ : InMux
    port map (
            O => \N__41623\,
            I => \N__41612\
        );

    \I__7717\ : Odrv4
    port map (
            O => \N__41620\,
            I => data_in_3_7
        );

    \I__7716\ : Odrv4
    port map (
            O => \N__41617\,
            I => data_in_3_7
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__41612\,
            I => data_in_3_7
        );

    \I__7714\ : CascadeMux
    port map (
            O => \N__41605\,
            I => \N__41601\
        );

    \I__7713\ : CascadeMux
    port map (
            O => \N__41604\,
            I => \N__41597\
        );

    \I__7712\ : InMux
    port map (
            O => \N__41601\,
            I => \N__41594\
        );

    \I__7711\ : InMux
    port map (
            O => \N__41600\,
            I => \N__41591\
        );

    \I__7710\ : InMux
    port map (
            O => \N__41597\,
            I => \N__41588\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__41594\,
            I => \N__41585\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__41591\,
            I => data_in_frame_16_6
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__41588\,
            I => data_in_frame_16_6
        );

    \I__7706\ : Odrv12
    port map (
            O => \N__41585\,
            I => data_in_frame_16_6
        );

    \I__7705\ : InMux
    port map (
            O => \N__41578\,
            I => \N__41574\
        );

    \I__7704\ : InMux
    port map (
            O => \N__41577\,
            I => \N__41571\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__41574\,
            I => \c0.data_in_frame_28_4\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__41571\,
            I => \c0.data_in_frame_28_4\
        );

    \I__7701\ : InMux
    port map (
            O => \N__41566\,
            I => \N__41563\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__41563\,
            I => \N__41560\
        );

    \I__7699\ : Span4Mux_h
    port map (
            O => \N__41560\,
            I => \N__41557\
        );

    \I__7698\ : Span4Mux_v
    port map (
            O => \N__41557\,
            I => \N__41554\
        );

    \I__7697\ : Odrv4
    port map (
            O => \N__41554\,
            I => \c0.n20931\
        );

    \I__7696\ : InMux
    port map (
            O => \N__41551\,
            I => \N__41548\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__41548\,
            I => \N__41544\
        );

    \I__7694\ : InMux
    port map (
            O => \N__41547\,
            I => \N__41541\
        );

    \I__7693\ : Span4Mux_v
    port map (
            O => \N__41544\,
            I => \N__41538\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__41541\,
            I => data_in_frame_18_6
        );

    \I__7691\ : Odrv4
    port map (
            O => \N__41538\,
            I => data_in_frame_18_6
        );

    \I__7690\ : InMux
    port map (
            O => \N__41533\,
            I => \N__41530\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__41530\,
            I => \N__41526\
        );

    \I__7688\ : InMux
    port map (
            O => \N__41529\,
            I => \N__41523\
        );

    \I__7687\ : Odrv4
    port map (
            O => \N__41526\,
            I => n4_adj_3595
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__41523\,
            I => n4_adj_3595
        );

    \I__7685\ : InMux
    port map (
            O => \N__41518\,
            I => \N__41515\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__41515\,
            I => \N__41512\
        );

    \I__7683\ : Span4Mux_v
    port map (
            O => \N__41512\,
            I => \N__41509\
        );

    \I__7682\ : Odrv4
    port map (
            O => \N__41509\,
            I => \c0.n14_adj_3434\
        );

    \I__7681\ : InMux
    port map (
            O => \N__41506\,
            I => \N__41500\
        );

    \I__7680\ : InMux
    port map (
            O => \N__41505\,
            I => \N__41500\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__41500\,
            I => \N__41497\
        );

    \I__7678\ : Span4Mux_v
    port map (
            O => \N__41497\,
            I => \N__41492\
        );

    \I__7677\ : InMux
    port map (
            O => \N__41496\,
            I => \N__41489\
        );

    \I__7676\ : InMux
    port map (
            O => \N__41495\,
            I => \N__41486\
        );

    \I__7675\ : Span4Mux_h
    port map (
            O => \N__41492\,
            I => \N__41483\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__41489\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__41486\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__7672\ : Odrv4
    port map (
            O => \N__41483\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__7671\ : InMux
    port map (
            O => \N__41476\,
            I => \N__41473\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__41473\,
            I => \N__41453\
        );

    \I__7669\ : InMux
    port map (
            O => \N__41472\,
            I => \N__41450\
        );

    \I__7668\ : InMux
    port map (
            O => \N__41471\,
            I => \N__41444\
        );

    \I__7667\ : InMux
    port map (
            O => \N__41470\,
            I => \N__41444\
        );

    \I__7666\ : InMux
    port map (
            O => \N__41469\,
            I => \N__41441\
        );

    \I__7665\ : InMux
    port map (
            O => \N__41468\,
            I => \N__41436\
        );

    \I__7664\ : InMux
    port map (
            O => \N__41467\,
            I => \N__41436\
        );

    \I__7663\ : InMux
    port map (
            O => \N__41466\,
            I => \N__41430\
        );

    \I__7662\ : InMux
    port map (
            O => \N__41465\,
            I => \N__41423\
        );

    \I__7661\ : InMux
    port map (
            O => \N__41464\,
            I => \N__41423\
        );

    \I__7660\ : InMux
    port map (
            O => \N__41463\,
            I => \N__41414\
        );

    \I__7659\ : InMux
    port map (
            O => \N__41462\,
            I => \N__41414\
        );

    \I__7658\ : InMux
    port map (
            O => \N__41461\,
            I => \N__41414\
        );

    \I__7657\ : InMux
    port map (
            O => \N__41460\,
            I => \N__41414\
        );

    \I__7656\ : InMux
    port map (
            O => \N__41459\,
            I => \N__41405\
        );

    \I__7655\ : InMux
    port map (
            O => \N__41458\,
            I => \N__41405\
        );

    \I__7654\ : InMux
    port map (
            O => \N__41457\,
            I => \N__41405\
        );

    \I__7653\ : InMux
    port map (
            O => \N__41456\,
            I => \N__41405\
        );

    \I__7652\ : Span4Mux_v
    port map (
            O => \N__41453\,
            I => \N__41400\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__41450\,
            I => \N__41397\
        );

    \I__7650\ : InMux
    port map (
            O => \N__41449\,
            I => \N__41394\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__41444\,
            I => \N__41390\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__41441\,
            I => \N__41387\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__41436\,
            I => \N__41384\
        );

    \I__7646\ : InMux
    port map (
            O => \N__41435\,
            I => \N__41381\
        );

    \I__7645\ : InMux
    port map (
            O => \N__41434\,
            I => \N__41378\
        );

    \I__7644\ : InMux
    port map (
            O => \N__41433\,
            I => \N__41375\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__41430\,
            I => \N__41372\
        );

    \I__7642\ : InMux
    port map (
            O => \N__41429\,
            I => \N__41369\
        );

    \I__7641\ : InMux
    port map (
            O => \N__41428\,
            I => \N__41366\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__41423\,
            I => \N__41358\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__41414\,
            I => \N__41358\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__41405\,
            I => \N__41358\
        );

    \I__7637\ : InMux
    port map (
            O => \N__41404\,
            I => \N__41355\
        );

    \I__7636\ : InMux
    port map (
            O => \N__41403\,
            I => \N__41352\
        );

    \I__7635\ : Span4Mux_v
    port map (
            O => \N__41400\,
            I => \N__41345\
        );

    \I__7634\ : Span4Mux_v
    port map (
            O => \N__41397\,
            I => \N__41345\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__41394\,
            I => \N__41345\
        );

    \I__7632\ : InMux
    port map (
            O => \N__41393\,
            I => \N__41342\
        );

    \I__7631\ : Span4Mux_h
    port map (
            O => \N__41390\,
            I => \N__41339\
        );

    \I__7630\ : Span4Mux_h
    port map (
            O => \N__41387\,
            I => \N__41330\
        );

    \I__7629\ : Span4Mux_v
    port map (
            O => \N__41384\,
            I => \N__41330\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__41381\,
            I => \N__41330\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__41378\,
            I => \N__41330\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__41375\,
            I => \N__41327\
        );

    \I__7625\ : Span4Mux_h
    port map (
            O => \N__41372\,
            I => \N__41320\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__41369\,
            I => \N__41320\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__41366\,
            I => \N__41320\
        );

    \I__7622\ : InMux
    port map (
            O => \N__41365\,
            I => \N__41317\
        );

    \I__7621\ : Span4Mux_v
    port map (
            O => \N__41358\,
            I => \N__41310\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__41355\,
            I => \N__41310\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__41352\,
            I => \N__41310\
        );

    \I__7618\ : Sp12to4
    port map (
            O => \N__41345\,
            I => \N__41305\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__41342\,
            I => \N__41305\
        );

    \I__7616\ : Span4Mux_h
    port map (
            O => \N__41339\,
            I => \N__41298\
        );

    \I__7615\ : Span4Mux_h
    port map (
            O => \N__41330\,
            I => \N__41298\
        );

    \I__7614\ : Span4Mux_h
    port map (
            O => \N__41327\,
            I => \N__41298\
        );

    \I__7613\ : Span4Mux_v
    port map (
            O => \N__41320\,
            I => \N__41291\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__41317\,
            I => \N__41291\
        );

    \I__7611\ : Span4Mux_h
    port map (
            O => \N__41310\,
            I => \N__41291\
        );

    \I__7610\ : Odrv12
    port map (
            O => \N__41305\,
            I => \c0.n14\
        );

    \I__7609\ : Odrv4
    port map (
            O => \N__41298\,
            I => \c0.n14\
        );

    \I__7608\ : Odrv4
    port map (
            O => \N__41291\,
            I => \c0.n14\
        );

    \I__7607\ : SRMux
    port map (
            O => \N__41284\,
            I => \N__41281\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__41281\,
            I => \N__41278\
        );

    \I__7605\ : Odrv12
    port map (
            O => \N__41278\,
            I => \c0.n18667\
        );

    \I__7604\ : CascadeMux
    port map (
            O => \N__41275\,
            I => \N__41272\
        );

    \I__7603\ : InMux
    port map (
            O => \N__41272\,
            I => \N__41269\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__41269\,
            I => \N__41266\
        );

    \I__7601\ : Span4Mux_h
    port map (
            O => \N__41266\,
            I => \N__41263\
        );

    \I__7600\ : Odrv4
    port map (
            O => \N__41263\,
            I => \c0.n94\
        );

    \I__7599\ : InMux
    port map (
            O => \N__41260\,
            I => \N__41257\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__41257\,
            I => \c0.n12_adj_3004\
        );

    \I__7597\ : InMux
    port map (
            O => \N__41254\,
            I => \N__41251\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__41251\,
            I => \c0.n20_adj_3539\
        );

    \I__7595\ : CascadeMux
    port map (
            O => \N__41248\,
            I => \c0.n12_adj_3001_cascade_\
        );

    \I__7594\ : CascadeMux
    port map (
            O => \N__41245\,
            I => \c0.n20403_cascade_\
        );

    \I__7593\ : InMux
    port map (
            O => \N__41242\,
            I => \N__41239\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__41239\,
            I => \c0.n10_adj_3514\
        );

    \I__7591\ : CascadeMux
    port map (
            O => \N__41236\,
            I => \c0.n20398_cascade_\
        );

    \I__7590\ : CascadeMux
    port map (
            O => \N__41233\,
            I => \N__41229\
        );

    \I__7589\ : InMux
    port map (
            O => \N__41232\,
            I => \N__41224\
        );

    \I__7588\ : InMux
    port map (
            O => \N__41229\,
            I => \N__41224\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__41224\,
            I => \N__41221\
        );

    \I__7586\ : Odrv4
    port map (
            O => \N__41221\,
            I => \c0.n4_adj_3071\
        );

    \I__7585\ : InMux
    port map (
            O => \N__41218\,
            I => \N__41213\
        );

    \I__7584\ : InMux
    port map (
            O => \N__41217\,
            I => \N__41208\
        );

    \I__7583\ : InMux
    port map (
            O => \N__41216\,
            I => \N__41208\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__41213\,
            I => \c0.n5_adj_3003\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__41208\,
            I => \c0.n5_adj_3003\
        );

    \I__7580\ : CascadeMux
    port map (
            O => \N__41203\,
            I => \c0.n36_adj_3267_cascade_\
        );

    \I__7579\ : InMux
    port map (
            O => \N__41200\,
            I => \N__41197\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__41197\,
            I => \c0.n6_adj_3005\
        );

    \I__7577\ : CascadeMux
    port map (
            O => \N__41194\,
            I => \N__41191\
        );

    \I__7576\ : InMux
    port map (
            O => \N__41191\,
            I => \N__41185\
        );

    \I__7575\ : InMux
    port map (
            O => \N__41190\,
            I => \N__41185\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__41185\,
            I => \c0.n13\
        );

    \I__7573\ : CascadeMux
    port map (
            O => \N__41182\,
            I => \c0.n36_adj_3547_cascade_\
        );

    \I__7572\ : InMux
    port map (
            O => \N__41179\,
            I => \N__41176\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__41176\,
            I => \N__41173\
        );

    \I__7570\ : Span4Mux_v
    port map (
            O => \N__41173\,
            I => \N__41170\
        );

    \I__7569\ : Odrv4
    port map (
            O => \N__41170\,
            I => \c0.n63_adj_3417\
        );

    \I__7568\ : CascadeMux
    port map (
            O => \N__41167\,
            I => \c0.n38_adj_3548_cascade_\
        );

    \I__7567\ : InMux
    port map (
            O => \N__41164\,
            I => \N__41161\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__41161\,
            I => \N__41158\
        );

    \I__7565\ : Span4Mux_h
    port map (
            O => \N__41158\,
            I => \N__41155\
        );

    \I__7564\ : Odrv4
    port map (
            O => \N__41155\,
            I => \c0.n34_adj_3411\
        );

    \I__7563\ : CascadeMux
    port map (
            O => \N__41152\,
            I => \c0.n18443_cascade_\
        );

    \I__7562\ : InMux
    port map (
            O => \N__41149\,
            I => \N__41146\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__41146\,
            I => \c0.n25_adj_3495\
        );

    \I__7560\ : InMux
    port map (
            O => \N__41143\,
            I => \N__41138\
        );

    \I__7559\ : InMux
    port map (
            O => \N__41142\,
            I => \N__41135\
        );

    \I__7558\ : InMux
    port map (
            O => \N__41141\,
            I => \N__41132\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__41138\,
            I => \N__41128\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__41135\,
            I => \N__41125\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__41132\,
            I => \N__41121\
        );

    \I__7554\ : InMux
    port map (
            O => \N__41131\,
            I => \N__41118\
        );

    \I__7553\ : Span4Mux_v
    port map (
            O => \N__41128\,
            I => \N__41113\
        );

    \I__7552\ : Span4Mux_v
    port map (
            O => \N__41125\,
            I => \N__41113\
        );

    \I__7551\ : InMux
    port map (
            O => \N__41124\,
            I => \N__41110\
        );

    \I__7550\ : Odrv4
    port map (
            O => \N__41121\,
            I => \c0.data_in_frame_9_4\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__41118\,
            I => \c0.data_in_frame_9_4\
        );

    \I__7548\ : Odrv4
    port map (
            O => \N__41113\,
            I => \c0.data_in_frame_9_4\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__41110\,
            I => \c0.data_in_frame_9_4\
        );

    \I__7546\ : CascadeMux
    port map (
            O => \N__41101\,
            I => \c0.n25_adj_3495_cascade_\
        );

    \I__7545\ : CascadeMux
    port map (
            O => \N__41098\,
            I => \N__41091\
        );

    \I__7544\ : CascadeMux
    port map (
            O => \N__41097\,
            I => \N__41088\
        );

    \I__7543\ : InMux
    port map (
            O => \N__41096\,
            I => \N__41083\
        );

    \I__7542\ : InMux
    port map (
            O => \N__41095\,
            I => \N__41080\
        );

    \I__7541\ : InMux
    port map (
            O => \N__41094\,
            I => \N__41077\
        );

    \I__7540\ : InMux
    port map (
            O => \N__41091\,
            I => \N__41068\
        );

    \I__7539\ : InMux
    port map (
            O => \N__41088\,
            I => \N__41068\
        );

    \I__7538\ : InMux
    port map (
            O => \N__41087\,
            I => \N__41068\
        );

    \I__7537\ : InMux
    port map (
            O => \N__41086\,
            I => \N__41068\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__41083\,
            I => n21222
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__41080\,
            I => n21222
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__41077\,
            I => n21222
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__41068\,
            I => n21222
        );

    \I__7532\ : InMux
    port map (
            O => \N__41059\,
            I => \N__41056\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__41056\,
            I => \N__41053\
        );

    \I__7530\ : Span4Mux_h
    port map (
            O => \N__41053\,
            I => \N__41050\
        );

    \I__7529\ : Span4Mux_h
    port map (
            O => \N__41050\,
            I => \N__41046\
        );

    \I__7528\ : InMux
    port map (
            O => \N__41049\,
            I => \N__41043\
        );

    \I__7527\ : Odrv4
    port map (
            O => \N__41046\,
            I => control_mode_1
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__41043\,
            I => control_mode_1
        );

    \I__7525\ : InMux
    port map (
            O => \N__41038\,
            I => \N__41035\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__41035\,
            I => \c0.n16_adj_3018\
        );

    \I__7523\ : CascadeMux
    port map (
            O => \N__41032\,
            I => \c0.n32_adj_3493_cascade_\
        );

    \I__7522\ : InMux
    port map (
            O => \N__41029\,
            I => \N__41024\
        );

    \I__7521\ : InMux
    port map (
            O => \N__41028\,
            I => \N__41019\
        );

    \I__7520\ : InMux
    port map (
            O => \N__41027\,
            I => \N__41019\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__41024\,
            I => \c0.n20209\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__41019\,
            I => \c0.n20209\
        );

    \I__7517\ : InMux
    port map (
            O => \N__41014\,
            I => \N__41011\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__41011\,
            I => \N__41008\
        );

    \I__7515\ : Odrv4
    port map (
            O => \N__41008\,
            I => \c0.n20204\
        );

    \I__7514\ : CascadeMux
    port map (
            O => \N__41005\,
            I => \c0.n19217_cascade_\
        );

    \I__7513\ : InMux
    port map (
            O => \N__41002\,
            I => \N__40996\
        );

    \I__7512\ : InMux
    port map (
            O => \N__41001\,
            I => \N__40996\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__40996\,
            I => \N__40992\
        );

    \I__7510\ : InMux
    port map (
            O => \N__40995\,
            I => \N__40989\
        );

    \I__7509\ : Odrv12
    port map (
            O => \N__40992\,
            I => \c0.n66\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__40989\,
            I => \c0.n66\
        );

    \I__7507\ : CascadeMux
    port map (
            O => \N__40984\,
            I => \c0.data_out_frame_28__0__N_708_cascade_\
        );

    \I__7506\ : InMux
    port map (
            O => \N__40981\,
            I => \N__40978\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__40978\,
            I => \c0.data_out_frame_28__0__N_708\
        );

    \I__7504\ : InMux
    port map (
            O => \N__40975\,
            I => \N__40972\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__40972\,
            I => \N__40969\
        );

    \I__7502\ : Span12Mux_v
    port map (
            O => \N__40969\,
            I => \N__40966\
        );

    \I__7501\ : Odrv12
    port map (
            O => \N__40966\,
            I => \c0.data_out_frame_29_0\
        );

    \I__7500\ : InMux
    port map (
            O => \N__40963\,
            I => \N__40960\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__40960\,
            I => \c0.data_out_frame_29_1\
        );

    \I__7498\ : InMux
    port map (
            O => \N__40957\,
            I => \N__40953\
        );

    \I__7497\ : InMux
    port map (
            O => \N__40956\,
            I => \N__40950\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__40953\,
            I => \N__40945\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__40950\,
            I => \N__40945\
        );

    \I__7494\ : Odrv4
    port map (
            O => \N__40945\,
            I => data_out_frame_28_1
        );

    \I__7493\ : InMux
    port map (
            O => \N__40942\,
            I => \N__40939\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__40939\,
            I => \N__40932\
        );

    \I__7491\ : InMux
    port map (
            O => \N__40938\,
            I => \N__40927\
        );

    \I__7490\ : InMux
    port map (
            O => \N__40937\,
            I => \N__40927\
        );

    \I__7489\ : CascadeMux
    port map (
            O => \N__40936\,
            I => \N__40920\
        );

    \I__7488\ : InMux
    port map (
            O => \N__40935\,
            I => \N__40916\
        );

    \I__7487\ : Span4Mux_v
    port map (
            O => \N__40932\,
            I => \N__40909\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__40927\,
            I => \N__40909\
        );

    \I__7485\ : InMux
    port map (
            O => \N__40926\,
            I => \N__40901\
        );

    \I__7484\ : InMux
    port map (
            O => \N__40925\,
            I => \N__40897\
        );

    \I__7483\ : InMux
    port map (
            O => \N__40924\,
            I => \N__40894\
        );

    \I__7482\ : InMux
    port map (
            O => \N__40923\,
            I => \N__40887\
        );

    \I__7481\ : InMux
    port map (
            O => \N__40920\,
            I => \N__40887\
        );

    \I__7480\ : InMux
    port map (
            O => \N__40919\,
            I => \N__40877\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__40916\,
            I => \N__40874\
        );

    \I__7478\ : InMux
    port map (
            O => \N__40915\,
            I => \N__40869\
        );

    \I__7477\ : InMux
    port map (
            O => \N__40914\,
            I => \N__40869\
        );

    \I__7476\ : Span4Mux_v
    port map (
            O => \N__40909\,
            I => \N__40866\
        );

    \I__7475\ : InMux
    port map (
            O => \N__40908\,
            I => \N__40861\
        );

    \I__7474\ : InMux
    port map (
            O => \N__40907\,
            I => \N__40861\
        );

    \I__7473\ : InMux
    port map (
            O => \N__40906\,
            I => \N__40858\
        );

    \I__7472\ : InMux
    port map (
            O => \N__40905\,
            I => \N__40850\
        );

    \I__7471\ : InMux
    port map (
            O => \N__40904\,
            I => \N__40847\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__40901\,
            I => \N__40841\
        );

    \I__7469\ : InMux
    port map (
            O => \N__40900\,
            I => \N__40838\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__40897\,
            I => \N__40833\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__40894\,
            I => \N__40833\
        );

    \I__7466\ : InMux
    port map (
            O => \N__40893\,
            I => \N__40830\
        );

    \I__7465\ : InMux
    port map (
            O => \N__40892\,
            I => \N__40827\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__40887\,
            I => \N__40820\
        );

    \I__7463\ : InMux
    port map (
            O => \N__40886\,
            I => \N__40817\
        );

    \I__7462\ : InMux
    port map (
            O => \N__40885\,
            I => \N__40814\
        );

    \I__7461\ : InMux
    port map (
            O => \N__40884\,
            I => \N__40811\
        );

    \I__7460\ : InMux
    port map (
            O => \N__40883\,
            I => \N__40806\
        );

    \I__7459\ : InMux
    port map (
            O => \N__40882\,
            I => \N__40806\
        );

    \I__7458\ : InMux
    port map (
            O => \N__40881\,
            I => \N__40801\
        );

    \I__7457\ : InMux
    port map (
            O => \N__40880\,
            I => \N__40801\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__40877\,
            I => \N__40794\
        );

    \I__7455\ : Span4Mux_v
    port map (
            O => \N__40874\,
            I => \N__40794\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__40869\,
            I => \N__40794\
        );

    \I__7453\ : Span4Mux_h
    port map (
            O => \N__40866\,
            I => \N__40787\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__40861\,
            I => \N__40787\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__40858\,
            I => \N__40787\
        );

    \I__7450\ : InMux
    port map (
            O => \N__40857\,
            I => \N__40784\
        );

    \I__7449\ : InMux
    port map (
            O => \N__40856\,
            I => \N__40781\
        );

    \I__7448\ : InMux
    port map (
            O => \N__40855\,
            I => \N__40774\
        );

    \I__7447\ : InMux
    port map (
            O => \N__40854\,
            I => \N__40774\
        );

    \I__7446\ : InMux
    port map (
            O => \N__40853\,
            I => \N__40774\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__40850\,
            I => \N__40771\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__40847\,
            I => \N__40768\
        );

    \I__7443\ : InMux
    port map (
            O => \N__40846\,
            I => \N__40761\
        );

    \I__7442\ : InMux
    port map (
            O => \N__40845\,
            I => \N__40761\
        );

    \I__7441\ : InMux
    port map (
            O => \N__40844\,
            I => \N__40761\
        );

    \I__7440\ : Span4Mux_h
    port map (
            O => \N__40841\,
            I => \N__40754\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__40838\,
            I => \N__40754\
        );

    \I__7438\ : Span4Mux_v
    port map (
            O => \N__40833\,
            I => \N__40754\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__40830\,
            I => \N__40749\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__40827\,
            I => \N__40749\
        );

    \I__7435\ : InMux
    port map (
            O => \N__40826\,
            I => \N__40746\
        );

    \I__7434\ : CascadeMux
    port map (
            O => \N__40825\,
            I => \N__40743\
        );

    \I__7433\ : InMux
    port map (
            O => \N__40824\,
            I => \N__40740\
        );

    \I__7432\ : InMux
    port map (
            O => \N__40823\,
            I => \N__40735\
        );

    \I__7431\ : Span4Mux_v
    port map (
            O => \N__40820\,
            I => \N__40732\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__40817\,
            I => \N__40729\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__40814\,
            I => \N__40716\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__40811\,
            I => \N__40716\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__40806\,
            I => \N__40716\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__40801\,
            I => \N__40716\
        );

    \I__7425\ : Span4Mux_h
    port map (
            O => \N__40794\,
            I => \N__40716\
        );

    \I__7424\ : Span4Mux_h
    port map (
            O => \N__40787\,
            I => \N__40716\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__40784\,
            I => \N__40707\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__40781\,
            I => \N__40707\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__40774\,
            I => \N__40707\
        );

    \I__7420\ : Span4Mux_v
    port map (
            O => \N__40771\,
            I => \N__40707\
        );

    \I__7419\ : Span4Mux_v
    port map (
            O => \N__40768\,
            I => \N__40696\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__40761\,
            I => \N__40696\
        );

    \I__7417\ : Span4Mux_v
    port map (
            O => \N__40754\,
            I => \N__40696\
        );

    \I__7416\ : Span4Mux_h
    port map (
            O => \N__40749\,
            I => \N__40696\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__40746\,
            I => \N__40696\
        );

    \I__7414\ : InMux
    port map (
            O => \N__40743\,
            I => \N__40693\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__40740\,
            I => \N__40690\
        );

    \I__7412\ : InMux
    port map (
            O => \N__40739\,
            I => \N__40687\
        );

    \I__7411\ : InMux
    port map (
            O => \N__40738\,
            I => \N__40684\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__40735\,
            I => \N__40679\
        );

    \I__7409\ : Span4Mux_h
    port map (
            O => \N__40732\,
            I => \N__40679\
        );

    \I__7408\ : Span4Mux_h
    port map (
            O => \N__40729\,
            I => \N__40674\
        );

    \I__7407\ : Span4Mux_v
    port map (
            O => \N__40716\,
            I => \N__40674\
        );

    \I__7406\ : Span4Mux_v
    port map (
            O => \N__40707\,
            I => \N__40669\
        );

    \I__7405\ : Span4Mux_v
    port map (
            O => \N__40696\,
            I => \N__40669\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__40693\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7403\ : Odrv4
    port map (
            O => \N__40690\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__40687\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__40684\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7400\ : Odrv4
    port map (
            O => \N__40679\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7399\ : Odrv4
    port map (
            O => \N__40674\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7398\ : Odrv4
    port map (
            O => \N__40669\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7397\ : InMux
    port map (
            O => \N__40654\,
            I => \N__40651\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__40651\,
            I => \N__40648\
        );

    \I__7395\ : Span4Mux_v
    port map (
            O => \N__40648\,
            I => \N__40645\
        );

    \I__7394\ : Odrv4
    port map (
            O => \N__40645\,
            I => \c0.n26_adj_3103\
        );

    \I__7393\ : CascadeMux
    port map (
            O => \N__40642\,
            I => \c0.n20246_cascade_\
        );

    \I__7392\ : CascadeMux
    port map (
            O => \N__40639\,
            I => \N__40636\
        );

    \I__7391\ : InMux
    port map (
            O => \N__40636\,
            I => \N__40633\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__40633\,
            I => \c0.n24_adj_3327\
        );

    \I__7389\ : CascadeMux
    port map (
            O => \N__40630\,
            I => \c0.n23_adj_3039_cascade_\
        );

    \I__7388\ : InMux
    port map (
            O => \N__40627\,
            I => \N__40624\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__40624\,
            I => \c0.n23_adj_3039\
        );

    \I__7386\ : InMux
    port map (
            O => \N__40621\,
            I => \N__40618\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__40618\,
            I => \c0.n30_adj_3042\
        );

    \I__7384\ : CascadeMux
    port map (
            O => \N__40615\,
            I => \N__40611\
        );

    \I__7383\ : InMux
    port map (
            O => \N__40614\,
            I => \N__40608\
        );

    \I__7382\ : InMux
    port map (
            O => \N__40611\,
            I => \N__40605\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__40608\,
            I => data_out_frame_29_2
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__40605\,
            I => data_out_frame_29_2
        );

    \I__7379\ : CascadeMux
    port map (
            O => \N__40600\,
            I => \c0.n18428_cascade_\
        );

    \I__7378\ : InMux
    port map (
            O => \N__40597\,
            I => \N__40594\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__40594\,
            I => \c0.n29_adj_3446\
        );

    \I__7376\ : InMux
    port map (
            O => \N__40591\,
            I => \N__40587\
        );

    \I__7375\ : InMux
    port map (
            O => \N__40590\,
            I => \N__40584\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__40587\,
            I => data_out_frame_28_2
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__40584\,
            I => data_out_frame_28_2
        );

    \I__7372\ : InMux
    port map (
            O => \N__40579\,
            I => \N__40576\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__40576\,
            I => \N__40570\
        );

    \I__7370\ : InMux
    port map (
            O => \N__40575\,
            I => \N__40567\
        );

    \I__7369\ : InMux
    port map (
            O => \N__40574\,
            I => \N__40562\
        );

    \I__7368\ : InMux
    port map (
            O => \N__40573\,
            I => \N__40562\
        );

    \I__7367\ : Odrv4
    port map (
            O => \N__40570\,
            I => data_in_0_5
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__40567\,
            I => data_in_0_5
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__40562\,
            I => data_in_0_5
        );

    \I__7364\ : InMux
    port map (
            O => \N__40555\,
            I => \N__40537\
        );

    \I__7363\ : InMux
    port map (
            O => \N__40554\,
            I => \N__40534\
        );

    \I__7362\ : InMux
    port map (
            O => \N__40553\,
            I => \N__40530\
        );

    \I__7361\ : InMux
    port map (
            O => \N__40552\,
            I => \N__40519\
        );

    \I__7360\ : InMux
    port map (
            O => \N__40551\,
            I => \N__40516\
        );

    \I__7359\ : InMux
    port map (
            O => \N__40550\,
            I => \N__40512\
        );

    \I__7358\ : InMux
    port map (
            O => \N__40549\,
            I => \N__40509\
        );

    \I__7357\ : InMux
    port map (
            O => \N__40548\,
            I => \N__40506\
        );

    \I__7356\ : InMux
    port map (
            O => \N__40547\,
            I => \N__40503\
        );

    \I__7355\ : InMux
    port map (
            O => \N__40546\,
            I => \N__40500\
        );

    \I__7354\ : InMux
    port map (
            O => \N__40545\,
            I => \N__40497\
        );

    \I__7353\ : InMux
    port map (
            O => \N__40544\,
            I => \N__40494\
        );

    \I__7352\ : InMux
    port map (
            O => \N__40543\,
            I => \N__40491\
        );

    \I__7351\ : InMux
    port map (
            O => \N__40542\,
            I => \N__40487\
        );

    \I__7350\ : InMux
    port map (
            O => \N__40541\,
            I => \N__40484\
        );

    \I__7349\ : InMux
    port map (
            O => \N__40540\,
            I => \N__40481\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__40537\,
            I => \N__40477\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__40534\,
            I => \N__40474\
        );

    \I__7346\ : InMux
    port map (
            O => \N__40533\,
            I => \N__40471\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__40530\,
            I => \N__40468\
        );

    \I__7344\ : InMux
    port map (
            O => \N__40529\,
            I => \N__40465\
        );

    \I__7343\ : InMux
    port map (
            O => \N__40528\,
            I => \N__40462\
        );

    \I__7342\ : InMux
    port map (
            O => \N__40527\,
            I => \N__40459\
        );

    \I__7341\ : InMux
    port map (
            O => \N__40526\,
            I => \N__40456\
        );

    \I__7340\ : InMux
    port map (
            O => \N__40525\,
            I => \N__40453\
        );

    \I__7339\ : InMux
    port map (
            O => \N__40524\,
            I => \N__40450\
        );

    \I__7338\ : InMux
    port map (
            O => \N__40523\,
            I => \N__40447\
        );

    \I__7337\ : InMux
    port map (
            O => \N__40522\,
            I => \N__40444\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__40519\,
            I => \N__40440\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__40516\,
            I => \N__40437\
        );

    \I__7334\ : InMux
    port map (
            O => \N__40515\,
            I => \N__40434\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__40512\,
            I => \N__40423\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__40509\,
            I => \N__40423\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__40506\,
            I => \N__40423\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__40503\,
            I => \N__40423\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__40500\,
            I => \N__40423\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__40497\,
            I => \N__40420\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__40494\,
            I => \N__40415\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__40491\,
            I => \N__40415\
        );

    \I__7325\ : InMux
    port map (
            O => \N__40490\,
            I => \N__40412\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__40487\,
            I => \N__40409\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__40484\,
            I => \N__40404\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__40481\,
            I => \N__40404\
        );

    \I__7321\ : InMux
    port map (
            O => \N__40480\,
            I => \N__40401\
        );

    \I__7320\ : Span4Mux_v
    port map (
            O => \N__40477\,
            I => \N__40396\
        );

    \I__7319\ : Span4Mux_v
    port map (
            O => \N__40474\,
            I => \N__40396\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__40471\,
            I => \N__40393\
        );

    \I__7317\ : Span4Mux_v
    port map (
            O => \N__40468\,
            I => \N__40374\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__40465\,
            I => \N__40374\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__40462\,
            I => \N__40374\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__40459\,
            I => \N__40374\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__40456\,
            I => \N__40374\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__40453\,
            I => \N__40374\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__40450\,
            I => \N__40374\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__40447\,
            I => \N__40374\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__40444\,
            I => \N__40374\
        );

    \I__7308\ : InMux
    port map (
            O => \N__40443\,
            I => \N__40371\
        );

    \I__7307\ : Span12Mux_s11_v
    port map (
            O => \N__40440\,
            I => \N__40368\
        );

    \I__7306\ : Span4Mux_h
    port map (
            O => \N__40437\,
            I => \N__40365\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__40434\,
            I => \N__40362\
        );

    \I__7304\ : Span4Mux_v
    port map (
            O => \N__40423\,
            I => \N__40353\
        );

    \I__7303\ : Span4Mux_h
    port map (
            O => \N__40420\,
            I => \N__40353\
        );

    \I__7302\ : Span4Mux_h
    port map (
            O => \N__40415\,
            I => \N__40353\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__40412\,
            I => \N__40353\
        );

    \I__7300\ : Span4Mux_v
    port map (
            O => \N__40409\,
            I => \N__40346\
        );

    \I__7299\ : Span4Mux_v
    port map (
            O => \N__40404\,
            I => \N__40346\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__40401\,
            I => \N__40346\
        );

    \I__7297\ : Span4Mux_h
    port map (
            O => \N__40396\,
            I => \N__40337\
        );

    \I__7296\ : Span4Mux_v
    port map (
            O => \N__40393\,
            I => \N__40337\
        );

    \I__7295\ : Span4Mux_v
    port map (
            O => \N__40374\,
            I => \N__40337\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__40371\,
            I => \N__40337\
        );

    \I__7293\ : Odrv12
    port map (
            O => \N__40368\,
            I => \c0.n5_adj_2999\
        );

    \I__7292\ : Odrv4
    port map (
            O => \N__40365\,
            I => \c0.n5_adj_2999\
        );

    \I__7291\ : Odrv12
    port map (
            O => \N__40362\,
            I => \c0.n5_adj_2999\
        );

    \I__7290\ : Odrv4
    port map (
            O => \N__40353\,
            I => \c0.n5_adj_2999\
        );

    \I__7289\ : Odrv4
    port map (
            O => \N__40346\,
            I => \c0.n5_adj_2999\
        );

    \I__7288\ : Odrv4
    port map (
            O => \N__40337\,
            I => \c0.n5_adj_2999\
        );

    \I__7287\ : InMux
    port map (
            O => \N__40324\,
            I => \N__40321\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__40321\,
            I => \N__40318\
        );

    \I__7285\ : Span4Mux_v
    port map (
            O => \N__40318\,
            I => \N__40313\
        );

    \I__7284\ : InMux
    port map (
            O => \N__40317\,
            I => \N__40310\
        );

    \I__7283\ : InMux
    port map (
            O => \N__40316\,
            I => \N__40307\
        );

    \I__7282\ : Span4Mux_h
    port map (
            O => \N__40313\,
            I => \N__40304\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__40310\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__40307\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__7279\ : Odrv4
    port map (
            O => \N__40304\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__7278\ : SRMux
    port map (
            O => \N__40297\,
            I => \N__40294\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__40294\,
            I => \N__40291\
        );

    \I__7276\ : Odrv12
    port map (
            O => \N__40291\,
            I => \c0.n18655\
        );

    \I__7275\ : InMux
    port map (
            O => \N__40288\,
            I => \N__40281\
        );

    \I__7274\ : InMux
    port map (
            O => \N__40287\,
            I => \N__40277\
        );

    \I__7273\ : InMux
    port map (
            O => \N__40286\,
            I => \N__40274\
        );

    \I__7272\ : InMux
    port map (
            O => \N__40285\,
            I => \N__40271\
        );

    \I__7271\ : InMux
    port map (
            O => \N__40284\,
            I => \N__40268\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__40281\,
            I => \N__40262\
        );

    \I__7269\ : InMux
    port map (
            O => \N__40280\,
            I => \N__40259\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__40277\,
            I => \N__40252\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__40274\,
            I => \N__40252\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__40271\,
            I => \N__40252\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__40268\,
            I => \N__40249\
        );

    \I__7264\ : InMux
    port map (
            O => \N__40267\,
            I => \N__40246\
        );

    \I__7263\ : InMux
    port map (
            O => \N__40266\,
            I => \N__40243\
        );

    \I__7262\ : CascadeMux
    port map (
            O => \N__40265\,
            I => \N__40240\
        );

    \I__7261\ : Span4Mux_h
    port map (
            O => \N__40262\,
            I => \N__40237\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__40259\,
            I => \N__40232\
        );

    \I__7259\ : Span4Mux_v
    port map (
            O => \N__40252\,
            I => \N__40232\
        );

    \I__7258\ : Span4Mux_h
    port map (
            O => \N__40249\,
            I => \N__40227\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__40246\,
            I => \N__40227\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__40243\,
            I => \N__40224\
        );

    \I__7255\ : InMux
    port map (
            O => \N__40240\,
            I => \N__40221\
        );

    \I__7254\ : Span4Mux_v
    port map (
            O => \N__40237\,
            I => \N__40216\
        );

    \I__7253\ : Span4Mux_v
    port map (
            O => \N__40232\,
            I => \N__40216\
        );

    \I__7252\ : Span4Mux_v
    port map (
            O => \N__40227\,
            I => \N__40213\
        );

    \I__7251\ : Sp12to4
    port map (
            O => \N__40224\,
            I => \N__40210\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__40221\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__7249\ : Odrv4
    port map (
            O => \N__40216\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__7248\ : Odrv4
    port map (
            O => \N__40213\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__7247\ : Odrv12
    port map (
            O => \N__40210\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__7246\ : InMux
    port map (
            O => \N__40201\,
            I => \N__40196\
        );

    \I__7245\ : InMux
    port map (
            O => \N__40200\,
            I => \N__40193\
        );

    \I__7244\ : InMux
    port map (
            O => \N__40199\,
            I => \N__40190\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__40196\,
            I => \N__40187\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__40193\,
            I => \N__40182\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__40190\,
            I => \N__40179\
        );

    \I__7240\ : Span4Mux_v
    port map (
            O => \N__40187\,
            I => \N__40176\
        );

    \I__7239\ : InMux
    port map (
            O => \N__40186\,
            I => \N__40170\
        );

    \I__7238\ : InMux
    port map (
            O => \N__40185\,
            I => \N__40170\
        );

    \I__7237\ : Span4Mux_h
    port map (
            O => \N__40182\,
            I => \N__40165\
        );

    \I__7236\ : Span4Mux_h
    port map (
            O => \N__40179\,
            I => \N__40165\
        );

    \I__7235\ : Span4Mux_v
    port map (
            O => \N__40176\,
            I => \N__40161\
        );

    \I__7234\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40158\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__40170\,
            I => \N__40155\
        );

    \I__7232\ : Sp12to4
    port map (
            O => \N__40165\,
            I => \N__40152\
        );

    \I__7231\ : InMux
    port map (
            O => \N__40164\,
            I => \N__40149\
        );

    \I__7230\ : Span4Mux_v
    port map (
            O => \N__40161\,
            I => \N__40146\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__40158\,
            I => \N__40143\
        );

    \I__7228\ : Span4Mux_h
    port map (
            O => \N__40155\,
            I => \N__40140\
        );

    \I__7227\ : Span12Mux_v
    port map (
            O => \N__40152\,
            I => \N__40137\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__40149\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__7225\ : Odrv4
    port map (
            O => \N__40146\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__7224\ : Odrv12
    port map (
            O => \N__40143\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__7223\ : Odrv4
    port map (
            O => \N__40140\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__7222\ : Odrv12
    port map (
            O => \N__40137\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__7221\ : CascadeMux
    port map (
            O => \N__40126\,
            I => \N__40122\
        );

    \I__7220\ : InMux
    port map (
            O => \N__40125\,
            I => \N__40119\
        );

    \I__7219\ : InMux
    port map (
            O => \N__40122\,
            I => \N__40115\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__40119\,
            I => \N__40112\
        );

    \I__7217\ : CascadeMux
    port map (
            O => \N__40118\,
            I => \N__40107\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__40115\,
            I => \N__40102\
        );

    \I__7215\ : Span4Mux_v
    port map (
            O => \N__40112\,
            I => \N__40102\
        );

    \I__7214\ : InMux
    port map (
            O => \N__40111\,
            I => \N__40099\
        );

    \I__7213\ : InMux
    port map (
            O => \N__40110\,
            I => \N__40096\
        );

    \I__7212\ : InMux
    port map (
            O => \N__40107\,
            I => \N__40093\
        );

    \I__7211\ : Span4Mux_v
    port map (
            O => \N__40102\,
            I => \N__40085\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__40099\,
            I => \N__40085\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__40096\,
            I => \N__40085\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__40093\,
            I => \N__40081\
        );

    \I__7207\ : InMux
    port map (
            O => \N__40092\,
            I => \N__40078\
        );

    \I__7206\ : Span4Mux_h
    port map (
            O => \N__40085\,
            I => \N__40075\
        );

    \I__7205\ : CascadeMux
    port map (
            O => \N__40084\,
            I => \N__40072\
        );

    \I__7204\ : Span4Mux_h
    port map (
            O => \N__40081\,
            I => \N__40068\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__40078\,
            I => \N__40063\
        );

    \I__7202\ : Sp12to4
    port map (
            O => \N__40075\,
            I => \N__40063\
        );

    \I__7201\ : InMux
    port map (
            O => \N__40072\,
            I => \N__40057\
        );

    \I__7200\ : InMux
    port map (
            O => \N__40071\,
            I => \N__40057\
        );

    \I__7199\ : Span4Mux_h
    port map (
            O => \N__40068\,
            I => \N__40054\
        );

    \I__7198\ : Span12Mux_v
    port map (
            O => \N__40063\,
            I => \N__40051\
        );

    \I__7197\ : InMux
    port map (
            O => \N__40062\,
            I => \N__40048\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__40057\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__7195\ : Odrv4
    port map (
            O => \N__40054\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__7194\ : Odrv12
    port map (
            O => \N__40051\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__40048\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__7192\ : CascadeMux
    port map (
            O => \N__40039\,
            I => \c0.n20224_cascade_\
        );

    \I__7191\ : CascadeMux
    port map (
            O => \N__40036\,
            I => \c0.n19_cascade_\
        );

    \I__7190\ : InMux
    port map (
            O => \N__40033\,
            I => \N__40027\
        );

    \I__7189\ : InMux
    port map (
            O => \N__40032\,
            I => \N__40027\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__40027\,
            I => \N__40022\
        );

    \I__7187\ : InMux
    port map (
            O => \N__40026\,
            I => \N__40017\
        );

    \I__7186\ : InMux
    port map (
            O => \N__40025\,
            I => \N__40017\
        );

    \I__7185\ : Odrv4
    port map (
            O => \N__40022\,
            I => data_in_2_3
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__40017\,
            I => data_in_2_3
        );

    \I__7183\ : InMux
    port map (
            O => \N__40012\,
            I => \N__40009\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__40009\,
            I => \N__40005\
        );

    \I__7181\ : InMux
    port map (
            O => \N__40008\,
            I => \N__40000\
        );

    \I__7180\ : Span4Mux_h
    port map (
            O => \N__40005\,
            I => \N__39997\
        );

    \I__7179\ : InMux
    port map (
            O => \N__40004\,
            I => \N__39994\
        );

    \I__7178\ : InMux
    port map (
            O => \N__40003\,
            I => \N__39991\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__40000\,
            I => data_in_1_3
        );

    \I__7176\ : Odrv4
    port map (
            O => \N__39997\,
            I => data_in_1_3
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__39994\,
            I => data_in_1_3
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__39991\,
            I => data_in_1_3
        );

    \I__7173\ : CascadeMux
    port map (
            O => \N__39982\,
            I => \N__39977\
        );

    \I__7172\ : InMux
    port map (
            O => \N__39981\,
            I => \N__39974\
        );

    \I__7171\ : InMux
    port map (
            O => \N__39980\,
            I => \N__39971\
        );

    \I__7170\ : InMux
    port map (
            O => \N__39977\,
            I => \N__39968\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__39974\,
            I => data_in_0_6
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__39971\,
            I => data_in_0_6
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__39968\,
            I => data_in_0_6
        );

    \I__7166\ : InMux
    port map (
            O => \N__39961\,
            I => \N__39955\
        );

    \I__7165\ : InMux
    port map (
            O => \N__39960\,
            I => \N__39955\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__39955\,
            I => \N__39951\
        );

    \I__7163\ : InMux
    port map (
            O => \N__39954\,
            I => \N__39948\
        );

    \I__7162\ : Span4Mux_h
    port map (
            O => \N__39951\,
            I => \N__39945\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__39948\,
            I => data_in_0_3
        );

    \I__7160\ : Odrv4
    port map (
            O => \N__39945\,
            I => data_in_0_3
        );

    \I__7159\ : InMux
    port map (
            O => \N__39940\,
            I => \N__39937\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__39937\,
            I => \c0.n18_adj_3246\
        );

    \I__7157\ : CascadeMux
    port map (
            O => \N__39934\,
            I => \c0.n20_cascade_\
        );

    \I__7156\ : InMux
    port map (
            O => \N__39931\,
            I => \N__39928\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__39928\,
            I => \c0.n16_adj_3247\
        );

    \I__7154\ : InMux
    port map (
            O => \N__39925\,
            I => \N__39919\
        );

    \I__7153\ : InMux
    port map (
            O => \N__39924\,
            I => \N__39919\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__39919\,
            I => \c0.n11311\
        );

    \I__7151\ : CascadeMux
    port map (
            O => \N__39916\,
            I => \N__39910\
        );

    \I__7150\ : InMux
    port map (
            O => \N__39915\,
            I => \N__39905\
        );

    \I__7149\ : InMux
    port map (
            O => \N__39914\,
            I => \N__39905\
        );

    \I__7148\ : InMux
    port map (
            O => \N__39913\,
            I => \N__39900\
        );

    \I__7147\ : InMux
    port map (
            O => \N__39910\,
            I => \N__39900\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__39905\,
            I => data_in_3_2
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__39900\,
            I => data_in_3_2
        );

    \I__7144\ : CascadeMux
    port map (
            O => \N__39895\,
            I => \N__39892\
        );

    \I__7143\ : InMux
    port map (
            O => \N__39892\,
            I => \N__39888\
        );

    \I__7142\ : InMux
    port map (
            O => \N__39891\,
            I => \N__39885\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__39888\,
            I => \N__39880\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__39885\,
            I => \N__39880\
        );

    \I__7139\ : Span4Mux_h
    port map (
            O => \N__39880\,
            I => \N__39876\
        );

    \I__7138\ : InMux
    port map (
            O => \N__39879\,
            I => \N__39873\
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__39876\,
            I => \c0.n105\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__39873\,
            I => \c0.n105\
        );

    \I__7135\ : InMux
    port map (
            O => \N__39868\,
            I => \N__39862\
        );

    \I__7134\ : InMux
    port map (
            O => \N__39867\,
            I => \N__39857\
        );

    \I__7133\ : InMux
    port map (
            O => \N__39866\,
            I => \N__39857\
        );

    \I__7132\ : InMux
    port map (
            O => \N__39865\,
            I => \N__39854\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__39862\,
            I => data_in_3_3
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__39857\,
            I => data_in_3_3
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__39854\,
            I => data_in_3_3
        );

    \I__7128\ : InMux
    port map (
            O => \N__39847\,
            I => \N__39839\
        );

    \I__7127\ : InMux
    port map (
            O => \N__39846\,
            I => \N__39839\
        );

    \I__7126\ : InMux
    port map (
            O => \N__39845\,
            I => \N__39834\
        );

    \I__7125\ : InMux
    port map (
            O => \N__39844\,
            I => \N__39834\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__39839\,
            I => data_in_3_1
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__39834\,
            I => data_in_3_1
        );

    \I__7122\ : CascadeMux
    port map (
            O => \N__39829\,
            I => \N__39825\
        );

    \I__7121\ : CascadeMux
    port map (
            O => \N__39828\,
            I => \N__39821\
        );

    \I__7120\ : InMux
    port map (
            O => \N__39825\,
            I => \N__39818\
        );

    \I__7119\ : InMux
    port map (
            O => \N__39824\,
            I => \N__39813\
        );

    \I__7118\ : InMux
    port map (
            O => \N__39821\,
            I => \N__39813\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__39818\,
            I => data_in_0_7
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__39813\,
            I => data_in_0_7
        );

    \I__7115\ : CascadeMux
    port map (
            O => \N__39808\,
            I => \N__39803\
        );

    \I__7114\ : InMux
    port map (
            O => \N__39807\,
            I => \N__39799\
        );

    \I__7113\ : InMux
    port map (
            O => \N__39806\,
            I => \N__39796\
        );

    \I__7112\ : InMux
    port map (
            O => \N__39803\,
            I => \N__39793\
        );

    \I__7111\ : InMux
    port map (
            O => \N__39802\,
            I => \N__39790\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__39799\,
            I => \N__39787\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__39796\,
            I => \N__39782\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__39793\,
            I => \N__39782\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__39790\,
            I => data_in_1_6
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__39787\,
            I => data_in_1_6
        );

    \I__7105\ : Odrv12
    port map (
            O => \N__39782\,
            I => data_in_1_6
        );

    \I__7104\ : InMux
    port map (
            O => \N__39775\,
            I => \N__39772\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__39772\,
            I => \c0.n18_adj_3229\
        );

    \I__7102\ : CascadeMux
    port map (
            O => \N__39769\,
            I => \N__39766\
        );

    \I__7101\ : InMux
    port map (
            O => \N__39766\,
            I => \N__39760\
        );

    \I__7100\ : InMux
    port map (
            O => \N__39765\,
            I => \N__39760\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__39760\,
            I => \N__39757\
        );

    \I__7098\ : Odrv4
    port map (
            O => \N__39757\,
            I => \c0.n11446\
        );

    \I__7097\ : CascadeMux
    port map (
            O => \N__39754\,
            I => \c0.n21108_cascade_\
        );

    \I__7096\ : InMux
    port map (
            O => \N__39751\,
            I => \N__39748\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__39748\,
            I => \c0.n12_adj_3248\
        );

    \I__7094\ : InMux
    port map (
            O => \N__39745\,
            I => \N__39740\
        );

    \I__7093\ : InMux
    port map (
            O => \N__39744\,
            I => \N__39736\
        );

    \I__7092\ : InMux
    port map (
            O => \N__39743\,
            I => \N__39733\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__39740\,
            I => \N__39730\
        );

    \I__7090\ : InMux
    port map (
            O => \N__39739\,
            I => \N__39727\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__39736\,
            I => \N__39724\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__39733\,
            I => \N__39717\
        );

    \I__7087\ : Span4Mux_v
    port map (
            O => \N__39730\,
            I => \N__39717\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__39727\,
            I => \N__39717\
        );

    \I__7085\ : Odrv12
    port map (
            O => \N__39724\,
            I => data_in_3_5
        );

    \I__7084\ : Odrv4
    port map (
            O => \N__39717\,
            I => data_in_3_5
        );

    \I__7083\ : InMux
    port map (
            O => \N__39712\,
            I => \N__39706\
        );

    \I__7082\ : InMux
    port map (
            O => \N__39711\,
            I => \N__39706\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__39706\,
            I => \c0.n20_adj_3250\
        );

    \I__7080\ : InMux
    port map (
            O => \N__39703\,
            I => \N__39699\
        );

    \I__7079\ : CascadeMux
    port map (
            O => \N__39702\,
            I => \N__39696\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__39699\,
            I => \N__39693\
        );

    \I__7077\ : InMux
    port map (
            O => \N__39696\,
            I => \N__39690\
        );

    \I__7076\ : Span4Mux_h
    port map (
            O => \N__39693\,
            I => \N__39687\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__39690\,
            I => \c0.data_in_frame_28_6\
        );

    \I__7074\ : Odrv4
    port map (
            O => \N__39687\,
            I => \c0.data_in_frame_28_6\
        );

    \I__7073\ : CascadeMux
    port map (
            O => \N__39682\,
            I => \c0.n17947_cascade_\
        );

    \I__7072\ : InMux
    port map (
            O => \N__39679\,
            I => \N__39676\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__39676\,
            I => \N__39673\
        );

    \I__7070\ : Odrv4
    port map (
            O => \N__39673\,
            I => \c0.n20793\
        );

    \I__7069\ : CascadeMux
    port map (
            O => \N__39670\,
            I => \c0.n10_adj_3242_cascade_\
        );

    \I__7068\ : InMux
    port map (
            O => \N__39667\,
            I => \N__39662\
        );

    \I__7067\ : InMux
    port map (
            O => \N__39666\,
            I => \N__39659\
        );

    \I__7066\ : InMux
    port map (
            O => \N__39665\,
            I => \N__39656\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__39662\,
            I => data_in_0_2
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__39659\,
            I => data_in_0_2
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__39656\,
            I => data_in_0_2
        );

    \I__7062\ : InMux
    port map (
            O => \N__39649\,
            I => \N__39646\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__39646\,
            I => \c0.n14_adj_3243\
        );

    \I__7060\ : CascadeMux
    port map (
            O => \N__39643\,
            I => \c0.n36_adj_3277_cascade_\
        );

    \I__7059\ : CascadeMux
    port map (
            O => \N__39640\,
            I => \c0.n20415_cascade_\
        );

    \I__7058\ : CascadeMux
    port map (
            O => \N__39637\,
            I => \c0.n14_adj_3407_cascade_\
        );

    \I__7057\ : InMux
    port map (
            O => \N__39634\,
            I => \N__39631\
        );

    \I__7056\ : LocalMux
    port map (
            O => \N__39631\,
            I => \c0.n100_adj_3403\
        );

    \I__7055\ : CascadeMux
    port map (
            O => \N__39628\,
            I => \N__39625\
        );

    \I__7054\ : InMux
    port map (
            O => \N__39625\,
            I => \N__39622\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__39622\,
            I => \N__39619\
        );

    \I__7052\ : Span4Mux_h
    port map (
            O => \N__39619\,
            I => \N__39616\
        );

    \I__7051\ : Span4Mux_v
    port map (
            O => \N__39616\,
            I => \N__39613\
        );

    \I__7050\ : Odrv4
    port map (
            O => \N__39613\,
            I => \c0.n18_adj_3412\
        );

    \I__7049\ : CascadeMux
    port map (
            O => \N__39610\,
            I => \c0.n20300_cascade_\
        );

    \I__7048\ : CascadeMux
    port map (
            O => \N__39607\,
            I => \N__39604\
        );

    \I__7047\ : InMux
    port map (
            O => \N__39604\,
            I => \N__39601\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__39601\,
            I => \c0.n20300\
        );

    \I__7045\ : CascadeMux
    port map (
            O => \N__39598\,
            I => \N__39591\
        );

    \I__7044\ : CascadeMux
    port map (
            O => \N__39597\,
            I => \N__39587\
        );

    \I__7043\ : InMux
    port map (
            O => \N__39596\,
            I => \N__39582\
        );

    \I__7042\ : InMux
    port map (
            O => \N__39595\,
            I => \N__39582\
        );

    \I__7041\ : InMux
    port map (
            O => \N__39594\,
            I => \N__39577\
        );

    \I__7040\ : InMux
    port map (
            O => \N__39591\,
            I => \N__39577\
        );

    \I__7039\ : InMux
    port map (
            O => \N__39590\,
            I => \N__39573\
        );

    \I__7038\ : InMux
    port map (
            O => \N__39587\,
            I => \N__39570\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__39582\,
            I => \N__39564\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__39577\,
            I => \N__39561\
        );

    \I__7035\ : InMux
    port map (
            O => \N__39576\,
            I => \N__39558\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__39573\,
            I => \N__39553\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__39570\,
            I => \N__39549\
        );

    \I__7032\ : InMux
    port map (
            O => \N__39569\,
            I => \N__39546\
        );

    \I__7031\ : InMux
    port map (
            O => \N__39568\,
            I => \N__39543\
        );

    \I__7030\ : InMux
    port map (
            O => \N__39567\,
            I => \N__39540\
        );

    \I__7029\ : Span4Mux_v
    port map (
            O => \N__39564\,
            I => \N__39537\
        );

    \I__7028\ : Span4Mux_h
    port map (
            O => \N__39561\,
            I => \N__39532\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__39558\,
            I => \N__39532\
        );

    \I__7026\ : InMux
    port map (
            O => \N__39557\,
            I => \N__39529\
        );

    \I__7025\ : InMux
    port map (
            O => \N__39556\,
            I => \N__39526\
        );

    \I__7024\ : Span4Mux_h
    port map (
            O => \N__39553\,
            I => \N__39523\
        );

    \I__7023\ : InMux
    port map (
            O => \N__39552\,
            I => \N__39520\
        );

    \I__7022\ : Span4Mux_h
    port map (
            O => \N__39549\,
            I => \N__39515\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__39546\,
            I => \N__39515\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__39543\,
            I => \N__39512\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__39540\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7018\ : Odrv4
    port map (
            O => \N__39537\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7017\ : Odrv4
    port map (
            O => \N__39532\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__39529\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__39526\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7014\ : Odrv4
    port map (
            O => \N__39523\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__39520\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7012\ : Odrv4
    port map (
            O => \N__39515\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7011\ : Odrv4
    port map (
            O => \N__39512\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7010\ : InMux
    port map (
            O => \N__39493\,
            I => \N__39487\
        );

    \I__7009\ : InMux
    port map (
            O => \N__39492\,
            I => \N__39483\
        );

    \I__7008\ : InMux
    port map (
            O => \N__39491\,
            I => \N__39478\
        );

    \I__7007\ : InMux
    port map (
            O => \N__39490\,
            I => \N__39478\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__39487\,
            I => \N__39475\
        );

    \I__7005\ : InMux
    port map (
            O => \N__39486\,
            I => \N__39472\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__39483\,
            I => \N__39469\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__39478\,
            I => \N__39466\
        );

    \I__7002\ : Span4Mux_v
    port map (
            O => \N__39475\,
            I => \N__39463\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__39472\,
            I => \N__39460\
        );

    \I__7000\ : Span4Mux_h
    port map (
            O => \N__39469\,
            I => \N__39457\
        );

    \I__6999\ : Sp12to4
    port map (
            O => \N__39466\,
            I => \N__39454\
        );

    \I__6998\ : Span4Mux_v
    port map (
            O => \N__39463\,
            I => \N__39449\
        );

    \I__6997\ : Span4Mux_h
    port map (
            O => \N__39460\,
            I => \N__39449\
        );

    \I__6996\ : Span4Mux_h
    port map (
            O => \N__39457\,
            I => \N__39446\
        );

    \I__6995\ : Span12Mux_v
    port map (
            O => \N__39454\,
            I => \N__39443\
        );

    \I__6994\ : Span4Mux_h
    port map (
            O => \N__39449\,
            I => \N__39440\
        );

    \I__6993\ : Odrv4
    port map (
            O => \N__39446\,
            I => \c0.n3235\
        );

    \I__6992\ : Odrv12
    port map (
            O => \N__39443\,
            I => \c0.n3235\
        );

    \I__6991\ : Odrv4
    port map (
            O => \N__39440\,
            I => \c0.n3235\
        );

    \I__6990\ : InMux
    port map (
            O => \N__39433\,
            I => \N__39429\
        );

    \I__6989\ : InMux
    port map (
            O => \N__39432\,
            I => \N__39426\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__39429\,
            I => \N__39423\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__39426\,
            I => \c0.rx.n15860\
        );

    \I__6986\ : Odrv4
    port map (
            O => \N__39423\,
            I => \c0.rx.n15860\
        );

    \I__6985\ : InMux
    port map (
            O => \N__39418\,
            I => \N__39415\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__39415\,
            I => \N__39412\
        );

    \I__6983\ : Span4Mux_v
    port map (
            O => \N__39412\,
            I => \N__39409\
        );

    \I__6982\ : Odrv4
    port map (
            O => \N__39409\,
            I => \c0.n19449\
        );

    \I__6981\ : InMux
    port map (
            O => \N__39406\,
            I => \N__39403\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__39403\,
            I => \N__39398\
        );

    \I__6979\ : InMux
    port map (
            O => \N__39402\,
            I => \N__39393\
        );

    \I__6978\ : InMux
    port map (
            O => \N__39401\,
            I => \N__39393\
        );

    \I__6977\ : Span12Mux_h
    port map (
            O => \N__39398\,
            I => \N__39390\
        );

    \I__6976\ : LocalMux
    port map (
            O => \N__39393\,
            I => \N__39387\
        );

    \I__6975\ : Odrv12
    port map (
            O => \N__39390\,
            I => n12492
        );

    \I__6974\ : Odrv4
    port map (
            O => \N__39387\,
            I => n12492
        );

    \I__6973\ : CascadeMux
    port map (
            O => \N__39382\,
            I => \N__39379\
        );

    \I__6972\ : InMux
    port map (
            O => \N__39379\,
            I => \N__39376\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__39376\,
            I => \N__39371\
        );

    \I__6970\ : InMux
    port map (
            O => \N__39375\,
            I => \N__39366\
        );

    \I__6969\ : InMux
    port map (
            O => \N__39374\,
            I => \N__39366\
        );

    \I__6968\ : Span4Mux_h
    port map (
            O => \N__39371\,
            I => \N__39363\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__39366\,
            I => \N__39360\
        );

    \I__6966\ : Sp12to4
    port map (
            O => \N__39363\,
            I => \N__39357\
        );

    \I__6965\ : Odrv12
    port map (
            O => \N__39360\,
            I => n12835
        );

    \I__6964\ : Odrv12
    port map (
            O => \N__39357\,
            I => n12835
        );

    \I__6963\ : InMux
    port map (
            O => \N__39352\,
            I => \N__39349\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__39349\,
            I => \N__39346\
        );

    \I__6961\ : Span4Mux_h
    port map (
            O => \N__39346\,
            I => \N__39339\
        );

    \I__6960\ : InMux
    port map (
            O => \N__39345\,
            I => \N__39336\
        );

    \I__6959\ : InMux
    port map (
            O => \N__39344\,
            I => \N__39328\
        );

    \I__6958\ : InMux
    port map (
            O => \N__39343\,
            I => \N__39328\
        );

    \I__6957\ : InMux
    port map (
            O => \N__39342\,
            I => \N__39328\
        );

    \I__6956\ : Span4Mux_v
    port map (
            O => \N__39339\,
            I => \N__39325\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__39336\,
            I => \N__39322\
        );

    \I__6954\ : InMux
    port map (
            O => \N__39335\,
            I => \N__39319\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__39328\,
            I => \N__39314\
        );

    \I__6952\ : Span4Mux_v
    port map (
            O => \N__39325\,
            I => \N__39314\
        );

    \I__6951\ : Odrv12
    port map (
            O => \N__39322\,
            I => \r_Bit_Index_0\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__39319\,
            I => \r_Bit_Index_0\
        );

    \I__6949\ : Odrv4
    port map (
            O => \N__39314\,
            I => \r_Bit_Index_0\
        );

    \I__6948\ : CascadeMux
    port map (
            O => \N__39307\,
            I => \c0.n22_adj_3276_cascade_\
        );

    \I__6947\ : InMux
    port map (
            O => \N__39304\,
            I => \N__39301\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__39301\,
            I => \N__39298\
        );

    \I__6945\ : Odrv12
    port map (
            O => \N__39298\,
            I => \c0.n21104\
        );

    \I__6944\ : CascadeMux
    port map (
            O => \N__39295\,
            I => \n3846_cascade_\
        );

    \I__6943\ : InMux
    port map (
            O => \N__39292\,
            I => \N__39286\
        );

    \I__6942\ : InMux
    port map (
            O => \N__39291\,
            I => \N__39280\
        );

    \I__6941\ : InMux
    port map (
            O => \N__39290\,
            I => \N__39277\
        );

    \I__6940\ : InMux
    port map (
            O => \N__39289\,
            I => \N__39274\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__39286\,
            I => \N__39271\
        );

    \I__6938\ : InMux
    port map (
            O => \N__39285\,
            I => \N__39264\
        );

    \I__6937\ : InMux
    port map (
            O => \N__39284\,
            I => \N__39264\
        );

    \I__6936\ : InMux
    port map (
            O => \N__39283\,
            I => \N__39264\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__39280\,
            I => \N__39261\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__39277\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__39274\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__6932\ : Odrv4
    port map (
            O => \N__39271\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__39264\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__6930\ : Odrv4
    port map (
            O => \N__39261\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__6929\ : InMux
    port map (
            O => \N__39250\,
            I => \N__39247\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__39247\,
            I => \c0.rx.n6_adj_2995\
        );

    \I__6927\ : InMux
    port map (
            O => \N__39244\,
            I => \N__39240\
        );

    \I__6926\ : InMux
    port map (
            O => \N__39243\,
            I => \N__39237\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__39240\,
            I => \c0.rx.n11455\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__39237\,
            I => \c0.rx.n11455\
        );

    \I__6923\ : InMux
    port map (
            O => \N__39232\,
            I => \N__39228\
        );

    \I__6922\ : InMux
    port map (
            O => \N__39231\,
            I => \N__39225\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__39228\,
            I => \N__39222\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__39225\,
            I => \N__39216\
        );

    \I__6919\ : Span4Mux_v
    port map (
            O => \N__39222\,
            I => \N__39216\
        );

    \I__6918\ : InMux
    port map (
            O => \N__39221\,
            I => \N__39213\
        );

    \I__6917\ : Span4Mux_h
    port map (
            O => \N__39216\,
            I => \N__39210\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__39213\,
            I => \c0.rx.r_SM_Main_2_N_2479_0\
        );

    \I__6915\ : Odrv4
    port map (
            O => \N__39210\,
            I => \c0.rx.r_SM_Main_2_N_2479_0\
        );

    \I__6914\ : InMux
    port map (
            O => \N__39205\,
            I => \N__39199\
        );

    \I__6913\ : InMux
    port map (
            O => \N__39204\,
            I => \N__39199\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__39199\,
            I => \N__39196\
        );

    \I__6911\ : Span4Mux_v
    port map (
            O => \N__39196\,
            I => \N__39187\
        );

    \I__6910\ : InMux
    port map (
            O => \N__39195\,
            I => \N__39184\
        );

    \I__6909\ : InMux
    port map (
            O => \N__39194\,
            I => \N__39177\
        );

    \I__6908\ : InMux
    port map (
            O => \N__39193\,
            I => \N__39177\
        );

    \I__6907\ : InMux
    port map (
            O => \N__39192\,
            I => \N__39177\
        );

    \I__6906\ : InMux
    port map (
            O => \N__39191\,
            I => \N__39172\
        );

    \I__6905\ : InMux
    port map (
            O => \N__39190\,
            I => \N__39172\
        );

    \I__6904\ : Odrv4
    port map (
            O => \N__39187\,
            I => n3792
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__39184\,
            I => n3792
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__39177\,
            I => n3792
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__39172\,
            I => n3792
        );

    \I__6900\ : InMux
    port map (
            O => \N__39163\,
            I => \N__39160\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__39160\,
            I => \N__39157\
        );

    \I__6898\ : Span4Mux_h
    port map (
            O => \N__39157\,
            I => \N__39154\
        );

    \I__6897\ : Odrv4
    port map (
            O => \N__39154\,
            I => n12911
        );

    \I__6896\ : InMux
    port map (
            O => \N__39151\,
            I => \N__39147\
        );

    \I__6895\ : InMux
    port map (
            O => \N__39150\,
            I => \N__39144\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__39147\,
            I => \N__39137\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__39144\,
            I => \N__39137\
        );

    \I__6892\ : CascadeMux
    port map (
            O => \N__39143\,
            I => \N__39133\
        );

    \I__6891\ : InMux
    port map (
            O => \N__39142\,
            I => \N__39130\
        );

    \I__6890\ : Span4Mux_h
    port map (
            O => \N__39137\,
            I => \N__39127\
        );

    \I__6889\ : InMux
    port map (
            O => \N__39136\,
            I => \N__39124\
        );

    \I__6888\ : InMux
    port map (
            O => \N__39133\,
            I => \N__39121\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__39130\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__6886\ : Odrv4
    port map (
            O => \N__39127\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__39124\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__39121\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__6883\ : InMux
    port map (
            O => \N__39112\,
            I => \N__39109\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__39109\,
            I => \c0.n16\
        );

    \I__6881\ : InMux
    port map (
            O => \N__39106\,
            I => \N__39103\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__39103\,
            I => \c0.n24\
        );

    \I__6879\ : CascadeMux
    port map (
            O => \N__39100\,
            I => \c0.n28_cascade_\
        );

    \I__6878\ : CascadeMux
    port map (
            O => \N__39097\,
            I => \c0.n12026_cascade_\
        );

    \I__6877\ : CascadeMux
    port map (
            O => \N__39094\,
            I => \c0.n10_cascade_\
        );

    \I__6876\ : CascadeMux
    port map (
            O => \N__39091\,
            I => \c0.n19449_cascade_\
        );

    \I__6875\ : InMux
    port map (
            O => \N__39088\,
            I => \N__39084\
        );

    \I__6874\ : InMux
    port map (
            O => \N__39087\,
            I => \N__39081\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__39084\,
            I => control_mode_0
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__39081\,
            I => control_mode_0
        );

    \I__6871\ : CascadeMux
    port map (
            O => \N__39076\,
            I => \N__39072\
        );

    \I__6870\ : InMux
    port map (
            O => \N__39075\,
            I => \N__39068\
        );

    \I__6869\ : InMux
    port map (
            O => \N__39072\,
            I => \N__39065\
        );

    \I__6868\ : InMux
    port map (
            O => \N__39071\,
            I => \N__39061\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__39068\,
            I => \N__39055\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__39065\,
            I => \N__39055\
        );

    \I__6865\ : InMux
    port map (
            O => \N__39064\,
            I => \N__39052\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__39061\,
            I => \N__39049\
        );

    \I__6863\ : InMux
    port map (
            O => \N__39060\,
            I => \N__39046\
        );

    \I__6862\ : Span4Mux_v
    port map (
            O => \N__39055\,
            I => \N__39043\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__39052\,
            I => \N__39040\
        );

    \I__6860\ : Span4Mux_h
    port map (
            O => \N__39049\,
            I => \N__39037\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__39046\,
            I => \N__39032\
        );

    \I__6858\ : Span4Mux_h
    port map (
            O => \N__39043\,
            I => \N__39032\
        );

    \I__6857\ : Span4Mux_v
    port map (
            O => \N__39040\,
            I => \N__39029\
        );

    \I__6856\ : Sp12to4
    port map (
            O => \N__39037\,
            I => \N__39026\
        );

    \I__6855\ : Span4Mux_v
    port map (
            O => \N__39032\,
            I => \N__39023\
        );

    \I__6854\ : Span4Mux_v
    port map (
            O => \N__39029\,
            I => \N__39020\
        );

    \I__6853\ : Span12Mux_v
    port map (
            O => \N__39026\,
            I => \N__39017\
        );

    \I__6852\ : Span4Mux_v
    port map (
            O => \N__39023\,
            I => \N__39014\
        );

    \I__6851\ : Span4Mux_v
    port map (
            O => \N__39020\,
            I => \N__39011\
        );

    \I__6850\ : Odrv12
    port map (
            O => \N__39017\,
            I => \FRAME_MATCHER_state_31_N_1800_2\
        );

    \I__6849\ : Odrv4
    port map (
            O => \N__39014\,
            I => \FRAME_MATCHER_state_31_N_1800_2\
        );

    \I__6848\ : Odrv4
    port map (
            O => \N__39011\,
            I => \FRAME_MATCHER_state_31_N_1800_2\
        );

    \I__6847\ : InMux
    port map (
            O => \N__39004\,
            I => \N__38998\
        );

    \I__6846\ : InMux
    port map (
            O => \N__39003\,
            I => \N__38998\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__38998\,
            I => \N__38993\
        );

    \I__6844\ : InMux
    port map (
            O => \N__38997\,
            I => \N__38990\
        );

    \I__6843\ : CascadeMux
    port map (
            O => \N__38996\,
            I => \N__38986\
        );

    \I__6842\ : Span4Mux_h
    port map (
            O => \N__38993\,
            I => \N__38979\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__38990\,
            I => \N__38979\
        );

    \I__6840\ : CascadeMux
    port map (
            O => \N__38989\,
            I => \N__38973\
        );

    \I__6839\ : InMux
    port map (
            O => \N__38986\,
            I => \N__38969\
        );

    \I__6838\ : CascadeMux
    port map (
            O => \N__38985\,
            I => \N__38965\
        );

    \I__6837\ : InMux
    port map (
            O => \N__38984\,
            I => \N__38961\
        );

    \I__6836\ : Span4Mux_v
    port map (
            O => \N__38979\,
            I => \N__38958\
        );

    \I__6835\ : InMux
    port map (
            O => \N__38978\,
            I => \N__38955\
        );

    \I__6834\ : CascadeMux
    port map (
            O => \N__38977\,
            I => \N__38952\
        );

    \I__6833\ : InMux
    port map (
            O => \N__38976\,
            I => \N__38947\
        );

    \I__6832\ : InMux
    port map (
            O => \N__38973\,
            I => \N__38947\
        );

    \I__6831\ : InMux
    port map (
            O => \N__38972\,
            I => \N__38944\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__38969\,
            I => \N__38941\
        );

    \I__6829\ : InMux
    port map (
            O => \N__38968\,
            I => \N__38938\
        );

    \I__6828\ : InMux
    port map (
            O => \N__38965\,
            I => \N__38935\
        );

    \I__6827\ : CascadeMux
    port map (
            O => \N__38964\,
            I => \N__38932\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__38961\,
            I => \N__38928\
        );

    \I__6825\ : Span4Mux_v
    port map (
            O => \N__38958\,
            I => \N__38922\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__38955\,
            I => \N__38919\
        );

    \I__6823\ : InMux
    port map (
            O => \N__38952\,
            I => \N__38916\
        );

    \I__6822\ : LocalMux
    port map (
            O => \N__38947\,
            I => \N__38913\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__38944\,
            I => \N__38910\
        );

    \I__6820\ : Span4Mux_v
    port map (
            O => \N__38941\,
            I => \N__38905\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__38938\,
            I => \N__38905\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__38935\,
            I => \N__38902\
        );

    \I__6817\ : InMux
    port map (
            O => \N__38932\,
            I => \N__38897\
        );

    \I__6816\ : InMux
    port map (
            O => \N__38931\,
            I => \N__38897\
        );

    \I__6815\ : Span12Mux_v
    port map (
            O => \N__38928\,
            I => \N__38894\
        );

    \I__6814\ : InMux
    port map (
            O => \N__38927\,
            I => \N__38891\
        );

    \I__6813\ : InMux
    port map (
            O => \N__38926\,
            I => \N__38888\
        );

    \I__6812\ : InMux
    port map (
            O => \N__38925\,
            I => \N__38885\
        );

    \I__6811\ : Span4Mux_h
    port map (
            O => \N__38922\,
            I => \N__38880\
        );

    \I__6810\ : Span4Mux_h
    port map (
            O => \N__38919\,
            I => \N__38880\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__38916\,
            I => \N__38875\
        );

    \I__6808\ : Span4Mux_h
    port map (
            O => \N__38913\,
            I => \N__38875\
        );

    \I__6807\ : Span4Mux_v
    port map (
            O => \N__38910\,
            I => \N__38870\
        );

    \I__6806\ : Span4Mux_v
    port map (
            O => \N__38905\,
            I => \N__38870\
        );

    \I__6805\ : Span12Mux_v
    port map (
            O => \N__38902\,
            I => \N__38865\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__38897\,
            I => \N__38865\
        );

    \I__6803\ : Odrv12
    port map (
            O => \N__38894\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__38891\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__38888\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__38885\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__6799\ : Odrv4
    port map (
            O => \N__38880\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__6798\ : Odrv4
    port map (
            O => \N__38875\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__6797\ : Odrv4
    port map (
            O => \N__38870\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__6796\ : Odrv12
    port map (
            O => \N__38865\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__6795\ : InMux
    port map (
            O => \N__38848\,
            I => \N__38845\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__38845\,
            I => \N__38842\
        );

    \I__6793\ : Span4Mux_v
    port map (
            O => \N__38842\,
            I => \N__38838\
        );

    \I__6792\ : InMux
    port map (
            O => \N__38841\,
            I => \N__38834\
        );

    \I__6791\ : Span4Mux_h
    port map (
            O => \N__38838\,
            I => \N__38831\
        );

    \I__6790\ : InMux
    port map (
            O => \N__38837\,
            I => \N__38828\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__38834\,
            I => \N__38825\
        );

    \I__6788\ : Sp12to4
    port map (
            O => \N__38831\,
            I => \N__38818\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__38828\,
            I => \N__38818\
        );

    \I__6786\ : Span12Mux_h
    port map (
            O => \N__38825\,
            I => \N__38818\
        );

    \I__6785\ : Span12Mux_v
    port map (
            O => \N__38818\,
            I => \N__38815\
        );

    \I__6784\ : Odrv12
    port map (
            O => \N__38815\,
            I => \c0.n15499\
        );

    \I__6783\ : InMux
    port map (
            O => \N__38812\,
            I => \N__38809\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__38809\,
            I => \c0.n13_adj_3016\
        );

    \I__6781\ : CascadeMux
    port map (
            O => \N__38806\,
            I => \N__38803\
        );

    \I__6780\ : InMux
    port map (
            O => \N__38803\,
            I => \N__38799\
        );

    \I__6779\ : InMux
    port map (
            O => \N__38802\,
            I => \N__38796\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__38799\,
            I => \N__38793\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__38796\,
            I => \N__38790\
        );

    \I__6776\ : Span4Mux_v
    port map (
            O => \N__38793\,
            I => \N__38787\
        );

    \I__6775\ : Span4Mux_h
    port map (
            O => \N__38790\,
            I => \N__38783\
        );

    \I__6774\ : Span4Mux_v
    port map (
            O => \N__38787\,
            I => \N__38780\
        );

    \I__6773\ : InMux
    port map (
            O => \N__38786\,
            I => \N__38777\
        );

    \I__6772\ : Odrv4
    port map (
            O => \N__38783\,
            I => \c0.FRAME_MATCHER_rx_data_ready_prev\
        );

    \I__6771\ : Odrv4
    port map (
            O => \N__38780\,
            I => \c0.FRAME_MATCHER_rx_data_ready_prev\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__38777\,
            I => \c0.FRAME_MATCHER_rx_data_ready_prev\
        );

    \I__6769\ : CascadeMux
    port map (
            O => \N__38770\,
            I => \c0.n19111_cascade_\
        );

    \I__6768\ : InMux
    port map (
            O => \N__38767\,
            I => \N__38764\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__38764\,
            I => \N__38760\
        );

    \I__6766\ : InMux
    port map (
            O => \N__38763\,
            I => \N__38757\
        );

    \I__6765\ : Odrv12
    port map (
            O => \N__38760\,
            I => \c0.n19493\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__38757\,
            I => \c0.n19493\
        );

    \I__6763\ : InMux
    port map (
            O => \N__38752\,
            I => \N__38748\
        );

    \I__6762\ : InMux
    port map (
            O => \N__38751\,
            I => \N__38745\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__38748\,
            I => control_mode_4
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__38745\,
            I => control_mode_4
        );

    \I__6759\ : InMux
    port map (
            O => \N__38740\,
            I => \N__38737\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__38737\,
            I => \N__38734\
        );

    \I__6757\ : Span4Mux_v
    port map (
            O => \N__38734\,
            I => \N__38730\
        );

    \I__6756\ : InMux
    port map (
            O => \N__38733\,
            I => \N__38727\
        );

    \I__6755\ : Odrv4
    port map (
            O => \N__38730\,
            I => control_mode_3
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__38727\,
            I => control_mode_3
        );

    \I__6753\ : InMux
    port map (
            O => \N__38722\,
            I => \N__38719\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__38719\,
            I => \N__38716\
        );

    \I__6751\ : Sp12to4
    port map (
            O => \N__38716\,
            I => \N__38712\
        );

    \I__6750\ : InMux
    port map (
            O => \N__38715\,
            I => \N__38709\
        );

    \I__6749\ : Odrv12
    port map (
            O => \N__38712\,
            I => control_mode_7
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__38709\,
            I => control_mode_7
        );

    \I__6747\ : CascadeMux
    port map (
            O => \N__38704\,
            I => \c0.n9_cascade_\
        );

    \I__6746\ : CascadeMux
    port map (
            O => \N__38701\,
            I => \c0.n16_adj_3008_cascade_\
        );

    \I__6745\ : InMux
    port map (
            O => \N__38698\,
            I => \N__38695\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__38695\,
            I => \c0.n9\
        );

    \I__6743\ : CascadeMux
    port map (
            O => \N__38692\,
            I => \c0.n19115_cascade_\
        );

    \I__6742\ : CascadeMux
    port map (
            O => \N__38689\,
            I => \N__38685\
        );

    \I__6741\ : InMux
    port map (
            O => \N__38688\,
            I => \N__38682\
        );

    \I__6740\ : InMux
    port map (
            O => \N__38685\,
            I => \N__38679\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__38682\,
            I => \c0.data_in_frame_10_1\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__38679\,
            I => \c0.data_in_frame_10_1\
        );

    \I__6737\ : InMux
    port map (
            O => \N__38674\,
            I => \N__38671\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__38671\,
            I => \N__38666\
        );

    \I__6735\ : InMux
    port map (
            O => \N__38670\,
            I => \N__38663\
        );

    \I__6734\ : InMux
    port map (
            O => \N__38669\,
            I => \N__38660\
        );

    \I__6733\ : Span4Mux_h
    port map (
            O => \N__38666\,
            I => \N__38657\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__38663\,
            I => \N__38654\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__38660\,
            I => \N__38651\
        );

    \I__6730\ : Span4Mux_v
    port map (
            O => \N__38657\,
            I => \N__38648\
        );

    \I__6729\ : Span12Mux_v
    port map (
            O => \N__38654\,
            I => \N__38643\
        );

    \I__6728\ : Span12Mux_h
    port map (
            O => \N__38651\,
            I => \N__38643\
        );

    \I__6727\ : Odrv4
    port map (
            O => \N__38648\,
            I => \c0.n63_adj_3146\
        );

    \I__6726\ : Odrv12
    port map (
            O => \N__38643\,
            I => \c0.n63_adj_3146\
        );

    \I__6725\ : CascadeMux
    port map (
            O => \N__38638\,
            I => \c0.n20_adj_3437_cascade_\
        );

    \I__6724\ : CascadeMux
    port map (
            O => \N__38635\,
            I => \n21222_cascade_\
        );

    \I__6723\ : InMux
    port map (
            O => \N__38632\,
            I => \N__38628\
        );

    \I__6722\ : InMux
    port map (
            O => \N__38631\,
            I => \N__38625\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__38628\,
            I => control_mode_6
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__38625\,
            I => control_mode_6
        );

    \I__6719\ : InMux
    port map (
            O => \N__38620\,
            I => \N__38616\
        );

    \I__6718\ : InMux
    port map (
            O => \N__38619\,
            I => \N__38613\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__38616\,
            I => control_mode_2
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__38613\,
            I => control_mode_2
        );

    \I__6715\ : CascadeMux
    port map (
            O => \N__38608\,
            I => \N__38604\
        );

    \I__6714\ : CascadeMux
    port map (
            O => \N__38607\,
            I => \N__38601\
        );

    \I__6713\ : InMux
    port map (
            O => \N__38604\,
            I => \N__38593\
        );

    \I__6712\ : InMux
    port map (
            O => \N__38601\,
            I => \N__38593\
        );

    \I__6711\ : InMux
    port map (
            O => \N__38600\,
            I => \N__38593\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__38593\,
            I => \c0.data_in_frame_5_0\
        );

    \I__6709\ : CascadeMux
    port map (
            O => \N__38590\,
            I => \N__38586\
        );

    \I__6708\ : CascadeMux
    port map (
            O => \N__38589\,
            I => \N__38583\
        );

    \I__6707\ : InMux
    port map (
            O => \N__38586\,
            I => \N__38578\
        );

    \I__6706\ : InMux
    port map (
            O => \N__38583\,
            I => \N__38578\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__38578\,
            I => \c0.data_in_frame_9_7\
        );

    \I__6704\ : InMux
    port map (
            O => \N__38575\,
            I => \N__38572\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__38572\,
            I => \c0.n38_adj_3328\
        );

    \I__6702\ : CascadeMux
    port map (
            O => \N__38569\,
            I => \c0.n21279_cascade_\
        );

    \I__6701\ : CascadeMux
    port map (
            O => \N__38566\,
            I => \c0.n21255_cascade_\
        );

    \I__6700\ : InMux
    port map (
            O => \N__38563\,
            I => \N__38560\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__38560\,
            I => \c0.n37_adj_3332\
        );

    \I__6698\ : CascadeMux
    port map (
            O => \N__38557\,
            I => \c0.n63_adj_3417_cascade_\
        );

    \I__6697\ : CascadeMux
    port map (
            O => \N__38554\,
            I => \c0.n5_adj_3040_cascade_\
        );

    \I__6696\ : InMux
    port map (
            O => \N__38551\,
            I => \N__38548\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__38548\,
            I => \N__38545\
        );

    \I__6694\ : Odrv4
    port map (
            O => \N__38545\,
            I => \c0.n30_adj_3264\
        );

    \I__6693\ : InMux
    port map (
            O => \N__38542\,
            I => \N__38539\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__38539\,
            I => \c0.n26_adj_3107\
        );

    \I__6691\ : CascadeMux
    port map (
            O => \N__38536\,
            I => \c0.n21281_cascade_\
        );

    \I__6690\ : InMux
    port map (
            O => \N__38533\,
            I => \N__38530\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__38530\,
            I => \c0.n108\
        );

    \I__6688\ : CascadeMux
    port map (
            O => \N__38527\,
            I => \c0.n108_cascade_\
        );

    \I__6687\ : InMux
    port map (
            O => \N__38524\,
            I => \N__38521\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__38521\,
            I => \N__38516\
        );

    \I__6685\ : InMux
    port map (
            O => \N__38520\,
            I => \N__38510\
        );

    \I__6684\ : InMux
    port map (
            O => \N__38519\,
            I => \N__38510\
        );

    \I__6683\ : Span4Mux_h
    port map (
            O => \N__38516\,
            I => \N__38507\
        );

    \I__6682\ : InMux
    port map (
            O => \N__38515\,
            I => \N__38504\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__38510\,
            I => \N__38501\
        );

    \I__6680\ : Odrv4
    port map (
            O => \N__38507\,
            I => \c0.n92_adj_3254\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__38504\,
            I => \c0.n92_adj_3254\
        );

    \I__6678\ : Odrv4
    port map (
            O => \N__38501\,
            I => \c0.n92_adj_3254\
        );

    \I__6677\ : InMux
    port map (
            O => \N__38494\,
            I => \N__38486\
        );

    \I__6676\ : InMux
    port map (
            O => \N__38493\,
            I => \N__38486\
        );

    \I__6675\ : InMux
    port map (
            O => \N__38492\,
            I => \N__38481\
        );

    \I__6674\ : InMux
    port map (
            O => \N__38491\,
            I => \N__38481\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__38486\,
            I => data_in_1_2
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__38481\,
            I => data_in_1_2
        );

    \I__6671\ : InMux
    port map (
            O => \N__38476\,
            I => \N__38473\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__38473\,
            I => \N__38470\
        );

    \I__6669\ : Span4Mux_v
    port map (
            O => \N__38470\,
            I => \N__38466\
        );

    \I__6668\ : InMux
    port map (
            O => \N__38469\,
            I => \N__38463\
        );

    \I__6667\ : Odrv4
    port map (
            O => \N__38466\,
            I => \c0.n121\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__38463\,
            I => \c0.n121\
        );

    \I__6665\ : InMux
    port map (
            O => \N__38458\,
            I => \N__38452\
        );

    \I__6664\ : InMux
    port map (
            O => \N__38457\,
            I => \N__38452\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__38452\,
            I => \c0.n103\
        );

    \I__6662\ : InMux
    port map (
            O => \N__38449\,
            I => \N__38446\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__38446\,
            I => \c0.n63_adj_3084\
        );

    \I__6660\ : InMux
    port map (
            O => \N__38443\,
            I => \N__38440\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__38440\,
            I => \c0.n19_adj_3252\
        );

    \I__6658\ : InMux
    port map (
            O => \N__38437\,
            I => \N__38431\
        );

    \I__6657\ : InMux
    port map (
            O => \N__38436\,
            I => \N__38431\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__38431\,
            I => \c0.n21_adj_3253\
        );

    \I__6655\ : CascadeMux
    port map (
            O => \N__38428\,
            I => \c0.n19_adj_3252_cascade_\
        );

    \I__6654\ : InMux
    port map (
            O => \N__38425\,
            I => \N__38419\
        );

    \I__6653\ : InMux
    port map (
            O => \N__38424\,
            I => \N__38419\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__38419\,
            I => \c0.n63_adj_3083\
        );

    \I__6651\ : InMux
    port map (
            O => \N__38416\,
            I => \N__38408\
        );

    \I__6650\ : InMux
    port map (
            O => \N__38415\,
            I => \N__38408\
        );

    \I__6649\ : InMux
    port map (
            O => \N__38414\,
            I => \N__38403\
        );

    \I__6648\ : InMux
    port map (
            O => \N__38413\,
            I => \N__38403\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__38408\,
            I => \c0.n7804\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__38403\,
            I => \c0.n7804\
        );

    \I__6645\ : InMux
    port map (
            O => \N__38398\,
            I => \N__38395\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__38395\,
            I => \N__38392\
        );

    \I__6643\ : Span12Mux_v
    port map (
            O => \N__38392\,
            I => \N__38389\
        );

    \I__6642\ : Odrv12
    port map (
            O => \N__38389\,
            I => \c0.n11_adj_3093\
        );

    \I__6641\ : CascadeMux
    port map (
            O => \N__38386\,
            I => \c0.n15701_cascade_\
        );

    \I__6640\ : CascadeMux
    port map (
            O => \N__38383\,
            I => \n11421_cascade_\
        );

    \I__6639\ : InMux
    port map (
            O => \N__38380\,
            I => \N__38377\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__38377\,
            I => \N__38374\
        );

    \I__6637\ : Span4Mux_v
    port map (
            O => \N__38374\,
            I => \N__38370\
        );

    \I__6636\ : InMux
    port map (
            O => \N__38373\,
            I => \N__38367\
        );

    \I__6635\ : Odrv4
    port map (
            O => \N__38370\,
            I => \c0.n11422\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__38367\,
            I => \c0.n11422\
        );

    \I__6633\ : InMux
    port map (
            O => \N__38362\,
            I => \N__38358\
        );

    \I__6632\ : InMux
    port map (
            O => \N__38361\,
            I => \N__38355\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__38358\,
            I => \N__38349\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__38355\,
            I => \N__38349\
        );

    \I__6629\ : InMux
    port map (
            O => \N__38354\,
            I => \N__38345\
        );

    \I__6628\ : Span4Mux_v
    port map (
            O => \N__38349\,
            I => \N__38342\
        );

    \I__6627\ : InMux
    port map (
            O => \N__38348\,
            I => \N__38339\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__38345\,
            I => \N__38336\
        );

    \I__6625\ : Span4Mux_h
    port map (
            O => \N__38342\,
            I => \N__38331\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__38339\,
            I => \N__38331\
        );

    \I__6623\ : Odrv4
    port map (
            O => \N__38336\,
            I => \c0.n3632\
        );

    \I__6622\ : Odrv4
    port map (
            O => \N__38331\,
            I => \c0.n3632\
        );

    \I__6621\ : InMux
    port map (
            O => \N__38326\,
            I => \N__38322\
        );

    \I__6620\ : InMux
    port map (
            O => \N__38325\,
            I => \N__38318\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__38322\,
            I => \N__38314\
        );

    \I__6618\ : InMux
    port map (
            O => \N__38321\,
            I => \N__38310\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__38318\,
            I => \N__38307\
        );

    \I__6616\ : InMux
    port map (
            O => \N__38317\,
            I => \N__38304\
        );

    \I__6615\ : Span4Mux_v
    port map (
            O => \N__38314\,
            I => \N__38301\
        );

    \I__6614\ : InMux
    port map (
            O => \N__38313\,
            I => \N__38298\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__38310\,
            I => \N__38293\
        );

    \I__6612\ : Span4Mux_v
    port map (
            O => \N__38307\,
            I => \N__38293\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__38304\,
            I => \c0.n9389\
        );

    \I__6610\ : Odrv4
    port map (
            O => \N__38301\,
            I => \c0.n9389\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__38298\,
            I => \c0.n9389\
        );

    \I__6608\ : Odrv4
    port map (
            O => \N__38293\,
            I => \c0.n9389\
        );

    \I__6607\ : InMux
    port map (
            O => \N__38284\,
            I => \N__38281\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__38281\,
            I => \N__38278\
        );

    \I__6605\ : Span4Mux_h
    port map (
            O => \N__38278\,
            I => \N__38274\
        );

    \I__6604\ : InMux
    port map (
            O => \N__38277\,
            I => \N__38271\
        );

    \I__6603\ : Odrv4
    port map (
            O => \N__38274\,
            I => \c0.n3\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__38271\,
            I => \c0.n3\
        );

    \I__6601\ : InMux
    port map (
            O => \N__38266\,
            I => \N__38262\
        );

    \I__6600\ : InMux
    port map (
            O => \N__38265\,
            I => \N__38259\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__38262\,
            I => \N__38255\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__38259\,
            I => \N__38252\
        );

    \I__6597\ : InMux
    port map (
            O => \N__38258\,
            I => \N__38249\
        );

    \I__6596\ : Span4Mux_v
    port map (
            O => \N__38255\,
            I => \N__38238\
        );

    \I__6595\ : Span4Mux_h
    port map (
            O => \N__38252\,
            I => \N__38238\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__38249\,
            I => \N__38238\
        );

    \I__6593\ : InMux
    port map (
            O => \N__38248\,
            I => \N__38235\
        );

    \I__6592\ : InMux
    port map (
            O => \N__38247\,
            I => \N__38230\
        );

    \I__6591\ : InMux
    port map (
            O => \N__38246\,
            I => \N__38230\
        );

    \I__6590\ : InMux
    port map (
            O => \N__38245\,
            I => \N__38227\
        );

    \I__6589\ : Span4Mux_h
    port map (
            O => \N__38238\,
            I => \N__38224\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__38235\,
            I => \N__38221\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__38230\,
            I => \c0.n11427\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__38227\,
            I => \c0.n11427\
        );

    \I__6585\ : Odrv4
    port map (
            O => \N__38224\,
            I => \c0.n11427\
        );

    \I__6584\ : Odrv12
    port map (
            O => \N__38221\,
            I => \c0.n11427\
        );

    \I__6583\ : InMux
    port map (
            O => \N__38212\,
            I => \N__38208\
        );

    \I__6582\ : InMux
    port map (
            O => \N__38211\,
            I => \N__38205\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__38208\,
            I => \c0.n15874\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__38205\,
            I => \c0.n15874\
        );

    \I__6579\ : InMux
    port map (
            O => \N__38200\,
            I => \N__38197\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__38197\,
            I => n12917
        );

    \I__6577\ : InMux
    port map (
            O => \N__38194\,
            I => \N__38190\
        );

    \I__6576\ : InMux
    port map (
            O => \N__38193\,
            I => \N__38187\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__38190\,
            I => \N__38181\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__38187\,
            I => \N__38181\
        );

    \I__6573\ : InMux
    port map (
            O => \N__38186\,
            I => \N__38178\
        );

    \I__6572\ : Span4Mux_h
    port map (
            O => \N__38181\,
            I => \N__38175\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__38178\,
            I => \c0.n11440\
        );

    \I__6570\ : Odrv4
    port map (
            O => \N__38175\,
            I => \c0.n11440\
        );

    \I__6569\ : CascadeMux
    port map (
            O => \N__38170\,
            I => \c0.n11317_cascade_\
        );

    \I__6568\ : CascadeMux
    port map (
            O => \N__38167\,
            I => \N__38164\
        );

    \I__6567\ : InMux
    port map (
            O => \N__38164\,
            I => \N__38161\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__38161\,
            I => \N__38157\
        );

    \I__6565\ : InMux
    port map (
            O => \N__38160\,
            I => \N__38154\
        );

    \I__6564\ : Span4Mux_v
    port map (
            O => \N__38157\,
            I => \N__38150\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__38154\,
            I => \N__38147\
        );

    \I__6562\ : InMux
    port map (
            O => \N__38153\,
            I => \N__38144\
        );

    \I__6561\ : Span4Mux_v
    port map (
            O => \N__38150\,
            I => \N__38141\
        );

    \I__6560\ : Span4Mux_h
    port map (
            O => \N__38147\,
            I => \N__38136\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__38144\,
            I => \N__38136\
        );

    \I__6558\ : Span4Mux_v
    port map (
            O => \N__38141\,
            I => \N__38131\
        );

    \I__6557\ : Sp12to4
    port map (
            O => \N__38136\,
            I => \N__38128\
        );

    \I__6556\ : InMux
    port map (
            O => \N__38135\,
            I => \N__38125\
        );

    \I__6555\ : InMux
    port map (
            O => \N__38134\,
            I => \N__38122\
        );

    \I__6554\ : Span4Mux_v
    port map (
            O => \N__38131\,
            I => \N__38119\
        );

    \I__6553\ : Span12Mux_v
    port map (
            O => \N__38128\,
            I => \N__38116\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__38125\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__38122\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__6550\ : Odrv4
    port map (
            O => \N__38119\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__6549\ : Odrv12
    port map (
            O => \N__38116\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__6548\ : InMux
    port map (
            O => \N__38107\,
            I => \N__38101\
        );

    \I__6547\ : InMux
    port map (
            O => \N__38106\,
            I => \N__38098\
        );

    \I__6546\ : InMux
    port map (
            O => \N__38105\,
            I => \N__38095\
        );

    \I__6545\ : InMux
    port map (
            O => \N__38104\,
            I => \N__38092\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__38101\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__38098\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__38095\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__38092\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__6540\ : InMux
    port map (
            O => \N__38083\,
            I => \N__38077\
        );

    \I__6539\ : InMux
    port map (
            O => \N__38082\,
            I => \N__38074\
        );

    \I__6538\ : InMux
    port map (
            O => \N__38081\,
            I => \N__38071\
        );

    \I__6537\ : InMux
    port map (
            O => \N__38080\,
            I => \N__38068\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__38077\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__38074\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__38071\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__38068\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__6532\ : InMux
    port map (
            O => \N__38059\,
            I => \N__38056\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__38056\,
            I => \N__38053\
        );

    \I__6530\ : Odrv4
    port map (
            O => \N__38053\,
            I => \c0.rx.n21267\
        );

    \I__6529\ : InMux
    port map (
            O => \N__38050\,
            I => \N__38047\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__38047\,
            I => \N__38042\
        );

    \I__6527\ : InMux
    port map (
            O => \N__38046\,
            I => \N__38039\
        );

    \I__6526\ : InMux
    port map (
            O => \N__38045\,
            I => \N__38036\
        );

    \I__6525\ : Span4Mux_h
    port map (
            O => \N__38042\,
            I => \N__38033\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__38039\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__38036\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__6522\ : Odrv4
    port map (
            O => \N__38033\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__6521\ : CascadeMux
    port map (
            O => \N__38026\,
            I => \N__38023\
        );

    \I__6520\ : InMux
    port map (
            O => \N__38023\,
            I => \N__38020\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__38020\,
            I => \N__38015\
        );

    \I__6518\ : InMux
    port map (
            O => \N__38019\,
            I => \N__38012\
        );

    \I__6517\ : InMux
    port map (
            O => \N__38018\,
            I => \N__38009\
        );

    \I__6516\ : Span4Mux_h
    port map (
            O => \N__38015\,
            I => \N__38006\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__38012\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__38009\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__6513\ : Odrv4
    port map (
            O => \N__38006\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__6512\ : InMux
    port map (
            O => \N__37999\,
            I => \N__37996\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__37996\,
            I => \N__37993\
        );

    \I__6510\ : Span4Mux_v
    port map (
            O => \N__37993\,
            I => \N__37989\
        );

    \I__6509\ : InMux
    port map (
            O => \N__37992\,
            I => \N__37986\
        );

    \I__6508\ : Span4Mux_v
    port map (
            O => \N__37989\,
            I => \N__37982\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__37986\,
            I => \N__37979\
        );

    \I__6506\ : InMux
    port map (
            O => \N__37985\,
            I => \N__37976\
        );

    \I__6505\ : Span4Mux_v
    port map (
            O => \N__37982\,
            I => \N__37973\
        );

    \I__6504\ : Odrv4
    port map (
            O => \N__37979\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__37976\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__6502\ : Odrv4
    port map (
            O => \N__37973\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__6501\ : InMux
    port map (
            O => \N__37966\,
            I => \N__37963\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__37963\,
            I => \c0.n42_adj_3256\
        );

    \I__6499\ : InMux
    port map (
            O => \N__37960\,
            I => \N__37956\
        );

    \I__6498\ : InMux
    port map (
            O => \N__37959\,
            I => \N__37953\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__37956\,
            I => \N__37950\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__37953\,
            I => \N__37947\
        );

    \I__6495\ : Odrv4
    port map (
            O => \N__37950\,
            I => \c0.n1_adj_3002\
        );

    \I__6494\ : Odrv4
    port map (
            O => \N__37947\,
            I => \c0.n1_adj_3002\
        );

    \I__6493\ : InMux
    port map (
            O => \N__37942\,
            I => \N__37939\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__37939\,
            I => \N__37936\
        );

    \I__6491\ : Odrv12
    port map (
            O => \N__37936\,
            I => \c0.n21053\
        );

    \I__6490\ : CascadeMux
    port map (
            O => \N__37933\,
            I => \c0.rx.n35_cascade_\
        );

    \I__6489\ : CascadeMux
    port map (
            O => \N__37930\,
            I => \N__37924\
        );

    \I__6488\ : CascadeMux
    port map (
            O => \N__37929\,
            I => \N__37917\
        );

    \I__6487\ : InMux
    port map (
            O => \N__37928\,
            I => \N__37914\
        );

    \I__6486\ : InMux
    port map (
            O => \N__37927\,
            I => \N__37907\
        );

    \I__6485\ : InMux
    port map (
            O => \N__37924\,
            I => \N__37907\
        );

    \I__6484\ : InMux
    port map (
            O => \N__37923\,
            I => \N__37900\
        );

    \I__6483\ : InMux
    port map (
            O => \N__37922\,
            I => \N__37900\
        );

    \I__6482\ : InMux
    port map (
            O => \N__37921\,
            I => \N__37900\
        );

    \I__6481\ : InMux
    port map (
            O => \N__37920\,
            I => \N__37895\
        );

    \I__6480\ : InMux
    port map (
            O => \N__37917\,
            I => \N__37895\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__37914\,
            I => \N__37892\
        );

    \I__6478\ : InMux
    port map (
            O => \N__37913\,
            I => \N__37887\
        );

    \I__6477\ : InMux
    port map (
            O => \N__37912\,
            I => \N__37887\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__37907\,
            I => \N__37884\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__37900\,
            I => \r_SM_Main_0\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__37895\,
            I => \r_SM_Main_0\
        );

    \I__6473\ : Odrv4
    port map (
            O => \N__37892\,
            I => \r_SM_Main_0\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__37887\,
            I => \r_SM_Main_0\
        );

    \I__6471\ : Odrv4
    port map (
            O => \N__37884\,
            I => \r_SM_Main_0\
        );

    \I__6470\ : CascadeMux
    port map (
            O => \N__37873\,
            I => \c0.rx.n12_cascade_\
        );

    \I__6469\ : InMux
    port map (
            O => \N__37870\,
            I => \N__37867\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__37867\,
            I => \N__37864\
        );

    \I__6467\ : Span4Mux_h
    port map (
            O => \N__37864\,
            I => \N__37859\
        );

    \I__6466\ : InMux
    port map (
            O => \N__37863\,
            I => \N__37854\
        );

    \I__6465\ : InMux
    port map (
            O => \N__37862\,
            I => \N__37846\
        );

    \I__6464\ : Span4Mux_v
    port map (
            O => \N__37859\,
            I => \N__37843\
        );

    \I__6463\ : InMux
    port map (
            O => \N__37858\,
            I => \N__37838\
        );

    \I__6462\ : InMux
    port map (
            O => \N__37857\,
            I => \N__37838\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__37854\,
            I => \N__37835\
        );

    \I__6460\ : InMux
    port map (
            O => \N__37853\,
            I => \N__37828\
        );

    \I__6459\ : InMux
    port map (
            O => \N__37852\,
            I => \N__37828\
        );

    \I__6458\ : InMux
    port map (
            O => \N__37851\,
            I => \N__37828\
        );

    \I__6457\ : InMux
    port map (
            O => \N__37850\,
            I => \N__37823\
        );

    \I__6456\ : InMux
    port map (
            O => \N__37849\,
            I => \N__37823\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__37846\,
            I => \r_SM_Main_1\
        );

    \I__6454\ : Odrv4
    port map (
            O => \N__37843\,
            I => \r_SM_Main_1\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__37838\,
            I => \r_SM_Main_1\
        );

    \I__6452\ : Odrv4
    port map (
            O => \N__37835\,
            I => \r_SM_Main_1\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__37828\,
            I => \r_SM_Main_1\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__37823\,
            I => \r_SM_Main_1\
        );

    \I__6449\ : InMux
    port map (
            O => \N__37810\,
            I => \N__37807\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__37807\,
            I => \N__37802\
        );

    \I__6447\ : InMux
    port map (
            O => \N__37806\,
            I => \N__37791\
        );

    \I__6446\ : InMux
    port map (
            O => \N__37805\,
            I => \N__37791\
        );

    \I__6445\ : Sp12to4
    port map (
            O => \N__37802\,
            I => \N__37788\
        );

    \I__6444\ : InMux
    port map (
            O => \N__37801\,
            I => \N__37785\
        );

    \I__6443\ : InMux
    port map (
            O => \N__37800\,
            I => \N__37780\
        );

    \I__6442\ : InMux
    port map (
            O => \N__37799\,
            I => \N__37780\
        );

    \I__6441\ : InMux
    port map (
            O => \N__37798\,
            I => \N__37777\
        );

    \I__6440\ : InMux
    port map (
            O => \N__37797\,
            I => \N__37772\
        );

    \I__6439\ : InMux
    port map (
            O => \N__37796\,
            I => \N__37772\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__37791\,
            I => \N__37769\
        );

    \I__6437\ : Odrv12
    port map (
            O => \N__37788\,
            I => \r_SM_Main_2\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__37785\,
            I => \r_SM_Main_2\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__37780\,
            I => \r_SM_Main_2\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__37777\,
            I => \r_SM_Main_2\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__37772\,
            I => \r_SM_Main_2\
        );

    \I__6432\ : Odrv4
    port map (
            O => \N__37769\,
            I => \r_SM_Main_2\
        );

    \I__6431\ : CascadeMux
    port map (
            O => \N__37756\,
            I => \c0.rx.n21406_cascade_\
        );

    \I__6430\ : CascadeMux
    port map (
            O => \N__37753\,
            I => \N__37750\
        );

    \I__6429\ : InMux
    port map (
            O => \N__37750\,
            I => \N__37745\
        );

    \I__6428\ : InMux
    port map (
            O => \N__37749\,
            I => \N__37741\
        );

    \I__6427\ : InMux
    port map (
            O => \N__37748\,
            I => \N__37738\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__37745\,
            I => \N__37735\
        );

    \I__6425\ : InMux
    port map (
            O => \N__37744\,
            I => \N__37732\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__37741\,
            I => \r_SM_Main_2_N_2473_2\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__37738\,
            I => \r_SM_Main_2_N_2473_2\
        );

    \I__6422\ : Odrv4
    port map (
            O => \N__37735\,
            I => \r_SM_Main_2_N_2473_2\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__37732\,
            I => \r_SM_Main_2_N_2473_2\
        );

    \I__6420\ : InMux
    port map (
            O => \N__37723\,
            I => \N__37719\
        );

    \I__6419\ : InMux
    port map (
            O => \N__37722\,
            I => \N__37716\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__37719\,
            I => \N__37710\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__37716\,
            I => \N__37707\
        );

    \I__6416\ : InMux
    port map (
            O => \N__37715\,
            I => \N__37704\
        );

    \I__6415\ : InMux
    port map (
            O => \N__37714\,
            I => \N__37699\
        );

    \I__6414\ : InMux
    port map (
            O => \N__37713\,
            I => \N__37699\
        );

    \I__6413\ : Sp12to4
    port map (
            O => \N__37710\,
            I => \N__37690\
        );

    \I__6412\ : Sp12to4
    port map (
            O => \N__37707\,
            I => \N__37690\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__37704\,
            I => \N__37690\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__37699\,
            I => \N__37690\
        );

    \I__6409\ : Odrv12
    port map (
            O => \N__37690\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__6408\ : InMux
    port map (
            O => \N__37687\,
            I => \N__37684\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__37684\,
            I => \N__37676\
        );

    \I__6406\ : InMux
    port map (
            O => \N__37683\,
            I => \N__37673\
        );

    \I__6405\ : InMux
    port map (
            O => \N__37682\,
            I => \N__37670\
        );

    \I__6404\ : InMux
    port map (
            O => \N__37681\,
            I => \N__37663\
        );

    \I__6403\ : InMux
    port map (
            O => \N__37680\,
            I => \N__37663\
        );

    \I__6402\ : InMux
    port map (
            O => \N__37679\,
            I => \N__37663\
        );

    \I__6401\ : Odrv4
    port map (
            O => \N__37676\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__37673\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__37670\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__37663\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__6397\ : InMux
    port map (
            O => \N__37654\,
            I => \N__37649\
        );

    \I__6396\ : CascadeMux
    port map (
            O => \N__37653\,
            I => \N__37644\
        );

    \I__6395\ : InMux
    port map (
            O => \N__37652\,
            I => \N__37641\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__37649\,
            I => \N__37638\
        );

    \I__6393\ : InMux
    port map (
            O => \N__37648\,
            I => \N__37633\
        );

    \I__6392\ : InMux
    port map (
            O => \N__37647\,
            I => \N__37633\
        );

    \I__6391\ : InMux
    port map (
            O => \N__37644\,
            I => \N__37630\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__37641\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__6389\ : Odrv4
    port map (
            O => \N__37638\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__37633\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__37630\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__6386\ : InMux
    port map (
            O => \N__37621\,
            I => \N__37618\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__37618\,
            I => \N__37614\
        );

    \I__6384\ : InMux
    port map (
            O => \N__37617\,
            I => \N__37611\
        );

    \I__6383\ : Span4Mux_h
    port map (
            O => \N__37614\,
            I => \N__37603\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__37611\,
            I => \N__37603\
        );

    \I__6381\ : InMux
    port map (
            O => \N__37610\,
            I => \N__37600\
        );

    \I__6380\ : InMux
    port map (
            O => \N__37609\,
            I => \N__37595\
        );

    \I__6379\ : InMux
    port map (
            O => \N__37608\,
            I => \N__37595\
        );

    \I__6378\ : Sp12to4
    port map (
            O => \N__37603\,
            I => \N__37588\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__37600\,
            I => \N__37588\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__37595\,
            I => \N__37588\
        );

    \I__6375\ : Odrv12
    port map (
            O => \N__37588\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__6374\ : InMux
    port map (
            O => \N__37585\,
            I => \N__37582\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__37582\,
            I => \c0.rx.n8\
        );

    \I__6372\ : InMux
    port map (
            O => \N__37579\,
            I => \N__37576\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__37576\,
            I => n12914
        );

    \I__6370\ : CascadeMux
    port map (
            O => \N__37573\,
            I => \c0.rx.n15906_cascade_\
        );

    \I__6369\ : InMux
    port map (
            O => \N__37570\,
            I => \N__37567\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__37567\,
            I => \c0.rx.n20851\
        );

    \I__6367\ : CascadeMux
    port map (
            O => \N__37564\,
            I => \N__37561\
        );

    \I__6366\ : InMux
    port map (
            O => \N__37561\,
            I => \N__37558\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__37558\,
            I => \c0.rx.n32\
        );

    \I__6364\ : SRMux
    port map (
            O => \N__37555\,
            I => \N__37552\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__37552\,
            I => \c0.rx.n20964\
        );

    \I__6362\ : InMux
    port map (
            O => \N__37549\,
            I => \N__37543\
        );

    \I__6361\ : InMux
    port map (
            O => \N__37548\,
            I => \N__37543\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__37543\,
            I => \c0.rx.n15906\
        );

    \I__6359\ : CascadeMux
    port map (
            O => \N__37540\,
            I => \r_SM_Main_2_N_2473_2_cascade_\
        );

    \I__6358\ : InMux
    port map (
            O => \N__37537\,
            I => \N__37534\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__37534\,
            I => \c0.rx.n15926\
        );

    \I__6356\ : InMux
    port map (
            O => \N__37531\,
            I => \N__37528\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__37528\,
            I => n9
        );

    \I__6354\ : InMux
    port map (
            O => \N__37525\,
            I => \N__37519\
        );

    \I__6353\ : InMux
    port map (
            O => \N__37524\,
            I => \N__37516\
        );

    \I__6352\ : InMux
    port map (
            O => \N__37523\,
            I => \N__37511\
        );

    \I__6351\ : InMux
    port map (
            O => \N__37522\,
            I => \N__37511\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__37519\,
            I => \N__37506\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__37516\,
            I => \N__37506\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__37511\,
            I => \N__37503\
        );

    \I__6347\ : Odrv12
    port map (
            O => \N__37506\,
            I => \c0.n9755\
        );

    \I__6346\ : Odrv4
    port map (
            O => \N__37503\,
            I => \c0.n9755\
        );

    \I__6345\ : CascadeMux
    port map (
            O => \N__37498\,
            I => \N__37495\
        );

    \I__6344\ : InMux
    port map (
            O => \N__37495\,
            I => \N__37492\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__37492\,
            I => \N__37489\
        );

    \I__6342\ : Span4Mux_h
    port map (
            O => \N__37489\,
            I => \N__37485\
        );

    \I__6341\ : InMux
    port map (
            O => \N__37488\,
            I => \N__37482\
        );

    \I__6340\ : Span4Mux_v
    port map (
            O => \N__37485\,
            I => \N__37479\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__37482\,
            I => data_out_frame_28_5
        );

    \I__6338\ : Odrv4
    port map (
            O => \N__37479\,
            I => data_out_frame_28_5
        );

    \I__6337\ : InMux
    port map (
            O => \N__37474\,
            I => \N__37471\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__37471\,
            I => \c0.n21308\
        );

    \I__6335\ : InMux
    port map (
            O => \N__37468\,
            I => \N__37455\
        );

    \I__6334\ : InMux
    port map (
            O => \N__37467\,
            I => \N__37455\
        );

    \I__6333\ : InMux
    port map (
            O => \N__37466\,
            I => \N__37452\
        );

    \I__6332\ : CascadeMux
    port map (
            O => \N__37465\,
            I => \N__37447\
        );

    \I__6331\ : InMux
    port map (
            O => \N__37464\,
            I => \N__37444\
        );

    \I__6330\ : InMux
    port map (
            O => \N__37463\,
            I => \N__37434\
        );

    \I__6329\ : InMux
    port map (
            O => \N__37462\,
            I => \N__37434\
        );

    \I__6328\ : InMux
    port map (
            O => \N__37461\,
            I => \N__37434\
        );

    \I__6327\ : InMux
    port map (
            O => \N__37460\,
            I => \N__37434\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__37455\,
            I => \N__37429\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__37452\,
            I => \N__37429\
        );

    \I__6324\ : CascadeMux
    port map (
            O => \N__37451\,
            I => \N__37425\
        );

    \I__6323\ : InMux
    port map (
            O => \N__37450\,
            I => \N__37419\
        );

    \I__6322\ : InMux
    port map (
            O => \N__37447\,
            I => \N__37416\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__37444\,
            I => \N__37413\
        );

    \I__6320\ : CascadeMux
    port map (
            O => \N__37443\,
            I => \N__37409\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__37434\,
            I => \N__37405\
        );

    \I__6318\ : Sp12to4
    port map (
            O => \N__37429\,
            I => \N__37402\
        );

    \I__6317\ : InMux
    port map (
            O => \N__37428\,
            I => \N__37391\
        );

    \I__6316\ : InMux
    port map (
            O => \N__37425\,
            I => \N__37391\
        );

    \I__6315\ : InMux
    port map (
            O => \N__37424\,
            I => \N__37391\
        );

    \I__6314\ : InMux
    port map (
            O => \N__37423\,
            I => \N__37391\
        );

    \I__6313\ : InMux
    port map (
            O => \N__37422\,
            I => \N__37391\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__37419\,
            I => \N__37388\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__37416\,
            I => \N__37385\
        );

    \I__6310\ : Span4Mux_v
    port map (
            O => \N__37413\,
            I => \N__37382\
        );

    \I__6309\ : InMux
    port map (
            O => \N__37412\,
            I => \N__37379\
        );

    \I__6308\ : InMux
    port map (
            O => \N__37409\,
            I => \N__37376\
        );

    \I__6307\ : InMux
    port map (
            O => \N__37408\,
            I => \N__37373\
        );

    \I__6306\ : Span4Mux_h
    port map (
            O => \N__37405\,
            I => \N__37370\
        );

    \I__6305\ : Span12Mux_v
    port map (
            O => \N__37402\,
            I => \N__37367\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__37391\,
            I => \N__37356\
        );

    \I__6303\ : Span4Mux_v
    port map (
            O => \N__37388\,
            I => \N__37356\
        );

    \I__6302\ : Span4Mux_h
    port map (
            O => \N__37385\,
            I => \N__37356\
        );

    \I__6301\ : Span4Mux_h
    port map (
            O => \N__37382\,
            I => \N__37356\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__37379\,
            I => \N__37356\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__37376\,
            I => byte_transmit_counter_4
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__37373\,
            I => byte_transmit_counter_4
        );

    \I__6297\ : Odrv4
    port map (
            O => \N__37370\,
            I => byte_transmit_counter_4
        );

    \I__6296\ : Odrv12
    port map (
            O => \N__37367\,
            I => byte_transmit_counter_4
        );

    \I__6295\ : Odrv4
    port map (
            O => \N__37356\,
            I => byte_transmit_counter_4
        );

    \I__6294\ : InMux
    port map (
            O => \N__37345\,
            I => \N__37337\
        );

    \I__6293\ : InMux
    port map (
            O => \N__37344\,
            I => \N__37330\
        );

    \I__6292\ : InMux
    port map (
            O => \N__37343\,
            I => \N__37330\
        );

    \I__6291\ : InMux
    port map (
            O => \N__37342\,
            I => \N__37323\
        );

    \I__6290\ : InMux
    port map (
            O => \N__37341\,
            I => \N__37323\
        );

    \I__6289\ : InMux
    port map (
            O => \N__37340\,
            I => \N__37323\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__37337\,
            I => \N__37320\
        );

    \I__6287\ : InMux
    port map (
            O => \N__37336\,
            I => \N__37317\
        );

    \I__6286\ : CascadeMux
    port map (
            O => \N__37335\,
            I => \N__37313\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__37330\,
            I => \N__37308\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__37323\,
            I => \N__37305\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__37320\,
            I => \N__37302\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__37317\,
            I => \N__37298\
        );

    \I__6281\ : InMux
    port map (
            O => \N__37316\,
            I => \N__37295\
        );

    \I__6280\ : InMux
    port map (
            O => \N__37313\,
            I => \N__37292\
        );

    \I__6279\ : InMux
    port map (
            O => \N__37312\,
            I => \N__37289\
        );

    \I__6278\ : InMux
    port map (
            O => \N__37311\,
            I => \N__37286\
        );

    \I__6277\ : Span4Mux_v
    port map (
            O => \N__37308\,
            I => \N__37283\
        );

    \I__6276\ : Span4Mux_h
    port map (
            O => \N__37305\,
            I => \N__37278\
        );

    \I__6275\ : Span4Mux_v
    port map (
            O => \N__37302\,
            I => \N__37278\
        );

    \I__6274\ : InMux
    port map (
            O => \N__37301\,
            I => \N__37275\
        );

    \I__6273\ : Span4Mux_v
    port map (
            O => \N__37298\,
            I => \N__37268\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__37295\,
            I => \N__37268\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__37292\,
            I => \N__37268\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__37289\,
            I => byte_transmit_counter_3
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__37286\,
            I => byte_transmit_counter_3
        );

    \I__6268\ : Odrv4
    port map (
            O => \N__37283\,
            I => byte_transmit_counter_3
        );

    \I__6267\ : Odrv4
    port map (
            O => \N__37278\,
            I => byte_transmit_counter_3
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__37275\,
            I => byte_transmit_counter_3
        );

    \I__6265\ : Odrv4
    port map (
            O => \N__37268\,
            I => byte_transmit_counter_3
        );

    \I__6264\ : CascadeMux
    port map (
            O => \N__37255\,
            I => \c0.n21310_cascade_\
        );

    \I__6263\ : InMux
    port map (
            O => \N__37252\,
            I => \N__37249\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__37249\,
            I => \N__37246\
        );

    \I__6261\ : Odrv12
    port map (
            O => \N__37246\,
            I => \c0.n21568\
        );

    \I__6260\ : InMux
    port map (
            O => \N__37243\,
            I => \N__37240\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__37240\,
            I => \N__37237\
        );

    \I__6258\ : Span4Mux_v
    port map (
            O => \N__37237\,
            I => \N__37234\
        );

    \I__6257\ : Odrv4
    port map (
            O => \N__37234\,
            I => n9_adj_3590
        );

    \I__6256\ : InMux
    port map (
            O => \N__37231\,
            I => \N__37228\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__37228\,
            I => \N__37225\
        );

    \I__6254\ : Span4Mux_v
    port map (
            O => \N__37225\,
            I => \N__37222\
        );

    \I__6253\ : Odrv4
    port map (
            O => \N__37222\,
            I => \c0.rx.n11302\
        );

    \I__6252\ : CascadeMux
    port map (
            O => \N__37219\,
            I => \c0.rx.n11302_cascade_\
        );

    \I__6251\ : InMux
    port map (
            O => \N__37216\,
            I => \N__37213\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__37213\,
            I => \N__37208\
        );

    \I__6249\ : CascadeMux
    port map (
            O => \N__37212\,
            I => \N__37205\
        );

    \I__6248\ : InMux
    port map (
            O => \N__37211\,
            I => \N__37202\
        );

    \I__6247\ : Span4Mux_h
    port map (
            O => \N__37208\,
            I => \N__37199\
        );

    \I__6246\ : InMux
    port map (
            O => \N__37205\,
            I => \N__37196\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__37202\,
            I => \N__37191\
        );

    \I__6244\ : Span4Mux_v
    port map (
            O => \N__37199\,
            I => \N__37191\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__37196\,
            I => \N__37188\
        );

    \I__6242\ : Odrv4
    port map (
            O => \N__37191\,
            I => encoder1_position_0
        );

    \I__6241\ : Odrv12
    port map (
            O => \N__37188\,
            I => encoder1_position_0
        );

    \I__6240\ : InMux
    port map (
            O => \N__37183\,
            I => \N__37179\
        );

    \I__6239\ : InMux
    port map (
            O => \N__37182\,
            I => \N__37176\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__37179\,
            I => \N__37173\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__37176\,
            I => data_out_frame_13_0
        );

    \I__6236\ : Odrv12
    port map (
            O => \N__37173\,
            I => data_out_frame_13_0
        );

    \I__6235\ : CascadeMux
    port map (
            O => \N__37168\,
            I => \c0.rx.n21451_cascade_\
        );

    \I__6234\ : InMux
    port map (
            O => \N__37165\,
            I => \N__37162\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__37162\,
            I => \N__37159\
        );

    \I__6232\ : Span4Mux_v
    port map (
            O => \N__37159\,
            I => \N__37156\
        );

    \I__6231\ : Odrv4
    port map (
            O => \N__37156\,
            I => n12920
        );

    \I__6230\ : InMux
    port map (
            O => \N__37153\,
            I => \N__37150\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__37150\,
            I => \N__37146\
        );

    \I__6228\ : InMux
    port map (
            O => \N__37149\,
            I => \N__37143\
        );

    \I__6227\ : Span12Mux_h
    port map (
            O => \N__37146\,
            I => \N__37138\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__37143\,
            I => \N__37138\
        );

    \I__6225\ : Odrv12
    port map (
            O => \N__37138\,
            I => \c0.n70\
        );

    \I__6224\ : InMux
    port map (
            O => \N__37135\,
            I => \N__37132\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__37132\,
            I => \N__37129\
        );

    \I__6222\ : Span4Mux_v
    port map (
            O => \N__37129\,
            I => \N__37125\
        );

    \I__6221\ : InMux
    port map (
            O => \N__37128\,
            I => \N__37122\
        );

    \I__6220\ : Span4Mux_v
    port map (
            O => \N__37125\,
            I => \N__37119\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__37122\,
            I => \N__37116\
        );

    \I__6218\ : Odrv4
    port map (
            O => \N__37119\,
            I => \c0.n15850\
        );

    \I__6217\ : Odrv4
    port map (
            O => \N__37116\,
            I => \c0.n15850\
        );

    \I__6216\ : CascadeMux
    port map (
            O => \N__37111\,
            I => \N__37108\
        );

    \I__6215\ : InMux
    port map (
            O => \N__37108\,
            I => \N__37105\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__37105\,
            I => \N__37102\
        );

    \I__6213\ : Span4Mux_v
    port map (
            O => \N__37102\,
            I => \N__37099\
        );

    \I__6212\ : Span4Mux_h
    port map (
            O => \N__37099\,
            I => \N__37096\
        );

    \I__6211\ : Odrv4
    port map (
            O => \N__37096\,
            I => \c0.n21231\
        );

    \I__6210\ : CascadeMux
    port map (
            O => \N__37093\,
            I => \N__37088\
        );

    \I__6209\ : CascadeMux
    port map (
            O => \N__37092\,
            I => \N__37085\
        );

    \I__6208\ : InMux
    port map (
            O => \N__37091\,
            I => \N__37082\
        );

    \I__6207\ : InMux
    port map (
            O => \N__37088\,
            I => \N__37077\
        );

    \I__6206\ : InMux
    port map (
            O => \N__37085\,
            I => \N__37077\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__37082\,
            I => \N__37074\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__37077\,
            I => \N__37071\
        );

    \I__6203\ : Span4Mux_h
    port map (
            O => \N__37074\,
            I => \N__37068\
        );

    \I__6202\ : Span4Mux_h
    port map (
            O => \N__37071\,
            I => \N__37065\
        );

    \I__6201\ : Odrv4
    port map (
            O => \N__37068\,
            I => \c0.n12254\
        );

    \I__6200\ : Odrv4
    port map (
            O => \N__37065\,
            I => \c0.n12254\
        );

    \I__6199\ : CascadeMux
    port map (
            O => \N__37060\,
            I => \N__37056\
        );

    \I__6198\ : InMux
    port map (
            O => \N__37059\,
            I => \N__37053\
        );

    \I__6197\ : InMux
    port map (
            O => \N__37056\,
            I => \N__37050\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__37053\,
            I => \N__37047\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__37050\,
            I => \N__37043\
        );

    \I__6194\ : Sp12to4
    port map (
            O => \N__37047\,
            I => \N__37040\
        );

    \I__6193\ : InMux
    port map (
            O => \N__37046\,
            I => \N__37037\
        );

    \I__6192\ : Span4Mux_h
    port map (
            O => \N__37043\,
            I => \N__37034\
        );

    \I__6191\ : Odrv12
    port map (
            O => \N__37040\,
            I => encoder1_position_12
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__37037\,
            I => encoder1_position_12
        );

    \I__6189\ : Odrv4
    port map (
            O => \N__37034\,
            I => encoder1_position_12
        );

    \I__6188\ : InMux
    port map (
            O => \N__37027\,
            I => \N__37024\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__37024\,
            I => \N__37020\
        );

    \I__6186\ : InMux
    port map (
            O => \N__37023\,
            I => \N__37017\
        );

    \I__6185\ : Span4Mux_v
    port map (
            O => \N__37020\,
            I => \N__37014\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__37017\,
            I => \N__37009\
        );

    \I__6183\ : Span4Mux_h
    port map (
            O => \N__37014\,
            I => \N__37009\
        );

    \I__6182\ : Odrv4
    port map (
            O => \N__37009\,
            I => data_out_frame_12_4
        );

    \I__6181\ : InMux
    port map (
            O => \N__37006\,
            I => \N__37002\
        );

    \I__6180\ : InMux
    port map (
            O => \N__37005\,
            I => \N__36999\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__37002\,
            I => data_out_frame_5_7
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__36999\,
            I => data_out_frame_5_7
        );

    \I__6177\ : InMux
    port map (
            O => \N__36994\,
            I => \N__36991\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__36991\,
            I => \c0.n5_adj_3475\
        );

    \I__6175\ : CascadeMux
    port map (
            O => \N__36988\,
            I => \N__36983\
        );

    \I__6174\ : CascadeMux
    port map (
            O => \N__36987\,
            I => \N__36980\
        );

    \I__6173\ : CascadeMux
    port map (
            O => \N__36986\,
            I => \N__36977\
        );

    \I__6172\ : InMux
    port map (
            O => \N__36983\,
            I => \N__36973\
        );

    \I__6171\ : InMux
    port map (
            O => \N__36980\,
            I => \N__36970\
        );

    \I__6170\ : InMux
    port map (
            O => \N__36977\,
            I => \N__36962\
        );

    \I__6169\ : InMux
    port map (
            O => \N__36976\,
            I => \N__36955\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__36973\,
            I => \N__36944\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__36970\,
            I => \N__36944\
        );

    \I__6166\ : InMux
    port map (
            O => \N__36969\,
            I => \N__36941\
        );

    \I__6165\ : InMux
    port map (
            O => \N__36968\,
            I => \N__36932\
        );

    \I__6164\ : InMux
    port map (
            O => \N__36967\,
            I => \N__36932\
        );

    \I__6163\ : InMux
    port map (
            O => \N__36966\,
            I => \N__36932\
        );

    \I__6162\ : InMux
    port map (
            O => \N__36965\,
            I => \N__36927\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__36962\,
            I => \N__36922\
        );

    \I__6160\ : InMux
    port map (
            O => \N__36961\,
            I => \N__36917\
        );

    \I__6159\ : InMux
    port map (
            O => \N__36960\,
            I => \N__36917\
        );

    \I__6158\ : InMux
    port map (
            O => \N__36959\,
            I => \N__36912\
        );

    \I__6157\ : InMux
    port map (
            O => \N__36958\,
            I => \N__36912\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__36955\,
            I => \N__36909\
        );

    \I__6155\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36905\
        );

    \I__6154\ : InMux
    port map (
            O => \N__36953\,
            I => \N__36902\
        );

    \I__6153\ : InMux
    port map (
            O => \N__36952\,
            I => \N__36897\
        );

    \I__6152\ : InMux
    port map (
            O => \N__36951\,
            I => \N__36897\
        );

    \I__6151\ : InMux
    port map (
            O => \N__36950\,
            I => \N__36894\
        );

    \I__6150\ : InMux
    port map (
            O => \N__36949\,
            I => \N__36891\
        );

    \I__6149\ : Span4Mux_h
    port map (
            O => \N__36944\,
            I => \N__36886\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__36941\,
            I => \N__36886\
        );

    \I__6147\ : InMux
    port map (
            O => \N__36940\,
            I => \N__36880\
        );

    \I__6146\ : InMux
    port map (
            O => \N__36939\,
            I => \N__36880\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__36932\,
            I => \N__36877\
        );

    \I__6144\ : InMux
    port map (
            O => \N__36931\,
            I => \N__36871\
        );

    \I__6143\ : InMux
    port map (
            O => \N__36930\,
            I => \N__36871\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__36927\,
            I => \N__36868\
        );

    \I__6141\ : CascadeMux
    port map (
            O => \N__36926\,
            I => \N__36865\
        );

    \I__6140\ : InMux
    port map (
            O => \N__36925\,
            I => \N__36861\
        );

    \I__6139\ : Span4Mux_v
    port map (
            O => \N__36922\,
            I => \N__36858\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__36917\,
            I => \N__36853\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__36912\,
            I => \N__36853\
        );

    \I__6136\ : Span4Mux_h
    port map (
            O => \N__36909\,
            I => \N__36850\
        );

    \I__6135\ : InMux
    port map (
            O => \N__36908\,
            I => \N__36847\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__36905\,
            I => \N__36844\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__36902\,
            I => \N__36839\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__36897\,
            I => \N__36839\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__36894\,
            I => \N__36834\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__36891\,
            I => \N__36834\
        );

    \I__6129\ : Span4Mux_v
    port map (
            O => \N__36886\,
            I => \N__36831\
        );

    \I__6128\ : InMux
    port map (
            O => \N__36885\,
            I => \N__36828\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__36880\,
            I => \N__36823\
        );

    \I__6126\ : Span4Mux_h
    port map (
            O => \N__36877\,
            I => \N__36823\
        );

    \I__6125\ : InMux
    port map (
            O => \N__36876\,
            I => \N__36820\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__36871\,
            I => \N__36815\
        );

    \I__6123\ : Span4Mux_v
    port map (
            O => \N__36868\,
            I => \N__36815\
        );

    \I__6122\ : InMux
    port map (
            O => \N__36865\,
            I => \N__36810\
        );

    \I__6121\ : InMux
    port map (
            O => \N__36864\,
            I => \N__36810\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__36861\,
            I => \N__36803\
        );

    \I__6119\ : Span4Mux_v
    port map (
            O => \N__36858\,
            I => \N__36803\
        );

    \I__6118\ : Span4Mux_v
    port map (
            O => \N__36853\,
            I => \N__36803\
        );

    \I__6117\ : Span4Mux_v
    port map (
            O => \N__36850\,
            I => \N__36800\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__36847\,
            I => \N__36789\
        );

    \I__6115\ : Span4Mux_v
    port map (
            O => \N__36844\,
            I => \N__36789\
        );

    \I__6114\ : Span4Mux_h
    port map (
            O => \N__36839\,
            I => \N__36789\
        );

    \I__6113\ : Span4Mux_h
    port map (
            O => \N__36834\,
            I => \N__36789\
        );

    \I__6112\ : Span4Mux_h
    port map (
            O => \N__36831\,
            I => \N__36789\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__36828\,
            I => \N__36778\
        );

    \I__6110\ : Span4Mux_v
    port map (
            O => \N__36823\,
            I => \N__36778\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__36820\,
            I => \N__36778\
        );

    \I__6108\ : Span4Mux_h
    port map (
            O => \N__36815\,
            I => \N__36778\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__36810\,
            I => \N__36778\
        );

    \I__6106\ : Odrv4
    port map (
            O => \N__36803\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__6105\ : Odrv4
    port map (
            O => \N__36800\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__6104\ : Odrv4
    port map (
            O => \N__36789\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__6103\ : Odrv4
    port map (
            O => \N__36778\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__6102\ : CascadeMux
    port map (
            O => \N__36769\,
            I => \c0.n21576_cascade_\
        );

    \I__6101\ : CascadeMux
    port map (
            O => \N__36766\,
            I => \N__36761\
        );

    \I__6100\ : InMux
    port map (
            O => \N__36765\,
            I => \N__36750\
        );

    \I__6099\ : InMux
    port map (
            O => \N__36764\,
            I => \N__36750\
        );

    \I__6098\ : InMux
    port map (
            O => \N__36761\,
            I => \N__36747\
        );

    \I__6097\ : CascadeMux
    port map (
            O => \N__36760\,
            I => \N__36743\
        );

    \I__6096\ : InMux
    port map (
            O => \N__36759\,
            I => \N__36740\
        );

    \I__6095\ : InMux
    port map (
            O => \N__36758\,
            I => \N__36737\
        );

    \I__6094\ : CascadeMux
    port map (
            O => \N__36757\,
            I => \N__36732\
        );

    \I__6093\ : InMux
    port map (
            O => \N__36756\,
            I => \N__36720\
        );

    \I__6092\ : InMux
    port map (
            O => \N__36755\,
            I => \N__36717\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__36750\,
            I => \N__36711\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__36747\,
            I => \N__36711\
        );

    \I__6089\ : InMux
    port map (
            O => \N__36746\,
            I => \N__36708\
        );

    \I__6088\ : InMux
    port map (
            O => \N__36743\,
            I => \N__36704\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__36740\,
            I => \N__36690\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__36737\,
            I => \N__36690\
        );

    \I__6085\ : InMux
    port map (
            O => \N__36736\,
            I => \N__36687\
        );

    \I__6084\ : InMux
    port map (
            O => \N__36735\,
            I => \N__36684\
        );

    \I__6083\ : InMux
    port map (
            O => \N__36732\,
            I => \N__36679\
        );

    \I__6082\ : InMux
    port map (
            O => \N__36731\,
            I => \N__36679\
        );

    \I__6081\ : InMux
    port map (
            O => \N__36730\,
            I => \N__36670\
        );

    \I__6080\ : InMux
    port map (
            O => \N__36729\,
            I => \N__36670\
        );

    \I__6079\ : InMux
    port map (
            O => \N__36728\,
            I => \N__36670\
        );

    \I__6078\ : InMux
    port map (
            O => \N__36727\,
            I => \N__36670\
        );

    \I__6077\ : InMux
    port map (
            O => \N__36726\,
            I => \N__36661\
        );

    \I__6076\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36661\
        );

    \I__6075\ : InMux
    port map (
            O => \N__36724\,
            I => \N__36661\
        );

    \I__6074\ : InMux
    port map (
            O => \N__36723\,
            I => \N__36661\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__36720\,
            I => \N__36656\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__36717\,
            I => \N__36656\
        );

    \I__6071\ : InMux
    port map (
            O => \N__36716\,
            I => \N__36653\
        );

    \I__6070\ : Span4Mux_h
    port map (
            O => \N__36711\,
            I => \N__36648\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__36708\,
            I => \N__36648\
        );

    \I__6068\ : InMux
    port map (
            O => \N__36707\,
            I => \N__36645\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__36704\,
            I => \N__36642\
        );

    \I__6066\ : InMux
    port map (
            O => \N__36703\,
            I => \N__36637\
        );

    \I__6065\ : InMux
    port map (
            O => \N__36702\,
            I => \N__36637\
        );

    \I__6064\ : InMux
    port map (
            O => \N__36701\,
            I => \N__36634\
        );

    \I__6063\ : InMux
    port map (
            O => \N__36700\,
            I => \N__36628\
        );

    \I__6062\ : InMux
    port map (
            O => \N__36699\,
            I => \N__36628\
        );

    \I__6061\ : InMux
    port map (
            O => \N__36698\,
            I => \N__36625\
        );

    \I__6060\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36618\
        );

    \I__6059\ : InMux
    port map (
            O => \N__36696\,
            I => \N__36613\
        );

    \I__6058\ : InMux
    port map (
            O => \N__36695\,
            I => \N__36613\
        );

    \I__6057\ : Span4Mux_v
    port map (
            O => \N__36690\,
            I => \N__36608\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__36687\,
            I => \N__36608\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__36684\,
            I => \N__36595\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__36679\,
            I => \N__36595\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__36670\,
            I => \N__36595\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__36661\,
            I => \N__36595\
        );

    \I__6051\ : Span4Mux_h
    port map (
            O => \N__36656\,
            I => \N__36595\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__36653\,
            I => \N__36595\
        );

    \I__6049\ : Span4Mux_h
    port map (
            O => \N__36648\,
            I => \N__36590\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__36645\,
            I => \N__36590\
        );

    \I__6047\ : Span4Mux_h
    port map (
            O => \N__36642\,
            I => \N__36585\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__36637\,
            I => \N__36580\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__36634\,
            I => \N__36580\
        );

    \I__6044\ : InMux
    port map (
            O => \N__36633\,
            I => \N__36577\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__36628\,
            I => \N__36574\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__36625\,
            I => \N__36571\
        );

    \I__6041\ : InMux
    port map (
            O => \N__36624\,
            I => \N__36564\
        );

    \I__6040\ : InMux
    port map (
            O => \N__36623\,
            I => \N__36564\
        );

    \I__6039\ : InMux
    port map (
            O => \N__36622\,
            I => \N__36564\
        );

    \I__6038\ : InMux
    port map (
            O => \N__36621\,
            I => \N__36561\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__36618\,
            I => \N__36552\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__36613\,
            I => \N__36552\
        );

    \I__6035\ : Span4Mux_v
    port map (
            O => \N__36608\,
            I => \N__36552\
        );

    \I__6034\ : Span4Mux_v
    port map (
            O => \N__36595\,
            I => \N__36552\
        );

    \I__6033\ : Span4Mux_v
    port map (
            O => \N__36590\,
            I => \N__36549\
        );

    \I__6032\ : InMux
    port map (
            O => \N__36589\,
            I => \N__36546\
        );

    \I__6031\ : InMux
    port map (
            O => \N__36588\,
            I => \N__36543\
        );

    \I__6030\ : Span4Mux_v
    port map (
            O => \N__36585\,
            I => \N__36538\
        );

    \I__6029\ : Span4Mux_h
    port map (
            O => \N__36580\,
            I => \N__36538\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__36577\,
            I => \N__36535\
        );

    \I__6027\ : Span4Mux_h
    port map (
            O => \N__36574\,
            I => \N__36526\
        );

    \I__6026\ : Span4Mux_v
    port map (
            O => \N__36571\,
            I => \N__36526\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__36564\,
            I => \N__36526\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__36561\,
            I => \N__36526\
        );

    \I__6023\ : Span4Mux_v
    port map (
            O => \N__36552\,
            I => \N__36521\
        );

    \I__6022\ : Span4Mux_h
    port map (
            O => \N__36549\,
            I => \N__36521\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__36546\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__36543\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6019\ : Odrv4
    port map (
            O => \N__36538\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6018\ : Odrv4
    port map (
            O => \N__36535\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6017\ : Odrv4
    port map (
            O => \N__36526\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6016\ : Odrv4
    port map (
            O => \N__36521\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6015\ : CascadeMux
    port map (
            O => \N__36508\,
            I => \c0.n21302_cascade_\
        );

    \I__6014\ : CascadeMux
    port map (
            O => \N__36505\,
            I => \c0.n21304_cascade_\
        );

    \I__6013\ : InMux
    port map (
            O => \N__36502\,
            I => \N__36499\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__36499\,
            I => \N__36496\
        );

    \I__6011\ : Span4Mux_h
    port map (
            O => \N__36496\,
            I => \N__36493\
        );

    \I__6010\ : Span4Mux_h
    port map (
            O => \N__36493\,
            I => \N__36490\
        );

    \I__6009\ : Odrv4
    port map (
            O => \N__36490\,
            I => \c0.n21572\
        );

    \I__6008\ : CascadeMux
    port map (
            O => \N__36487\,
            I => \N__36484\
        );

    \I__6007\ : InMux
    port map (
            O => \N__36484\,
            I => \N__36478\
        );

    \I__6006\ : InMux
    port map (
            O => \N__36483\,
            I => \N__36478\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__36478\,
            I => data_out_frame_5_4
        );

    \I__6004\ : InMux
    port map (
            O => \N__36475\,
            I => \N__36472\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__36472\,
            I => \N__36469\
        );

    \I__6002\ : Span4Mux_v
    port map (
            O => \N__36469\,
            I => \N__36466\
        );

    \I__6001\ : Span4Mux_h
    port map (
            O => \N__36466\,
            I => \N__36463\
        );

    \I__6000\ : Odrv4
    port map (
            O => \N__36463\,
            I => \c0.n21465\
        );

    \I__5999\ : InMux
    port map (
            O => \N__36460\,
            I => \N__36456\
        );

    \I__5998\ : InMux
    port map (
            O => \N__36459\,
            I => \N__36453\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__36456\,
            I => \c0.data_out_frame_5_0\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__36453\,
            I => \c0.data_out_frame_5_0\
        );

    \I__5995\ : InMux
    port map (
            O => \N__36448\,
            I => \N__36445\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__36445\,
            I => \N__36442\
        );

    \I__5993\ : Span4Mux_v
    port map (
            O => \N__36442\,
            I => \N__36438\
        );

    \I__5992\ : InMux
    port map (
            O => \N__36441\,
            I => \N__36435\
        );

    \I__5991\ : Odrv4
    port map (
            O => \N__36438\,
            I => control_mode_5
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__36435\,
            I => control_mode_5
        );

    \I__5989\ : InMux
    port map (
            O => \N__36430\,
            I => \N__36427\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__36427\,
            I => \N__36424\
        );

    \I__5987\ : Span4Mux_v
    port map (
            O => \N__36424\,
            I => \N__36421\
        );

    \I__5986\ : Odrv4
    port map (
            O => \N__36421\,
            I => \c0.n21638\
        );

    \I__5985\ : CascadeMux
    port map (
            O => \N__36418\,
            I => \N__36415\
        );

    \I__5984\ : InMux
    port map (
            O => \N__36415\,
            I => \N__36412\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__36412\,
            I => \N__36409\
        );

    \I__5982\ : Span4Mux_h
    port map (
            O => \N__36409\,
            I => \N__36406\
        );

    \I__5981\ : Odrv4
    port map (
            O => \N__36406\,
            I => \c0.n11_adj_3462\
        );

    \I__5980\ : InMux
    port map (
            O => \N__36403\,
            I => \N__36399\
        );

    \I__5979\ : InMux
    port map (
            O => \N__36402\,
            I => \N__36396\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__36399\,
            I => \N__36393\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__36396\,
            I => data_out_frame_5_2
        );

    \I__5976\ : Odrv12
    port map (
            O => \N__36393\,
            I => data_out_frame_5_2
        );

    \I__5975\ : InMux
    port map (
            O => \N__36388\,
            I => \N__36385\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__36385\,
            I => \N__36382\
        );

    \I__5973\ : Span4Mux_h
    port map (
            O => \N__36382\,
            I => \N__36379\
        );

    \I__5972\ : Odrv4
    port map (
            O => \N__36379\,
            I => \c0.rx.n9\
        );

    \I__5971\ : InMux
    port map (
            O => \N__36376\,
            I => \N__36373\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__36373\,
            I => \c0.n11_adj_3325\
        );

    \I__5969\ : InMux
    port map (
            O => \N__36370\,
            I => \N__36366\
        );

    \I__5968\ : CascadeMux
    port map (
            O => \N__36369\,
            I => \N__36363\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__36366\,
            I => \N__36360\
        );

    \I__5966\ : InMux
    port map (
            O => \N__36363\,
            I => \N__36357\
        );

    \I__5965\ : Span4Mux_v
    port map (
            O => \N__36360\,
            I => \N__36353\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__36357\,
            I => \N__36350\
        );

    \I__5963\ : InMux
    port map (
            O => \N__36356\,
            I => \N__36347\
        );

    \I__5962\ : Span4Mux_h
    port map (
            O => \N__36353\,
            I => \N__36344\
        );

    \I__5961\ : Span4Mux_h
    port map (
            O => \N__36350\,
            I => \N__36341\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__36347\,
            I => encoder1_position_8
        );

    \I__5959\ : Odrv4
    port map (
            O => \N__36344\,
            I => encoder1_position_8
        );

    \I__5958\ : Odrv4
    port map (
            O => \N__36341\,
            I => encoder1_position_8
        );

    \I__5957\ : CascadeMux
    port map (
            O => \N__36334\,
            I => \N__36331\
        );

    \I__5956\ : InMux
    port map (
            O => \N__36331\,
            I => \N__36325\
        );

    \I__5955\ : InMux
    port map (
            O => \N__36330\,
            I => \N__36325\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__36325\,
            I => data_out_frame_12_0
        );

    \I__5953\ : CascadeMux
    port map (
            O => \N__36322\,
            I => \N__36319\
        );

    \I__5952\ : InMux
    port map (
            O => \N__36319\,
            I => \N__36315\
        );

    \I__5951\ : InMux
    port map (
            O => \N__36318\,
            I => \N__36312\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__36315\,
            I => \N__36308\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__36312\,
            I => \N__36305\
        );

    \I__5948\ : InMux
    port map (
            O => \N__36311\,
            I => \N__36302\
        );

    \I__5947\ : Span4Mux_h
    port map (
            O => \N__36308\,
            I => \N__36299\
        );

    \I__5946\ : Odrv4
    port map (
            O => \N__36305\,
            I => encoder1_position_23
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__36302\,
            I => encoder1_position_23
        );

    \I__5944\ : Odrv4
    port map (
            O => \N__36299\,
            I => encoder1_position_23
        );

    \I__5943\ : CascadeMux
    port map (
            O => \N__36292\,
            I => \N__36288\
        );

    \I__5942\ : InMux
    port map (
            O => \N__36291\,
            I => \N__36285\
        );

    \I__5941\ : InMux
    port map (
            O => \N__36288\,
            I => \N__36282\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__36285\,
            I => data_out_frame_11_7
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__36282\,
            I => data_out_frame_11_7
        );

    \I__5938\ : InMux
    port map (
            O => \N__36277\,
            I => \N__36274\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__36274\,
            I => \N__36271\
        );

    \I__5936\ : Span4Mux_v
    port map (
            O => \N__36271\,
            I => \N__36268\
        );

    \I__5935\ : Span4Mux_h
    port map (
            O => \N__36268\,
            I => \N__36265\
        );

    \I__5934\ : Odrv4
    port map (
            O => \N__36265\,
            I => n2317
        );

    \I__5933\ : InMux
    port map (
            O => \N__36262\,
            I => \N__36251\
        );

    \I__5932\ : InMux
    port map (
            O => \N__36261\,
            I => \N__36240\
        );

    \I__5931\ : InMux
    port map (
            O => \N__36260\,
            I => \N__36240\
        );

    \I__5930\ : InMux
    port map (
            O => \N__36259\,
            I => \N__36231\
        );

    \I__5929\ : InMux
    port map (
            O => \N__36258\,
            I => \N__36231\
        );

    \I__5928\ : InMux
    port map (
            O => \N__36257\,
            I => \N__36231\
        );

    \I__5927\ : InMux
    port map (
            O => \N__36256\,
            I => \N__36231\
        );

    \I__5926\ : InMux
    port map (
            O => \N__36255\,
            I => \N__36218\
        );

    \I__5925\ : InMux
    port map (
            O => \N__36254\,
            I => \N__36215\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__36251\,
            I => \N__36212\
        );

    \I__5923\ : InMux
    port map (
            O => \N__36250\,
            I => \N__36207\
        );

    \I__5922\ : InMux
    port map (
            O => \N__36249\,
            I => \N__36207\
        );

    \I__5921\ : InMux
    port map (
            O => \N__36248\,
            I => \N__36204\
        );

    \I__5920\ : InMux
    port map (
            O => \N__36247\,
            I => \N__36201\
        );

    \I__5919\ : InMux
    port map (
            O => \N__36246\,
            I => \N__36196\
        );

    \I__5918\ : InMux
    port map (
            O => \N__36245\,
            I => \N__36196\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__36240\,
            I => \N__36191\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__36231\,
            I => \N__36191\
        );

    \I__5915\ : InMux
    port map (
            O => \N__36230\,
            I => \N__36184\
        );

    \I__5914\ : InMux
    port map (
            O => \N__36229\,
            I => \N__36184\
        );

    \I__5913\ : InMux
    port map (
            O => \N__36228\,
            I => \N__36184\
        );

    \I__5912\ : InMux
    port map (
            O => \N__36227\,
            I => \N__36181\
        );

    \I__5911\ : InMux
    port map (
            O => \N__36226\,
            I => \N__36169\
        );

    \I__5910\ : InMux
    port map (
            O => \N__36225\,
            I => \N__36169\
        );

    \I__5909\ : InMux
    port map (
            O => \N__36224\,
            I => \N__36166\
        );

    \I__5908\ : InMux
    port map (
            O => \N__36223\,
            I => \N__36159\
        );

    \I__5907\ : InMux
    port map (
            O => \N__36222\,
            I => \N__36159\
        );

    \I__5906\ : InMux
    port map (
            O => \N__36221\,
            I => \N__36159\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__36218\,
            I => \N__36150\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__36215\,
            I => \N__36150\
        );

    \I__5903\ : Span4Mux_v
    port map (
            O => \N__36212\,
            I => \N__36150\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__36207\,
            I => \N__36150\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__36204\,
            I => \N__36141\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__36201\,
            I => \N__36141\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__36196\,
            I => \N__36141\
        );

    \I__5898\ : Span4Mux_v
    port map (
            O => \N__36191\,
            I => \N__36141\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__36184\,
            I => \N__36138\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__36181\,
            I => \N__36135\
        );

    \I__5895\ : InMux
    port map (
            O => \N__36180\,
            I => \N__36120\
        );

    \I__5894\ : InMux
    port map (
            O => \N__36179\,
            I => \N__36120\
        );

    \I__5893\ : InMux
    port map (
            O => \N__36178\,
            I => \N__36120\
        );

    \I__5892\ : InMux
    port map (
            O => \N__36177\,
            I => \N__36120\
        );

    \I__5891\ : InMux
    port map (
            O => \N__36176\,
            I => \N__36120\
        );

    \I__5890\ : InMux
    port map (
            O => \N__36175\,
            I => \N__36120\
        );

    \I__5889\ : InMux
    port map (
            O => \N__36174\,
            I => \N__36120\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__36169\,
            I => \N__36117\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__36166\,
            I => \N__36112\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__36159\,
            I => \N__36112\
        );

    \I__5885\ : Span4Mux_v
    port map (
            O => \N__36150\,
            I => \N__36107\
        );

    \I__5884\ : Span4Mux_v
    port map (
            O => \N__36141\,
            I => \N__36107\
        );

    \I__5883\ : Span4Mux_h
    port map (
            O => \N__36138\,
            I => \N__36102\
        );

    \I__5882\ : Span4Mux_h
    port map (
            O => \N__36135\,
            I => \N__36102\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__36120\,
            I => \N__36095\
        );

    \I__5880\ : Span4Mux_h
    port map (
            O => \N__36117\,
            I => \N__36095\
        );

    \I__5879\ : Span4Mux_v
    port map (
            O => \N__36112\,
            I => \N__36095\
        );

    \I__5878\ : Sp12to4
    port map (
            O => \N__36107\,
            I => \N__36092\
        );

    \I__5877\ : Span4Mux_v
    port map (
            O => \N__36102\,
            I => \N__36089\
        );

    \I__5876\ : Odrv4
    port map (
            O => \N__36095\,
            I => count_enable_adj_3586
        );

    \I__5875\ : Odrv12
    port map (
            O => \N__36092\,
            I => count_enable_adj_3586
        );

    \I__5874\ : Odrv4
    port map (
            O => \N__36089\,
            I => count_enable_adj_3586
        );

    \I__5873\ : InMux
    port map (
            O => \N__36082\,
            I => \N__36079\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__36079\,
            I => \N__36075\
        );

    \I__5871\ : InMux
    port map (
            O => \N__36078\,
            I => \N__36071\
        );

    \I__5870\ : Span4Mux_h
    port map (
            O => \N__36075\,
            I => \N__36068\
        );

    \I__5869\ : InMux
    port map (
            O => \N__36074\,
            I => \N__36065\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__36071\,
            I => \N__36062\
        );

    \I__5867\ : Span4Mux_h
    port map (
            O => \N__36068\,
            I => \N__36059\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__36065\,
            I => \N__36054\
        );

    \I__5865\ : Span4Mux_v
    port map (
            O => \N__36062\,
            I => \N__36054\
        );

    \I__5864\ : Odrv4
    port map (
            O => \N__36059\,
            I => encoder1_position_28
        );

    \I__5863\ : Odrv4
    port map (
            O => \N__36054\,
            I => encoder1_position_28
        );

    \I__5862\ : InMux
    port map (
            O => \N__36049\,
            I => \N__36045\
        );

    \I__5861\ : InMux
    port map (
            O => \N__36048\,
            I => \N__36042\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__36045\,
            I => data_out_frame_5_6
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__36042\,
            I => data_out_frame_5_6
        );

    \I__5858\ : InMux
    port map (
            O => \N__36037\,
            I => \N__36034\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__36034\,
            I => \N__36030\
        );

    \I__5856\ : InMux
    port map (
            O => \N__36033\,
            I => \N__36027\
        );

    \I__5855\ : Span4Mux_h
    port map (
            O => \N__36030\,
            I => \N__36024\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__36027\,
            I => data_out_frame_29_3
        );

    \I__5853\ : Odrv4
    port map (
            O => \N__36024\,
            I => data_out_frame_29_3
        );

    \I__5852\ : InMux
    port map (
            O => \N__36019\,
            I => \N__36015\
        );

    \I__5851\ : InMux
    port map (
            O => \N__36018\,
            I => \N__36012\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__36015\,
            I => \c0.data_out_frame_28_3\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__36012\,
            I => \c0.data_out_frame_28_3\
        );

    \I__5848\ : CascadeMux
    port map (
            O => \N__36007\,
            I => \N__36004\
        );

    \I__5847\ : InMux
    port map (
            O => \N__36004\,
            I => \N__36001\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__36001\,
            I => \N__35996\
        );

    \I__5845\ : InMux
    port map (
            O => \N__36000\,
            I => \N__35993\
        );

    \I__5844\ : CascadeMux
    port map (
            O => \N__35999\,
            I => \N__35990\
        );

    \I__5843\ : Span4Mux_v
    port map (
            O => \N__35996\,
            I => \N__35985\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__35993\,
            I => \N__35985\
        );

    \I__5841\ : InMux
    port map (
            O => \N__35990\,
            I => \N__35982\
        );

    \I__5840\ : Span4Mux_v
    port map (
            O => \N__35985\,
            I => \N__35979\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__35982\,
            I => \N__35976\
        );

    \I__5838\ : Span4Mux_h
    port map (
            O => \N__35979\,
            I => \N__35973\
        );

    \I__5837\ : Span12Mux_h
    port map (
            O => \N__35976\,
            I => \N__35970\
        );

    \I__5836\ : Odrv4
    port map (
            O => \N__35973\,
            I => \c0.n9753\
        );

    \I__5835\ : Odrv12
    port map (
            O => \N__35970\,
            I => \c0.n9753\
        );

    \I__5834\ : CascadeMux
    port map (
            O => \N__35965\,
            I => \c0.n26_adj_3382_cascade_\
        );

    \I__5833\ : InMux
    port map (
            O => \N__35962\,
            I => \N__35959\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__35959\,
            I => \N__35956\
        );

    \I__5831\ : Odrv4
    port map (
            O => \N__35956\,
            I => \c0.n21314\
        );

    \I__5830\ : InMux
    port map (
            O => \N__35953\,
            I => \N__35950\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__35950\,
            I => \N__35947\
        );

    \I__5828\ : Span4Mux_v
    port map (
            O => \N__35947\,
            I => \N__35944\
        );

    \I__5827\ : Odrv4
    port map (
            O => \N__35944\,
            I => \c0.n21316\
        );

    \I__5826\ : InMux
    port map (
            O => \N__35941\,
            I => \N__35938\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__35938\,
            I => \N__35935\
        );

    \I__5824\ : Span12Mux_v
    port map (
            O => \N__35935\,
            I => \N__35932\
        );

    \I__5823\ : Odrv12
    port map (
            O => \N__35932\,
            I => \c0.n21562\
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__35929\,
            I => \c0.n21322_cascade_\
        );

    \I__5821\ : InMux
    port map (
            O => \N__35926\,
            I => \N__35923\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__35923\,
            I => \N__35920\
        );

    \I__5819\ : Span4Mux_v
    port map (
            O => \N__35920\,
            I => \N__35917\
        );

    \I__5818\ : Odrv4
    port map (
            O => \N__35917\,
            I => n10_adj_3594
        );

    \I__5817\ : InMux
    port map (
            O => \N__35914\,
            I => \N__35910\
        );

    \I__5816\ : InMux
    port map (
            O => \N__35913\,
            I => \N__35907\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__35910\,
            I => data_out_frame_7_2
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__35907\,
            I => data_out_frame_7_2
        );

    \I__5813\ : InMux
    port map (
            O => \N__35902\,
            I => \N__35899\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__35899\,
            I => \c0.n5_adj_3106\
        );

    \I__5811\ : InMux
    port map (
            O => \N__35896\,
            I => \N__35892\
        );

    \I__5810\ : CascadeMux
    port map (
            O => \N__35895\,
            I => \N__35888\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__35892\,
            I => \N__35885\
        );

    \I__5808\ : InMux
    port map (
            O => \N__35891\,
            I => \N__35882\
        );

    \I__5807\ : InMux
    port map (
            O => \N__35888\,
            I => \N__35879\
        );

    \I__5806\ : Odrv12
    port map (
            O => \N__35885\,
            I => encoder0_position_26
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__35882\,
            I => encoder0_position_26
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__35879\,
            I => encoder0_position_26
        );

    \I__5803\ : InMux
    port map (
            O => \N__35872\,
            I => \N__35868\
        );

    \I__5802\ : InMux
    port map (
            O => \N__35871\,
            I => \N__35865\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__35868\,
            I => data_out_frame_6_2
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__35865\,
            I => data_out_frame_6_2
        );

    \I__5799\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35854\
        );

    \I__5798\ : InMux
    port map (
            O => \N__35859\,
            I => \N__35854\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__35854\,
            I => \c0.data_out_frame_0_2\
        );

    \I__5796\ : CascadeMux
    port map (
            O => \N__35851\,
            I => \c0.n21473_cascade_\
        );

    \I__5795\ : InMux
    port map (
            O => \N__35848\,
            I => \N__35845\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__35845\,
            I => \N__35842\
        );

    \I__5793\ : Odrv4
    port map (
            O => \N__35842\,
            I => \c0.n6_adj_3105\
        );

    \I__5792\ : CascadeMux
    port map (
            O => \N__35839\,
            I => \N__35836\
        );

    \I__5791\ : InMux
    port map (
            O => \N__35836\,
            I => \N__35833\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__35833\,
            I => \N__35830\
        );

    \I__5789\ : Span4Mux_v
    port map (
            O => \N__35830\,
            I => \N__35826\
        );

    \I__5788\ : InMux
    port map (
            O => \N__35829\,
            I => \N__35823\
        );

    \I__5787\ : Span4Mux_h
    port map (
            O => \N__35826\,
            I => \N__35820\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__35823\,
            I => data_out_frame_28_6
        );

    \I__5785\ : Odrv4
    port map (
            O => \N__35820\,
            I => data_out_frame_28_6
        );

    \I__5784\ : InMux
    port map (
            O => \N__35815\,
            I => \N__35811\
        );

    \I__5783\ : InMux
    port map (
            O => \N__35814\,
            I => \N__35808\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__35811\,
            I => \c0.data_out_frame_0_3\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__35808\,
            I => \c0.data_out_frame_0_3\
        );

    \I__5780\ : SRMux
    port map (
            O => \N__35803\,
            I => \N__35800\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__35800\,
            I => \N__35797\
        );

    \I__5778\ : Span4Mux_h
    port map (
            O => \N__35797\,
            I => \N__35794\
        );

    \I__5777\ : Odrv4
    port map (
            O => \N__35794\,
            I => \c0.n6_adj_3150\
        );

    \I__5776\ : InMux
    port map (
            O => \N__35791\,
            I => \N__35788\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__35788\,
            I => \N__35785\
        );

    \I__5774\ : Span4Mux_h
    port map (
            O => \N__35785\,
            I => \N__35782\
        );

    \I__5773\ : Odrv4
    port map (
            O => \N__35782\,
            I => n2333
        );

    \I__5772\ : InMux
    port map (
            O => \N__35779\,
            I => \N__35776\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__35776\,
            I => \N__35773\
        );

    \I__5770\ : Span4Mux_h
    port map (
            O => \N__35773\,
            I => \N__35770\
        );

    \I__5769\ : Odrv4
    port map (
            O => \N__35770\,
            I => \c0.n21319\
        );

    \I__5768\ : InMux
    port map (
            O => \N__35767\,
            I => \N__35764\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__35764\,
            I => \N__35761\
        );

    \I__5766\ : Span4Mux_v
    port map (
            O => \N__35761\,
            I => \N__35757\
        );

    \I__5765\ : CascadeMux
    port map (
            O => \N__35760\,
            I => \N__35753\
        );

    \I__5764\ : Span4Mux_h
    port map (
            O => \N__35757\,
            I => \N__35750\
        );

    \I__5763\ : InMux
    port map (
            O => \N__35756\,
            I => \N__35747\
        );

    \I__5762\ : InMux
    port map (
            O => \N__35753\,
            I => \N__35744\
        );

    \I__5761\ : Odrv4
    port map (
            O => \N__35750\,
            I => encoder0_position_18
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__35747\,
            I => encoder0_position_18
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__35744\,
            I => encoder0_position_18
        );

    \I__5758\ : InMux
    port map (
            O => \N__35737\,
            I => \N__35734\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__35734\,
            I => \c0.n21317\
        );

    \I__5756\ : InMux
    port map (
            O => \N__35731\,
            I => \N__35725\
        );

    \I__5755\ : InMux
    port map (
            O => \N__35730\,
            I => \N__35706\
        );

    \I__5754\ : InMux
    port map (
            O => \N__35729\,
            I => \N__35701\
        );

    \I__5753\ : InMux
    port map (
            O => \N__35728\,
            I => \N__35701\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__35725\,
            I => \N__35698\
        );

    \I__5751\ : InMux
    port map (
            O => \N__35724\,
            I => \N__35695\
        );

    \I__5750\ : InMux
    port map (
            O => \N__35723\,
            I => \N__35692\
        );

    \I__5749\ : InMux
    port map (
            O => \N__35722\,
            I => \N__35689\
        );

    \I__5748\ : InMux
    port map (
            O => \N__35721\,
            I => \N__35684\
        );

    \I__5747\ : InMux
    port map (
            O => \N__35720\,
            I => \N__35681\
        );

    \I__5746\ : InMux
    port map (
            O => \N__35719\,
            I => \N__35678\
        );

    \I__5745\ : InMux
    port map (
            O => \N__35718\,
            I => \N__35663\
        );

    \I__5744\ : InMux
    port map (
            O => \N__35717\,
            I => \N__35663\
        );

    \I__5743\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35663\
        );

    \I__5742\ : InMux
    port map (
            O => \N__35715\,
            I => \N__35663\
        );

    \I__5741\ : InMux
    port map (
            O => \N__35714\,
            I => \N__35663\
        );

    \I__5740\ : InMux
    port map (
            O => \N__35713\,
            I => \N__35663\
        );

    \I__5739\ : InMux
    port map (
            O => \N__35712\,
            I => \N__35663\
        );

    \I__5738\ : InMux
    port map (
            O => \N__35711\,
            I => \N__35656\
        );

    \I__5737\ : InMux
    port map (
            O => \N__35710\,
            I => \N__35656\
        );

    \I__5736\ : InMux
    port map (
            O => \N__35709\,
            I => \N__35656\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__35706\,
            I => \N__35645\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__35701\,
            I => \N__35645\
        );

    \I__5733\ : Span4Mux_h
    port map (
            O => \N__35698\,
            I => \N__35645\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__35695\,
            I => \N__35645\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__35692\,
            I => \N__35645\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__35689\,
            I => \N__35642\
        );

    \I__5729\ : InMux
    port map (
            O => \N__35688\,
            I => \N__35629\
        );

    \I__5728\ : InMux
    port map (
            O => \N__35687\,
            I => \N__35626\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__35684\,
            I => \N__35621\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__35681\,
            I => \N__35621\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__35678\,
            I => \N__35614\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__35663\,
            I => \N__35614\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__35656\,
            I => \N__35614\
        );

    \I__5722\ : Span4Mux_v
    port map (
            O => \N__35645\,
            I => \N__35609\
        );

    \I__5721\ : Span4Mux_h
    port map (
            O => \N__35642\,
            I => \N__35609\
        );

    \I__5720\ : InMux
    port map (
            O => \N__35641\,
            I => \N__35604\
        );

    \I__5719\ : InMux
    port map (
            O => \N__35640\,
            I => \N__35604\
        );

    \I__5718\ : InMux
    port map (
            O => \N__35639\,
            I => \N__35587\
        );

    \I__5717\ : InMux
    port map (
            O => \N__35638\,
            I => \N__35587\
        );

    \I__5716\ : InMux
    port map (
            O => \N__35637\,
            I => \N__35587\
        );

    \I__5715\ : InMux
    port map (
            O => \N__35636\,
            I => \N__35587\
        );

    \I__5714\ : InMux
    port map (
            O => \N__35635\,
            I => \N__35587\
        );

    \I__5713\ : InMux
    port map (
            O => \N__35634\,
            I => \N__35587\
        );

    \I__5712\ : InMux
    port map (
            O => \N__35633\,
            I => \N__35587\
        );

    \I__5711\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35587\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__35629\,
            I => \N__35582\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__35626\,
            I => \N__35582\
        );

    \I__5708\ : Span4Mux_h
    port map (
            O => \N__35621\,
            I => \N__35577\
        );

    \I__5707\ : Span4Mux_v
    port map (
            O => \N__35614\,
            I => \N__35577\
        );

    \I__5706\ : Span4Mux_h
    port map (
            O => \N__35609\,
            I => \N__35574\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__35604\,
            I => count_enable
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__35587\,
            I => count_enable
        );

    \I__5703\ : Odrv12
    port map (
            O => \N__35582\,
            I => count_enable
        );

    \I__5702\ : Odrv4
    port map (
            O => \N__35577\,
            I => count_enable
        );

    \I__5701\ : Odrv4
    port map (
            O => \N__35574\,
            I => count_enable
        );

    \I__5700\ : InMux
    port map (
            O => \N__35563\,
            I => \N__35560\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__35560\,
            I => \N__35557\
        );

    \I__5698\ : Span4Mux_h
    port map (
            O => \N__35557\,
            I => \N__35554\
        );

    \I__5697\ : Span4Mux_h
    port map (
            O => \N__35554\,
            I => \N__35551\
        );

    \I__5696\ : Odrv4
    port map (
            O => \N__35551\,
            I => n2252
        );

    \I__5695\ : InMux
    port map (
            O => \N__35548\,
            I => \N__35544\
        );

    \I__5694\ : CascadeMux
    port map (
            O => \N__35547\,
            I => \N__35541\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__35544\,
            I => \N__35538\
        );

    \I__5692\ : InMux
    port map (
            O => \N__35541\,
            I => \N__35535\
        );

    \I__5691\ : Span4Mux_v
    port map (
            O => \N__35538\,
            I => \N__35530\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__35535\,
            I => \N__35530\
        );

    \I__5689\ : Span4Mux_h
    port map (
            O => \N__35530\,
            I => \N__35526\
        );

    \I__5688\ : InMux
    port map (
            O => \N__35529\,
            I => \N__35523\
        );

    \I__5687\ : Span4Mux_h
    port map (
            O => \N__35526\,
            I => \N__35520\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__35523\,
            I => encoder0_position_27
        );

    \I__5685\ : Odrv4
    port map (
            O => \N__35520\,
            I => encoder0_position_27
        );

    \I__5684\ : InMux
    port map (
            O => \N__35515\,
            I => \N__35511\
        );

    \I__5683\ : InMux
    port map (
            O => \N__35514\,
            I => \N__35508\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__35511\,
            I => data_out_frame_7_3
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__35508\,
            I => data_out_frame_7_3
        );

    \I__5680\ : InMux
    port map (
            O => \N__35503\,
            I => \N__35500\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__35500\,
            I => \N__35496\
        );

    \I__5678\ : InMux
    port map (
            O => \N__35499\,
            I => \N__35493\
        );

    \I__5677\ : Span4Mux_h
    port map (
            O => \N__35496\,
            I => \N__35490\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__35493\,
            I => data_out_frame_6_3
        );

    \I__5675\ : Odrv4
    port map (
            O => \N__35490\,
            I => data_out_frame_6_3
        );

    \I__5674\ : InMux
    port map (
            O => \N__35485\,
            I => \N__35482\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__35482\,
            I => \c0.n5_adj_3380\
        );

    \I__5672\ : InMux
    port map (
            O => \N__35479\,
            I => \N__35476\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__35476\,
            I => \c0.n21320\
        );

    \I__5670\ : InMux
    port map (
            O => \N__35473\,
            I => \N__35468\
        );

    \I__5669\ : InMux
    port map (
            O => \N__35472\,
            I => \N__35465\
        );

    \I__5668\ : InMux
    port map (
            O => \N__35471\,
            I => \N__35462\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__35468\,
            I => \N__35459\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__35465\,
            I => \N__35456\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__35462\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__5664\ : Odrv4
    port map (
            O => \N__35459\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__5663\ : Odrv4
    port map (
            O => \N__35456\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__5662\ : SRMux
    port map (
            O => \N__35449\,
            I => \N__35446\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__35446\,
            I => \N__35443\
        );

    \I__5660\ : Span4Mux_h
    port map (
            O => \N__35443\,
            I => \N__35440\
        );

    \I__5659\ : Odrv4
    port map (
            O => \N__35440\,
            I => \c0.n18675\
        );

    \I__5658\ : InMux
    port map (
            O => \N__35437\,
            I => \N__35433\
        );

    \I__5657\ : InMux
    port map (
            O => \N__35436\,
            I => \N__35430\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__35433\,
            I => \N__35427\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__35430\,
            I => \N__35424\
        );

    \I__5654\ : Span4Mux_h
    port map (
            O => \N__35427\,
            I => \N__35420\
        );

    \I__5653\ : Span4Mux_h
    port map (
            O => \N__35424\,
            I => \N__35415\
        );

    \I__5652\ : InMux
    port map (
            O => \N__35423\,
            I => \N__35412\
        );

    \I__5651\ : Sp12to4
    port map (
            O => \N__35420\,
            I => \N__35409\
        );

    \I__5650\ : InMux
    port map (
            O => \N__35419\,
            I => \N__35406\
        );

    \I__5649\ : InMux
    port map (
            O => \N__35418\,
            I => \N__35403\
        );

    \I__5648\ : Span4Mux_v
    port map (
            O => \N__35415\,
            I => \N__35398\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__35412\,
            I => \N__35398\
        );

    \I__5646\ : Span12Mux_v
    port map (
            O => \N__35409\,
            I => \N__35395\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__35406\,
            I => \N__35392\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__35403\,
            I => \N__35387\
        );

    \I__5643\ : Span4Mux_h
    port map (
            O => \N__35398\,
            I => \N__35387\
        );

    \I__5642\ : Odrv12
    port map (
            O => \N__35395\,
            I => n11289
        );

    \I__5641\ : Odrv4
    port map (
            O => \N__35392\,
            I => n11289
        );

    \I__5640\ : Odrv4
    port map (
            O => \N__35387\,
            I => n11289
        );

    \I__5639\ : InMux
    port map (
            O => \N__35380\,
            I => \N__35377\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__35377\,
            I => \N__35372\
        );

    \I__5637\ : InMux
    port map (
            O => \N__35376\,
            I => \N__35369\
        );

    \I__5636\ : InMux
    port map (
            O => \N__35375\,
            I => \N__35366\
        );

    \I__5635\ : Span4Mux_v
    port map (
            O => \N__35372\,
            I => \N__35363\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__35369\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__35366\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__5632\ : Odrv4
    port map (
            O => \N__35363\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__5631\ : CascadeMux
    port map (
            O => \N__35356\,
            I => \n2108_cascade_\
        );

    \I__5630\ : SRMux
    port map (
            O => \N__35353\,
            I => \N__35350\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__35350\,
            I => \N__35347\
        );

    \I__5628\ : Odrv12
    port map (
            O => \N__35347\,
            I => \c0.n6_adj_3170\
        );

    \I__5627\ : SRMux
    port map (
            O => \N__35344\,
            I => \N__35341\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__35341\,
            I => \N__35338\
        );

    \I__5625\ : Span4Mux_h
    port map (
            O => \N__35338\,
            I => \N__35335\
        );

    \I__5624\ : Odrv4
    port map (
            O => \N__35335\,
            I => \c0.n6_adj_3165\
        );

    \I__5623\ : InMux
    port map (
            O => \N__35332\,
            I => \N__35329\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__35329\,
            I => \N__35324\
        );

    \I__5621\ : InMux
    port map (
            O => \N__35328\,
            I => \N__35321\
        );

    \I__5620\ : InMux
    port map (
            O => \N__35327\,
            I => \N__35318\
        );

    \I__5619\ : Span4Mux_v
    port map (
            O => \N__35324\,
            I => \N__35315\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__35321\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__35318\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__5616\ : Odrv4
    port map (
            O => \N__35315\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__5615\ : SRMux
    port map (
            O => \N__35308\,
            I => \N__35305\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__35305\,
            I => \c0.n6_adj_3168\
        );

    \I__5613\ : CascadeMux
    port map (
            O => \N__35302\,
            I => \N__35299\
        );

    \I__5612\ : InMux
    port map (
            O => \N__35299\,
            I => \N__35296\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__35296\,
            I => \N__35293\
        );

    \I__5610\ : Span4Mux_h
    port map (
            O => \N__35293\,
            I => \N__35288\
        );

    \I__5609\ : InMux
    port map (
            O => \N__35292\,
            I => \N__35285\
        );

    \I__5608\ : InMux
    port map (
            O => \N__35291\,
            I => \N__35282\
        );

    \I__5607\ : Span4Mux_v
    port map (
            O => \N__35288\,
            I => \N__35279\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__35285\,
            I => \c0.FRAME_MATCHER_i_28\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__35282\,
            I => \c0.FRAME_MATCHER_i_28\
        );

    \I__5604\ : Odrv4
    port map (
            O => \N__35279\,
            I => \c0.FRAME_MATCHER_i_28\
        );

    \I__5603\ : SRMux
    port map (
            O => \N__35272\,
            I => \N__35269\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__35269\,
            I => \N__35266\
        );

    \I__5601\ : Odrv12
    port map (
            O => \N__35266\,
            I => \c0.n6_adj_3166\
        );

    \I__5600\ : SRMux
    port map (
            O => \N__35263\,
            I => \N__35260\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__35260\,
            I => \N__35257\
        );

    \I__5598\ : Span4Mux_s1_v
    port map (
            O => \N__35257\,
            I => \N__35254\
        );

    \I__5597\ : Odrv4
    port map (
            O => \N__35254\,
            I => \c0.n6_adj_3159\
        );

    \I__5596\ : InMux
    port map (
            O => \N__35251\,
            I => \N__35248\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__35248\,
            I => \N__35243\
        );

    \I__5594\ : InMux
    port map (
            O => \N__35247\,
            I => \N__35240\
        );

    \I__5593\ : InMux
    port map (
            O => \N__35246\,
            I => \N__35237\
        );

    \I__5592\ : Span4Mux_v
    port map (
            O => \N__35243\,
            I => \N__35234\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__35240\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__35237\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__5589\ : Odrv4
    port map (
            O => \N__35234\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__5588\ : SRMux
    port map (
            O => \N__35227\,
            I => \N__35224\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__35224\,
            I => \N__35221\
        );

    \I__5586\ : Odrv12
    port map (
            O => \N__35221\,
            I => \c0.n6_adj_3164\
        );

    \I__5585\ : SRMux
    port map (
            O => \N__35218\,
            I => \N__35215\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__35215\,
            I => \N__35212\
        );

    \I__5583\ : Odrv12
    port map (
            O => \N__35212\,
            I => \c0.n18653\
        );

    \I__5582\ : InMux
    port map (
            O => \N__35209\,
            I => \N__35204\
        );

    \I__5581\ : InMux
    port map (
            O => \N__35208\,
            I => \N__35201\
        );

    \I__5580\ : InMux
    port map (
            O => \N__35207\,
            I => \N__35198\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__35204\,
            I => \N__35195\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__35201\,
            I => \N__35192\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__35198\,
            I => \N__35189\
        );

    \I__5576\ : Span4Mux_v
    port map (
            O => \N__35195\,
            I => \N__35186\
        );

    \I__5575\ : Span4Mux_h
    port map (
            O => \N__35192\,
            I => \N__35183\
        );

    \I__5574\ : Span4Mux_h
    port map (
            O => \N__35189\,
            I => \N__35180\
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__35186\,
            I => \c0.FRAME_MATCHER_state_31_N_1736_2\
        );

    \I__5572\ : Odrv4
    port map (
            O => \N__35183\,
            I => \c0.FRAME_MATCHER_state_31_N_1736_2\
        );

    \I__5571\ : Odrv4
    port map (
            O => \N__35180\,
            I => \c0.FRAME_MATCHER_state_31_N_1736_2\
        );

    \I__5570\ : InMux
    port map (
            O => \N__35173\,
            I => \N__35170\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__35170\,
            I => \N__35167\
        );

    \I__5568\ : Odrv4
    port map (
            O => \N__35167\,
            I => \c0.FRAME_MATCHER_state_31_N_1736_1\
        );

    \I__5567\ : SRMux
    port map (
            O => \N__35164\,
            I => \N__35161\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__35161\,
            I => \N__35158\
        );

    \I__5565\ : Odrv4
    port map (
            O => \N__35158\,
            I => \c0.n6_adj_3176\
        );

    \I__5564\ : InMux
    port map (
            O => \N__35155\,
            I => \N__35151\
        );

    \I__5563\ : InMux
    port map (
            O => \N__35154\,
            I => \N__35147\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__35151\,
            I => \N__35144\
        );

    \I__5561\ : InMux
    port map (
            O => \N__35150\,
            I => \N__35141\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__35147\,
            I => \c0.n11433\
        );

    \I__5559\ : Odrv4
    port map (
            O => \N__35144\,
            I => \c0.n11433\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__35141\,
            I => \c0.n11433\
        );

    \I__5557\ : CascadeMux
    port map (
            O => \N__35134\,
            I => \N__35130\
        );

    \I__5556\ : CascadeMux
    port map (
            O => \N__35133\,
            I => \N__35127\
        );

    \I__5555\ : InMux
    port map (
            O => \N__35130\,
            I => \N__35124\
        );

    \I__5554\ : InMux
    port map (
            O => \N__35127\,
            I => \N__35120\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__35124\,
            I => \N__35117\
        );

    \I__5552\ : InMux
    port map (
            O => \N__35123\,
            I => \N__35114\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__35120\,
            I => \N__35111\
        );

    \I__5550\ : Span4Mux_h
    port map (
            O => \N__35117\,
            I => \N__35104\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__35114\,
            I => \N__35104\
        );

    \I__5548\ : Span4Mux_v
    port map (
            O => \N__35111\,
            I => \N__35104\
        );

    \I__5547\ : Span4Mux_v
    port map (
            O => \N__35104\,
            I => \N__35101\
        );

    \I__5546\ : Span4Mux_v
    port map (
            O => \N__35101\,
            I => \N__35098\
        );

    \I__5545\ : Odrv4
    port map (
            O => \N__35098\,
            I => \c0.n700\
        );

    \I__5544\ : InMux
    port map (
            O => \N__35095\,
            I => \N__35092\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__35092\,
            I => \N__35089\
        );

    \I__5542\ : Span4Mux_h
    port map (
            O => \N__35089\,
            I => \N__35086\
        );

    \I__5541\ : Odrv4
    port map (
            O => \N__35086\,
            I => \c0.n1\
        );

    \I__5540\ : InMux
    port map (
            O => \N__35083\,
            I => \N__35080\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__35080\,
            I => \N__35075\
        );

    \I__5538\ : InMux
    port map (
            O => \N__35079\,
            I => \N__35072\
        );

    \I__5537\ : InMux
    port map (
            O => \N__35078\,
            I => \N__35069\
        );

    \I__5536\ : Span4Mux_v
    port map (
            O => \N__35075\,
            I => \N__35066\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__35072\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__35069\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__5533\ : Odrv4
    port map (
            O => \N__35066\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__5532\ : CascadeMux
    port map (
            O => \N__35059\,
            I => \N__35056\
        );

    \I__5531\ : InMux
    port map (
            O => \N__35056\,
            I => \N__35052\
        );

    \I__5530\ : InMux
    port map (
            O => \N__35055\,
            I => \N__35049\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__35052\,
            I => \N__35046\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__35049\,
            I => \N__35043\
        );

    \I__5527\ : Span4Mux_v
    port map (
            O => \N__35046\,
            I => \N__35039\
        );

    \I__5526\ : Span4Mux_v
    port map (
            O => \N__35043\,
            I => \N__35036\
        );

    \I__5525\ : InMux
    port map (
            O => \N__35042\,
            I => \N__35033\
        );

    \I__5524\ : Span4Mux_v
    port map (
            O => \N__35039\,
            I => \N__35030\
        );

    \I__5523\ : Odrv4
    port map (
            O => \N__35036\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__35033\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__5521\ : Odrv4
    port map (
            O => \N__35030\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__5520\ : InMux
    port map (
            O => \N__35023\,
            I => \N__35020\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__35020\,
            I => \N__35017\
        );

    \I__5518\ : Odrv12
    port map (
            O => \N__35017\,
            I => \c0.n44_adj_3255\
        );

    \I__5517\ : InMux
    port map (
            O => \N__35014\,
            I => \N__35009\
        );

    \I__5516\ : InMux
    port map (
            O => \N__35013\,
            I => \N__35006\
        );

    \I__5515\ : InMux
    port map (
            O => \N__35012\,
            I => \N__35003\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__35009\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__35006\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__35003\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__5511\ : SRMux
    port map (
            O => \N__34996\,
            I => \N__34993\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__34993\,
            I => \N__34990\
        );

    \I__5509\ : Span4Mux_v
    port map (
            O => \N__34990\,
            I => \N__34987\
        );

    \I__5508\ : Span4Mux_h
    port map (
            O => \N__34987\,
            I => \N__34984\
        );

    \I__5507\ : Odrv4
    port map (
            O => \N__34984\,
            I => \c0.n6_adj_3174\
        );

    \I__5506\ : InMux
    port map (
            O => \N__34981\,
            I => \N__34978\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__34978\,
            I => \N__34975\
        );

    \I__5504\ : Odrv12
    port map (
            O => \N__34975\,
            I => \c0.n21273\
        );

    \I__5503\ : CascadeMux
    port map (
            O => \N__34972\,
            I => \c0.n5_adj_3306_cascade_\
        );

    \I__5502\ : CascadeMux
    port map (
            O => \N__34969\,
            I => \N__34966\
        );

    \I__5501\ : InMux
    port map (
            O => \N__34966\,
            I => \N__34960\
        );

    \I__5500\ : InMux
    port map (
            O => \N__34965\,
            I => \N__34960\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__34960\,
            I => \c0.n2_adj_3302\
        );

    \I__5498\ : CascadeMux
    port map (
            O => \N__34957\,
            I => \c0.n11433_cascade_\
        );

    \I__5497\ : CascadeMux
    port map (
            O => \N__34954\,
            I => \c0.n8_adj_3228_cascade_\
        );

    \I__5496\ : InMux
    port map (
            O => \N__34951\,
            I => \N__34947\
        );

    \I__5495\ : InMux
    port map (
            O => \N__34950\,
            I => \N__34944\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__34947\,
            I => \N__34941\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__34944\,
            I => \c0.n2103\
        );

    \I__5492\ : Odrv4
    port map (
            O => \N__34941\,
            I => \c0.n2103\
        );

    \I__5491\ : CascadeMux
    port map (
            O => \N__34936\,
            I => \c0.n2103_cascade_\
        );

    \I__5490\ : InMux
    port map (
            O => \N__34933\,
            I => \N__34928\
        );

    \I__5489\ : InMux
    port map (
            O => \N__34932\,
            I => \N__34925\
        );

    \I__5488\ : InMux
    port map (
            O => \N__34931\,
            I => \N__34922\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__34928\,
            I => \N__34919\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__34925\,
            I => \N__34916\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__34922\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__5484\ : Odrv12
    port map (
            O => \N__34919\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__5483\ : Odrv4
    port map (
            O => \N__34916\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__5482\ : CascadeMux
    port map (
            O => \N__34909\,
            I => \c0.n41_adj_3258_cascade_\
        );

    \I__5481\ : InMux
    port map (
            O => \N__34906\,
            I => \N__34903\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__34903\,
            I => \c0.n43_adj_3257\
        );

    \I__5479\ : InMux
    port map (
            O => \N__34900\,
            I => \N__34897\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__34897\,
            I => \N__34893\
        );

    \I__5477\ : InMux
    port map (
            O => \N__34896\,
            I => \N__34889\
        );

    \I__5476\ : Span4Mux_v
    port map (
            O => \N__34893\,
            I => \N__34886\
        );

    \I__5475\ : InMux
    port map (
            O => \N__34892\,
            I => \N__34883\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__34889\,
            I => \N__34878\
        );

    \I__5473\ : Span4Mux_v
    port map (
            O => \N__34886\,
            I => \N__34878\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__34883\,
            I => \c0.FRAME_MATCHER_i_10\
        );

    \I__5471\ : Odrv4
    port map (
            O => \N__34878\,
            I => \c0.FRAME_MATCHER_i_10\
        );

    \I__5470\ : InMux
    port map (
            O => \N__34873\,
            I => \N__34870\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__34870\,
            I => \N__34865\
        );

    \I__5468\ : InMux
    port map (
            O => \N__34869\,
            I => \N__34862\
        );

    \I__5467\ : InMux
    port map (
            O => \N__34868\,
            I => \N__34859\
        );

    \I__5466\ : Span4Mux_v
    port map (
            O => \N__34865\,
            I => \N__34856\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__34862\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__34859\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__5463\ : Odrv4
    port map (
            O => \N__34856\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__5462\ : InMux
    port map (
            O => \N__34849\,
            I => \N__34845\
        );

    \I__5461\ : InMux
    port map (
            O => \N__34848\,
            I => \N__34842\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__34845\,
            I => \N__34839\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__34842\,
            I => \N__34836\
        );

    \I__5458\ : Span4Mux_v
    port map (
            O => \N__34839\,
            I => \N__34832\
        );

    \I__5457\ : Span4Mux_v
    port map (
            O => \N__34836\,
            I => \N__34829\
        );

    \I__5456\ : InMux
    port map (
            O => \N__34835\,
            I => \N__34826\
        );

    \I__5455\ : Span4Mux_v
    port map (
            O => \N__34832\,
            I => \N__34823\
        );

    \I__5454\ : Odrv4
    port map (
            O => \N__34829\,
            I => \c0.FRAME_MATCHER_i_13\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__34826\,
            I => \c0.FRAME_MATCHER_i_13\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__34823\,
            I => \c0.FRAME_MATCHER_i_13\
        );

    \I__5451\ : InMux
    port map (
            O => \N__34816\,
            I => \N__34813\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__34813\,
            I => \N__34810\
        );

    \I__5449\ : Span4Mux_v
    port map (
            O => \N__34810\,
            I => \N__34806\
        );

    \I__5448\ : InMux
    port map (
            O => \N__34809\,
            I => \N__34803\
        );

    \I__5447\ : Span4Mux_v
    port map (
            O => \N__34806\,
            I => \N__34799\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__34803\,
            I => \N__34796\
        );

    \I__5445\ : InMux
    port map (
            O => \N__34802\,
            I => \N__34793\
        );

    \I__5444\ : Span4Mux_v
    port map (
            O => \N__34799\,
            I => \N__34790\
        );

    \I__5443\ : Odrv4
    port map (
            O => \N__34796\,
            I => \c0.FRAME_MATCHER_i_9\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__34793\,
            I => \c0.FRAME_MATCHER_i_9\
        );

    \I__5441\ : Odrv4
    port map (
            O => \N__34790\,
            I => \c0.FRAME_MATCHER_i_9\
        );

    \I__5440\ : InMux
    port map (
            O => \N__34783\,
            I => \N__34780\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__34780\,
            I => \c0.n40_adj_3259\
        );

    \I__5438\ : InMux
    port map (
            O => \N__34777\,
            I => \N__34774\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__34774\,
            I => \c0.n45_adj_3262\
        );

    \I__5436\ : CascadeMux
    port map (
            O => \N__34771\,
            I => \c0.n39_adj_3260_cascade_\
        );

    \I__5435\ : InMux
    port map (
            O => \N__34768\,
            I => \N__34765\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__34765\,
            I => \c0.n50_adj_3261\
        );

    \I__5433\ : InMux
    port map (
            O => \N__34762\,
            I => \N__34759\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__34759\,
            I => \N__34754\
        );

    \I__5431\ : InMux
    port map (
            O => \N__34758\,
            I => \N__34749\
        );

    \I__5430\ : InMux
    port map (
            O => \N__34757\,
            I => \N__34749\
        );

    \I__5429\ : Odrv4
    port map (
            O => \N__34754\,
            I => \c0.n11432\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__34749\,
            I => \c0.n11432\
        );

    \I__5427\ : CascadeMux
    port map (
            O => \N__34744\,
            I => \c0.n14_adj_3080_cascade_\
        );

    \I__5426\ : InMux
    port map (
            O => \N__34741\,
            I => \N__34738\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__34738\,
            I => \N__34735\
        );

    \I__5424\ : Span4Mux_h
    port map (
            O => \N__34735\,
            I => \N__34732\
        );

    \I__5423\ : Odrv4
    port map (
            O => \N__34732\,
            I => \c0.n10_adj_3081\
        );

    \I__5422\ : CascadeMux
    port map (
            O => \N__34729\,
            I => \N__34724\
        );

    \I__5421\ : InMux
    port map (
            O => \N__34728\,
            I => \N__34721\
        );

    \I__5420\ : InMux
    port map (
            O => \N__34727\,
            I => \N__34718\
        );

    \I__5419\ : InMux
    port map (
            O => \N__34724\,
            I => \N__34715\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__34721\,
            I => \N__34712\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__34718\,
            I => \N__34707\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__34715\,
            I => \N__34707\
        );

    \I__5415\ : Span4Mux_h
    port map (
            O => \N__34712\,
            I => \N__34704\
        );

    \I__5414\ : Odrv4
    port map (
            O => \N__34707\,
            I => \c0.n4812\
        );

    \I__5413\ : Odrv4
    port map (
            O => \N__34704\,
            I => \c0.n4812\
        );

    \I__5412\ : InMux
    port map (
            O => \N__34699\,
            I => \N__34696\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__34696\,
            I => \c0.n19119\
        );

    \I__5410\ : CascadeMux
    port map (
            O => \N__34693\,
            I => \c0.n19119_cascade_\
        );

    \I__5409\ : CascadeMux
    port map (
            O => \N__34690\,
            I => \N__34680\
        );

    \I__5408\ : CascadeMux
    port map (
            O => \N__34689\,
            I => \N__34677\
        );

    \I__5407\ : CascadeMux
    port map (
            O => \N__34688\,
            I => \N__34674\
        );

    \I__5406\ : CascadeMux
    port map (
            O => \N__34687\,
            I => \N__34671\
        );

    \I__5405\ : CascadeMux
    port map (
            O => \N__34686\,
            I => \N__34668\
        );

    \I__5404\ : CascadeMux
    port map (
            O => \N__34685\,
            I => \N__34665\
        );

    \I__5403\ : CascadeMux
    port map (
            O => \N__34684\,
            I => \N__34662\
        );

    \I__5402\ : CascadeMux
    port map (
            O => \N__34683\,
            I => \N__34659\
        );

    \I__5401\ : InMux
    port map (
            O => \N__34680\,
            I => \N__34650\
        );

    \I__5400\ : InMux
    port map (
            O => \N__34677\,
            I => \N__34650\
        );

    \I__5399\ : InMux
    port map (
            O => \N__34674\,
            I => \N__34650\
        );

    \I__5398\ : InMux
    port map (
            O => \N__34671\,
            I => \N__34650\
        );

    \I__5397\ : InMux
    port map (
            O => \N__34668\,
            I => \N__34641\
        );

    \I__5396\ : InMux
    port map (
            O => \N__34665\,
            I => \N__34641\
        );

    \I__5395\ : InMux
    port map (
            O => \N__34662\,
            I => \N__34641\
        );

    \I__5394\ : InMux
    port map (
            O => \N__34659\,
            I => \N__34641\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__34650\,
            I => \c0.rx.n3\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__34641\,
            I => \c0.rx.n3\
        );

    \I__5391\ : InMux
    port map (
            O => \N__34636\,
            I => \c0.rx.n17273\
        );

    \I__5390\ : InMux
    port map (
            O => \N__34633\,
            I => \N__34630\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__34630\,
            I => \c0.rx.n7\
        );

    \I__5388\ : CascadeMux
    port map (
            O => \N__34627\,
            I => \N__34624\
        );

    \I__5387\ : InMux
    port map (
            O => \N__34624\,
            I => \N__34621\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__34621\,
            I => \N__34618\
        );

    \I__5385\ : Span4Mux_v
    port map (
            O => \N__34618\,
            I => \N__34615\
        );

    \I__5384\ : Span4Mux_v
    port map (
            O => \N__34615\,
            I => \N__34611\
        );

    \I__5383\ : InMux
    port map (
            O => \N__34614\,
            I => \N__34607\
        );

    \I__5382\ : Span4Mux_v
    port map (
            O => \N__34611\,
            I => \N__34604\
        );

    \I__5381\ : InMux
    port map (
            O => \N__34610\,
            I => \N__34601\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__34607\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__5379\ : Odrv4
    port map (
            O => \N__34604\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__34601\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__5377\ : InMux
    port map (
            O => \N__34594\,
            I => \N__34591\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__34591\,
            I => \N__34586\
        );

    \I__5375\ : InMux
    port map (
            O => \N__34590\,
            I => \N__34583\
        );

    \I__5374\ : InMux
    port map (
            O => \N__34589\,
            I => \N__34580\
        );

    \I__5373\ : Odrv4
    port map (
            O => \N__34586\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__34583\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__34580\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__5370\ : SRMux
    port map (
            O => \N__34573\,
            I => \N__34570\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__34570\,
            I => \N__34567\
        );

    \I__5368\ : Span4Mux_h
    port map (
            O => \N__34567\,
            I => \N__34564\
        );

    \I__5367\ : Span4Mux_v
    port map (
            O => \N__34564\,
            I => \N__34561\
        );

    \I__5366\ : Odrv4
    port map (
            O => \N__34561\,
            I => \c0.n6_adj_3161\
        );

    \I__5365\ : InMux
    port map (
            O => \N__34558\,
            I => \N__34552\
        );

    \I__5364\ : InMux
    port map (
            O => \N__34557\,
            I => \N__34552\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__34552\,
            I => \N__34548\
        );

    \I__5362\ : InMux
    port map (
            O => \N__34551\,
            I => \N__34545\
        );

    \I__5361\ : Span4Mux_v
    port map (
            O => \N__34548\,
            I => \N__34542\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__34545\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__5359\ : Odrv4
    port map (
            O => \N__34542\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__5358\ : SRMux
    port map (
            O => \N__34537\,
            I => \N__34534\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__34534\,
            I => \N__34531\
        );

    \I__5356\ : Span4Mux_v
    port map (
            O => \N__34531\,
            I => \N__34528\
        );

    \I__5355\ : Span4Mux_v
    port map (
            O => \N__34528\,
            I => \N__34525\
        );

    \I__5354\ : Odrv4
    port map (
            O => \N__34525\,
            I => \c0.n6_adj_3172\
        );

    \I__5353\ : SRMux
    port map (
            O => \N__34522\,
            I => \N__34519\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__34519\,
            I => \N__34516\
        );

    \I__5351\ : Span4Mux_h
    port map (
            O => \N__34516\,
            I => \N__34513\
        );

    \I__5350\ : Span4Mux_v
    port map (
            O => \N__34513\,
            I => \N__34510\
        );

    \I__5349\ : Odrv4
    port map (
            O => \N__34510\,
            I => \c0.n6_adj_3194\
        );

    \I__5348\ : InMux
    port map (
            O => \N__34507\,
            I => \N__34501\
        );

    \I__5347\ : InMux
    port map (
            O => \N__34506\,
            I => \N__34501\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__34501\,
            I => \N__34498\
        );

    \I__5345\ : Span4Mux_v
    port map (
            O => \N__34498\,
            I => \N__34494\
        );

    \I__5344\ : InMux
    port map (
            O => \N__34497\,
            I => \N__34491\
        );

    \I__5343\ : Span4Mux_v
    port map (
            O => \N__34494\,
            I => \N__34488\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__34491\,
            I => \c0.FRAME_MATCHER_i_12\
        );

    \I__5341\ : Odrv4
    port map (
            O => \N__34488\,
            I => \c0.FRAME_MATCHER_i_12\
        );

    \I__5340\ : InMux
    port map (
            O => \N__34483\,
            I => \N__34478\
        );

    \I__5339\ : InMux
    port map (
            O => \N__34482\,
            I => \N__34475\
        );

    \I__5338\ : InMux
    port map (
            O => \N__34481\,
            I => \N__34472\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__34478\,
            I => \c0.FRAME_MATCHER_i_20\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__34475\,
            I => \c0.FRAME_MATCHER_i_20\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__34472\,
            I => \c0.FRAME_MATCHER_i_20\
        );

    \I__5334\ : CascadeMux
    port map (
            O => \N__34465\,
            I => \N__34461\
        );

    \I__5333\ : InMux
    port map (
            O => \N__34464\,
            I => \N__34456\
        );

    \I__5332\ : InMux
    port map (
            O => \N__34461\,
            I => \N__34456\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__34456\,
            I => \N__34452\
        );

    \I__5330\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34449\
        );

    \I__5329\ : Span4Mux_v
    port map (
            O => \N__34452\,
            I => \N__34446\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__34449\,
            I => \c0.FRAME_MATCHER_i_14\
        );

    \I__5327\ : Odrv4
    port map (
            O => \N__34446\,
            I => \c0.FRAME_MATCHER_i_14\
        );

    \I__5326\ : InMux
    port map (
            O => \N__34441\,
            I => \N__34437\
        );

    \I__5325\ : InMux
    port map (
            O => \N__34440\,
            I => \N__34434\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__34437\,
            I => \N__34431\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__34434\,
            I => \N__34428\
        );

    \I__5322\ : Span4Mux_v
    port map (
            O => \N__34431\,
            I => \N__34425\
        );

    \I__5321\ : Span12Mux_h
    port map (
            O => \N__34428\,
            I => \N__34421\
        );

    \I__5320\ : Span4Mux_v
    port map (
            O => \N__34425\,
            I => \N__34418\
        );

    \I__5319\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34415\
        );

    \I__5318\ : Span12Mux_v
    port map (
            O => \N__34421\,
            I => \N__34412\
        );

    \I__5317\ : Odrv4
    port map (
            O => \N__34418\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__34415\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__5315\ : Odrv12
    port map (
            O => \N__34412\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__5314\ : SRMux
    port map (
            O => \N__34405\,
            I => \N__34402\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__34402\,
            I => \N__34399\
        );

    \I__5312\ : Span4Mux_v
    port map (
            O => \N__34399\,
            I => \N__34396\
        );

    \I__5311\ : Span4Mux_v
    port map (
            O => \N__34396\,
            I => \N__34393\
        );

    \I__5310\ : Odrv4
    port map (
            O => \N__34393\,
            I => \c0.n6_adj_3160\
        );

    \I__5309\ : InMux
    port map (
            O => \N__34390\,
            I => \N__34387\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__34387\,
            I => \N__34383\
        );

    \I__5307\ : InMux
    port map (
            O => \N__34386\,
            I => \N__34379\
        );

    \I__5306\ : Span4Mux_h
    port map (
            O => \N__34383\,
            I => \N__34376\
        );

    \I__5305\ : InMux
    port map (
            O => \N__34382\,
            I => \N__34373\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__34379\,
            I => \N__34370\
        );

    \I__5303\ : Odrv4
    port map (
            O => \N__34376\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__34373\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__5301\ : Odrv4
    port map (
            O => \N__34370\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__5300\ : CascadeMux
    port map (
            O => \N__34363\,
            I => \N__34360\
        );

    \I__5299\ : InMux
    port map (
            O => \N__34360\,
            I => \N__34357\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__34357\,
            I => \N__34352\
        );

    \I__5297\ : InMux
    port map (
            O => \N__34356\,
            I => \N__34349\
        );

    \I__5296\ : InMux
    port map (
            O => \N__34355\,
            I => \N__34346\
        );

    \I__5295\ : Span4Mux_v
    port map (
            O => \N__34352\,
            I => \N__34343\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__34349\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__34346\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__5292\ : Odrv4
    port map (
            O => \N__34343\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__5291\ : InMux
    port map (
            O => \N__34336\,
            I => \N__34332\
        );

    \I__5290\ : InMux
    port map (
            O => \N__34335\,
            I => \N__34329\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__34332\,
            I => \N__34324\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__34329\,
            I => \N__34324\
        );

    \I__5287\ : Span4Mux_v
    port map (
            O => \N__34324\,
            I => \N__34320\
        );

    \I__5286\ : InMux
    port map (
            O => \N__34323\,
            I => \N__34317\
        );

    \I__5285\ : Span4Mux_v
    port map (
            O => \N__34320\,
            I => \N__34314\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__34317\,
            I => \c0.FRAME_MATCHER_i_11\
        );

    \I__5283\ : Odrv4
    port map (
            O => \N__34314\,
            I => \c0.FRAME_MATCHER_i_11\
        );

    \I__5282\ : InMux
    port map (
            O => \N__34309\,
            I => \N__34306\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__34306\,
            I => n13179
        );

    \I__5280\ : InMux
    port map (
            O => \N__34303\,
            I => \bfn_15_19_0_\
        );

    \I__5279\ : InMux
    port map (
            O => \N__34300\,
            I => \c0.rx.n17267\
        );

    \I__5278\ : InMux
    port map (
            O => \N__34297\,
            I => \N__34294\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__34294\,
            I => n12908
        );

    \I__5276\ : InMux
    port map (
            O => \N__34291\,
            I => \c0.rx.n17268\
        );

    \I__5275\ : InMux
    port map (
            O => \N__34288\,
            I => \c0.rx.n17269\
        );

    \I__5274\ : InMux
    port map (
            O => \N__34285\,
            I => \c0.rx.n17270\
        );

    \I__5273\ : InMux
    port map (
            O => \N__34282\,
            I => \c0.rx.n17271\
        );

    \I__5272\ : InMux
    port map (
            O => \N__34279\,
            I => \c0.rx.n17272\
        );

    \I__5271\ : CascadeMux
    port map (
            O => \N__34276\,
            I => \c0.rx.n14601_cascade_\
        );

    \I__5270\ : InMux
    port map (
            O => \N__34273\,
            I => \N__34270\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__34270\,
            I => \N__34267\
        );

    \I__5268\ : Odrv12
    port map (
            O => \N__34267\,
            I => n12301
        );

    \I__5267\ : InMux
    port map (
            O => \N__34264\,
            I => \N__34261\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__34261\,
            I => \N__34258\
        );

    \I__5265\ : Span4Mux_h
    port map (
            O => \N__34258\,
            I => \N__34255\
        );

    \I__5264\ : Odrv4
    port map (
            O => \N__34255\,
            I => \c0.n15685\
        );

    \I__5263\ : CascadeMux
    port map (
            O => \N__34252\,
            I => \N__34249\
        );

    \I__5262\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34246\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__34246\,
            I => \N__34243\
        );

    \I__5260\ : Span4Mux_h
    port map (
            O => \N__34243\,
            I => \N__34240\
        );

    \I__5259\ : Odrv4
    port map (
            O => \N__34240\,
            I => \c0.rx.n6\
        );

    \I__5258\ : CascadeMux
    port map (
            O => \N__34237\,
            I => \n12492_cascade_\
        );

    \I__5257\ : InMux
    port map (
            O => \N__34234\,
            I => \N__34230\
        );

    \I__5256\ : CascadeMux
    port map (
            O => \N__34233\,
            I => \N__34223\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__34230\,
            I => \N__34217\
        );

    \I__5254\ : InMux
    port map (
            O => \N__34229\,
            I => \N__34212\
        );

    \I__5253\ : InMux
    port map (
            O => \N__34228\,
            I => \N__34212\
        );

    \I__5252\ : InMux
    port map (
            O => \N__34227\,
            I => \N__34209\
        );

    \I__5251\ : InMux
    port map (
            O => \N__34226\,
            I => \N__34204\
        );

    \I__5250\ : InMux
    port map (
            O => \N__34223\,
            I => \N__34204\
        );

    \I__5249\ : InMux
    port map (
            O => \N__34222\,
            I => \N__34197\
        );

    \I__5248\ : InMux
    port map (
            O => \N__34221\,
            I => \N__34197\
        );

    \I__5247\ : InMux
    port map (
            O => \N__34220\,
            I => \N__34197\
        );

    \I__5246\ : Span4Mux_v
    port map (
            O => \N__34217\,
            I => \N__34194\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__34212\,
            I => \c0.r_Bit_Index_0\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__34209\,
            I => \c0.r_Bit_Index_0\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__34204\,
            I => \c0.r_Bit_Index_0\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__34197\,
            I => \c0.r_Bit_Index_0\
        );

    \I__5241\ : Odrv4
    port map (
            O => \N__34194\,
            I => \c0.r_Bit_Index_0\
        );

    \I__5240\ : IoInMux
    port map (
            O => \N__34183\,
            I => \N__34179\
        );

    \I__5239\ : InMux
    port map (
            O => \N__34182\,
            I => \N__34176\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__34179\,
            I => \N__34170\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__34176\,
            I => \N__34170\
        );

    \I__5236\ : InMux
    port map (
            O => \N__34175\,
            I => \N__34165\
        );

    \I__5235\ : Span4Mux_s3_h
    port map (
            O => \N__34170\,
            I => \N__34162\
        );

    \I__5234\ : InMux
    port map (
            O => \N__34169\,
            I => \N__34155\
        );

    \I__5233\ : InMux
    port map (
            O => \N__34168\,
            I => \N__34155\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__34165\,
            I => \N__34152\
        );

    \I__5231\ : Sp12to4
    port map (
            O => \N__34162\,
            I => \N__34149\
        );

    \I__5230\ : InMux
    port map (
            O => \N__34161\,
            I => \N__34146\
        );

    \I__5229\ : InMux
    port map (
            O => \N__34160\,
            I => \N__34143\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__34155\,
            I => \N__34138\
        );

    \I__5227\ : Span4Mux_h
    port map (
            O => \N__34152\,
            I => \N__34138\
        );

    \I__5226\ : Span12Mux_v
    port map (
            O => \N__34149\,
            I => \N__34135\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__34146\,
            I => \N__34130\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__34143\,
            I => \N__34130\
        );

    \I__5223\ : Span4Mux_h
    port map (
            O => \N__34138\,
            I => \N__34127\
        );

    \I__5222\ : Odrv12
    port map (
            O => \N__34135\,
            I => tx_o
        );

    \I__5221\ : Odrv4
    port map (
            O => \N__34130\,
            I => tx_o
        );

    \I__5220\ : Odrv4
    port map (
            O => \N__34127\,
            I => tx_o
        );

    \I__5219\ : CascadeMux
    port map (
            O => \N__34120\,
            I => \N__34116\
        );

    \I__5218\ : CascadeMux
    port map (
            O => \N__34119\,
            I => \N__34113\
        );

    \I__5217\ : InMux
    port map (
            O => \N__34116\,
            I => \N__34110\
        );

    \I__5216\ : InMux
    port map (
            O => \N__34113\,
            I => \N__34107\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__34110\,
            I => \N__34104\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__34107\,
            I => \r_Tx_Data_1\
        );

    \I__5213\ : Odrv4
    port map (
            O => \N__34104\,
            I => \r_Tx_Data_1\
        );

    \I__5212\ : InMux
    port map (
            O => \N__34099\,
            I => \N__34089\
        );

    \I__5211\ : InMux
    port map (
            O => \N__34098\,
            I => \N__34086\
        );

    \I__5210\ : InMux
    port map (
            O => \N__34097\,
            I => \N__34078\
        );

    \I__5209\ : InMux
    port map (
            O => \N__34096\,
            I => \N__34078\
        );

    \I__5208\ : InMux
    port map (
            O => \N__34095\,
            I => \N__34069\
        );

    \I__5207\ : InMux
    port map (
            O => \N__34094\,
            I => \N__34069\
        );

    \I__5206\ : InMux
    port map (
            O => \N__34093\,
            I => \N__34069\
        );

    \I__5205\ : InMux
    port map (
            O => \N__34092\,
            I => \N__34069\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__34089\,
            I => \N__34066\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__34086\,
            I => \N__34056\
        );

    \I__5202\ : InMux
    port map (
            O => \N__34085\,
            I => \N__34053\
        );

    \I__5201\ : InMux
    port map (
            O => \N__34084\,
            I => \N__34050\
        );

    \I__5200\ : InMux
    port map (
            O => \N__34083\,
            I => \N__34047\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__34078\,
            I => \N__34040\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__34069\,
            I => \N__34040\
        );

    \I__5197\ : Span4Mux_h
    port map (
            O => \N__34066\,
            I => \N__34040\
        );

    \I__5196\ : InMux
    port map (
            O => \N__34065\,
            I => \N__34037\
        );

    \I__5195\ : InMux
    port map (
            O => \N__34064\,
            I => \N__34034\
        );

    \I__5194\ : InMux
    port map (
            O => \N__34063\,
            I => \N__34031\
        );

    \I__5193\ : InMux
    port map (
            O => \N__34062\,
            I => \N__34028\
        );

    \I__5192\ : InMux
    port map (
            O => \N__34061\,
            I => \N__34021\
        );

    \I__5191\ : InMux
    port map (
            O => \N__34060\,
            I => \N__34021\
        );

    \I__5190\ : InMux
    port map (
            O => \N__34059\,
            I => \N__34021\
        );

    \I__5189\ : Span4Mux_h
    port map (
            O => \N__34056\,
            I => \N__34018\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__34053\,
            I => \N__34011\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__34050\,
            I => \N__34011\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__34047\,
            I => \N__34011\
        );

    \I__5185\ : Span4Mux_h
    port map (
            O => \N__34040\,
            I => \N__34008\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__34037\,
            I => \c0.r_SM_Main_2\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__34034\,
            I => \c0.r_SM_Main_2\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__34031\,
            I => \c0.r_SM_Main_2\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__34028\,
            I => \c0.r_SM_Main_2\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__34021\,
            I => \c0.r_SM_Main_2\
        );

    \I__5179\ : Odrv4
    port map (
            O => \N__34018\,
            I => \c0.r_SM_Main_2\
        );

    \I__5178\ : Odrv4
    port map (
            O => \N__34011\,
            I => \c0.r_SM_Main_2\
        );

    \I__5177\ : Odrv4
    port map (
            O => \N__34008\,
            I => \c0.r_SM_Main_2\
        );

    \I__5176\ : InMux
    port map (
            O => \N__33991\,
            I => \N__33988\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__33988\,
            I => \N__33985\
        );

    \I__5174\ : Span4Mux_v
    port map (
            O => \N__33985\,
            I => \N__33982\
        );

    \I__5173\ : Odrv4
    port map (
            O => \N__33982\,
            I => \c0.n21611\
        );

    \I__5172\ : InMux
    port map (
            O => \N__33979\,
            I => \N__33976\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__33976\,
            I => \N__33973\
        );

    \I__5170\ : Span4Mux_h
    port map (
            O => \N__33973\,
            I => \N__33970\
        );

    \I__5169\ : Span4Mux_h
    port map (
            O => \N__33970\,
            I => \N__33966\
        );

    \I__5168\ : CascadeMux
    port map (
            O => \N__33969\,
            I => \N__33962\
        );

    \I__5167\ : Span4Mux_v
    port map (
            O => \N__33966\,
            I => \N__33959\
        );

    \I__5166\ : InMux
    port map (
            O => \N__33965\,
            I => \N__33956\
        );

    \I__5165\ : InMux
    port map (
            O => \N__33962\,
            I => \N__33953\
        );

    \I__5164\ : Odrv4
    port map (
            O => \N__33959\,
            I => encoder0_position_23
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__33956\,
            I => encoder0_position_23
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__33953\,
            I => encoder0_position_23
        );

    \I__5161\ : InMux
    port map (
            O => \N__33946\,
            I => \N__33942\
        );

    \I__5160\ : InMux
    port map (
            O => \N__33945\,
            I => \N__33939\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__33942\,
            I => \N__33936\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__33939\,
            I => data_out_frame_7_7
        );

    \I__5157\ : Odrv12
    port map (
            O => \N__33936\,
            I => data_out_frame_7_7
        );

    \I__5156\ : InMux
    port map (
            O => \N__33931\,
            I => \N__33927\
        );

    \I__5155\ : InMux
    port map (
            O => \N__33930\,
            I => \N__33924\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__33927\,
            I => \N__33921\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__33924\,
            I => \r_Tx_Data_7\
        );

    \I__5152\ : Odrv4
    port map (
            O => \N__33921\,
            I => \r_Tx_Data_7\
        );

    \I__5151\ : InMux
    port map (
            O => \N__33916\,
            I => \N__33910\
        );

    \I__5150\ : InMux
    port map (
            O => \N__33915\,
            I => \N__33910\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__33910\,
            I => data_out_frame_7_5
        );

    \I__5148\ : InMux
    port map (
            O => \N__33907\,
            I => \N__33903\
        );

    \I__5147\ : InMux
    port map (
            O => \N__33906\,
            I => \N__33900\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__33903\,
            I => \N__33897\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__33900\,
            I => data_out_frame_6_5
        );

    \I__5144\ : Odrv4
    port map (
            O => \N__33897\,
            I => data_out_frame_6_5
        );

    \I__5143\ : InMux
    port map (
            O => \N__33892\,
            I => \N__33889\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__33889\,
            I => \c0.n5_adj_3447\
        );

    \I__5141\ : CascadeMux
    port map (
            O => \N__33886\,
            I => \N__33882\
        );

    \I__5140\ : CascadeMux
    port map (
            O => \N__33885\,
            I => \N__33874\
        );

    \I__5139\ : InMux
    port map (
            O => \N__33882\,
            I => \N__33870\
        );

    \I__5138\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33865\
        );

    \I__5137\ : InMux
    port map (
            O => \N__33880\,
            I => \N__33865\
        );

    \I__5136\ : InMux
    port map (
            O => \N__33879\,
            I => \N__33862\
        );

    \I__5135\ : CascadeMux
    port map (
            O => \N__33878\,
            I => \N__33858\
        );

    \I__5134\ : CascadeMux
    port map (
            O => \N__33877\,
            I => \N__33855\
        );

    \I__5133\ : InMux
    port map (
            O => \N__33874\,
            I => \N__33852\
        );

    \I__5132\ : InMux
    port map (
            O => \N__33873\,
            I => \N__33849\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__33870\,
            I => \N__33845\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__33865\,
            I => \N__33840\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__33862\,
            I => \N__33840\
        );

    \I__5128\ : InMux
    port map (
            O => \N__33861\,
            I => \N__33835\
        );

    \I__5127\ : InMux
    port map (
            O => \N__33858\,
            I => \N__33835\
        );

    \I__5126\ : InMux
    port map (
            O => \N__33855\,
            I => \N__33832\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__33852\,
            I => \N__33827\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__33849\,
            I => \N__33827\
        );

    \I__5123\ : InMux
    port map (
            O => \N__33848\,
            I => \N__33824\
        );

    \I__5122\ : Span4Mux_h
    port map (
            O => \N__33845\,
            I => \N__33821\
        );

    \I__5121\ : Span4Mux_v
    port map (
            O => \N__33840\,
            I => \N__33818\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__33835\,
            I => byte_transmit_counter_5
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__33832\,
            I => byte_transmit_counter_5
        );

    \I__5118\ : Odrv12
    port map (
            O => \N__33827\,
            I => byte_transmit_counter_5
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__33824\,
            I => byte_transmit_counter_5
        );

    \I__5116\ : Odrv4
    port map (
            O => \N__33821\,
            I => byte_transmit_counter_5
        );

    \I__5115\ : Odrv4
    port map (
            O => \N__33818\,
            I => byte_transmit_counter_5
        );

    \I__5114\ : CascadeMux
    port map (
            O => \N__33805\,
            I => \N__33802\
        );

    \I__5113\ : InMux
    port map (
            O => \N__33802\,
            I => \N__33792\
        );

    \I__5112\ : InMux
    port map (
            O => \N__33801\,
            I => \N__33792\
        );

    \I__5111\ : InMux
    port map (
            O => \N__33800\,
            I => \N__33789\
        );

    \I__5110\ : InMux
    port map (
            O => \N__33799\,
            I => \N__33786\
        );

    \I__5109\ : InMux
    port map (
            O => \N__33798\,
            I => \N__33780\
        );

    \I__5108\ : InMux
    port map (
            O => \N__33797\,
            I => \N__33780\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__33792\,
            I => \N__33775\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__33789\,
            I => \N__33775\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__33786\,
            I => \N__33772\
        );

    \I__5104\ : InMux
    port map (
            O => \N__33785\,
            I => \N__33769\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__33780\,
            I => \N__33766\
        );

    \I__5102\ : Span4Mux_h
    port map (
            O => \N__33775\,
            I => \N__33762\
        );

    \I__5101\ : Span4Mux_h
    port map (
            O => \N__33772\,
            I => \N__33757\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__33769\,
            I => \N__33757\
        );

    \I__5099\ : Span4Mux_h
    port map (
            O => \N__33766\,
            I => \N__33754\
        );

    \I__5098\ : InMux
    port map (
            O => \N__33765\,
            I => \N__33751\
        );

    \I__5097\ : Odrv4
    port map (
            O => \N__33762\,
            I => n9377
        );

    \I__5096\ : Odrv4
    port map (
            O => \N__33757\,
            I => n9377
        );

    \I__5095\ : Odrv4
    port map (
            O => \N__33754\,
            I => n9377
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__33751\,
            I => n9377
        );

    \I__5093\ : CascadeMux
    port map (
            O => \N__33742\,
            I => \N__33739\
        );

    \I__5092\ : InMux
    port map (
            O => \N__33739\,
            I => \N__33736\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__33736\,
            I => \N__33732\
        );

    \I__5090\ : InMux
    port map (
            O => \N__33735\,
            I => \N__33729\
        );

    \I__5089\ : Span4Mux_v
    port map (
            O => \N__33732\,
            I => \N__33726\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__33729\,
            I => data_out_frame_5_5
        );

    \I__5087\ : Odrv4
    port map (
            O => \N__33726\,
            I => data_out_frame_5_5
        );

    \I__5086\ : CascadeMux
    port map (
            O => \N__33721\,
            I => \N__33718\
        );

    \I__5085\ : InMux
    port map (
            O => \N__33718\,
            I => \N__33715\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__33715\,
            I => \c0.n21546\
        );

    \I__5083\ : SRMux
    port map (
            O => \N__33712\,
            I => \N__33709\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__33709\,
            I => \N__33706\
        );

    \I__5081\ : Odrv4
    port map (
            O => \N__33706\,
            I => \c0.n6_adj_3192\
        );

    \I__5080\ : InMux
    port map (
            O => \N__33703\,
            I => \N__33699\
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__33702\,
            I => \N__33696\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__33699\,
            I => \N__33693\
        );

    \I__5077\ : InMux
    port map (
            O => \N__33696\,
            I => \N__33690\
        );

    \I__5076\ : Span4Mux_h
    port map (
            O => \N__33693\,
            I => \N__33686\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__33690\,
            I => \N__33683\
        );

    \I__5074\ : InMux
    port map (
            O => \N__33689\,
            I => \N__33680\
        );

    \I__5073\ : Span4Mux_v
    port map (
            O => \N__33686\,
            I => \N__33675\
        );

    \I__5072\ : Span4Mux_h
    port map (
            O => \N__33683\,
            I => \N__33675\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__33680\,
            I => encoder1_position_1
        );

    \I__5070\ : Odrv4
    port map (
            O => \N__33675\,
            I => encoder1_position_1
        );

    \I__5069\ : InMux
    port map (
            O => \N__33670\,
            I => \N__33666\
        );

    \I__5068\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33663\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__33666\,
            I => \N__33660\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__33663\,
            I => data_out_frame_13_1
        );

    \I__5065\ : Odrv4
    port map (
            O => \N__33660\,
            I => data_out_frame_13_1
        );

    \I__5064\ : SRMux
    port map (
            O => \N__33655\,
            I => \N__33652\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__33652\,
            I => \N__33649\
        );

    \I__5062\ : Odrv4
    port map (
            O => \N__33649\,
            I => \c0.n6_adj_3190\
        );

    \I__5061\ : CascadeMux
    port map (
            O => \N__33646\,
            I => \N__33643\
        );

    \I__5060\ : InMux
    port map (
            O => \N__33643\,
            I => \N__33639\
        );

    \I__5059\ : InMux
    port map (
            O => \N__33642\,
            I => \N__33636\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__33639\,
            I => \N__33633\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__33636\,
            I => data_out_frame_11_2
        );

    \I__5056\ : Odrv12
    port map (
            O => \N__33633\,
            I => data_out_frame_11_2
        );

    \I__5055\ : InMux
    port map (
            O => \N__33628\,
            I => \N__33624\
        );

    \I__5054\ : InMux
    port map (
            O => \N__33627\,
            I => \N__33621\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__33624\,
            I => \N__33616\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__33621\,
            I => \N__33616\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__33616\,
            I => data_out_frame_10_0
        );

    \I__5050\ : CascadeMux
    port map (
            O => \N__33613\,
            I => \N__33610\
        );

    \I__5049\ : InMux
    port map (
            O => \N__33610\,
            I => \N__33607\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__33607\,
            I => \N__33603\
        );

    \I__5047\ : InMux
    port map (
            O => \N__33606\,
            I => \N__33600\
        );

    \I__5046\ : Span12Mux_h
    port map (
            O => \N__33603\,
            I => \N__33597\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__33600\,
            I => data_out_frame_11_0
        );

    \I__5044\ : Odrv12
    port map (
            O => \N__33597\,
            I => data_out_frame_11_0
        );

    \I__5043\ : InMux
    port map (
            O => \N__33592\,
            I => \N__33588\
        );

    \I__5042\ : InMux
    port map (
            O => \N__33591\,
            I => \N__33585\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__33588\,
            I => \N__33582\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__33585\,
            I => data_out_frame_8_0
        );

    \I__5039\ : Odrv4
    port map (
            O => \N__33582\,
            I => data_out_frame_8_0
        );

    \I__5038\ : CascadeMux
    port map (
            O => \N__33577\,
            I => \c0.n21617_cascade_\
        );

    \I__5037\ : InMux
    port map (
            O => \N__33574\,
            I => \N__33570\
        );

    \I__5036\ : InMux
    port map (
            O => \N__33573\,
            I => \N__33567\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__33570\,
            I => \N__33564\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__33567\,
            I => data_out_frame_9_0
        );

    \I__5033\ : Odrv12
    port map (
            O => \N__33564\,
            I => data_out_frame_9_0
        );

    \I__5032\ : CascadeMux
    port map (
            O => \N__33559\,
            I => \c0.n21620_cascade_\
        );

    \I__5031\ : InMux
    port map (
            O => \N__33556\,
            I => \N__33553\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__33553\,
            I => \N__33550\
        );

    \I__5029\ : Span4Mux_h
    port map (
            O => \N__33550\,
            I => \N__33547\
        );

    \I__5028\ : Odrv4
    port map (
            O => \N__33547\,
            I => \c0.n21574\
        );

    \I__5027\ : InMux
    port map (
            O => \N__33544\,
            I => \N__33541\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__33541\,
            I => \N__33537\
        );

    \I__5025\ : InMux
    port map (
            O => \N__33540\,
            I => \N__33534\
        );

    \I__5024\ : Span4Mux_h
    port map (
            O => \N__33537\,
            I => \N__33531\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__33534\,
            I => \c0.byte_transmit_counter_6\
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__33531\,
            I => \c0.byte_transmit_counter_6\
        );

    \I__5021\ : InMux
    port map (
            O => \N__33526\,
            I => \N__33523\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__33523\,
            I => \N__33519\
        );

    \I__5019\ : InMux
    port map (
            O => \N__33522\,
            I => \N__33516\
        );

    \I__5018\ : Span4Mux_h
    port map (
            O => \N__33519\,
            I => \N__33513\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__33516\,
            I => \c0.byte_transmit_counter_7\
        );

    \I__5016\ : Odrv4
    port map (
            O => \N__33513\,
            I => \c0.byte_transmit_counter_7\
        );

    \I__5015\ : InMux
    port map (
            O => \N__33508\,
            I => \N__33502\
        );

    \I__5014\ : InMux
    port map (
            O => \N__33507\,
            I => \N__33502\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__33502\,
            I => \N__33499\
        );

    \I__5012\ : Odrv12
    port map (
            O => \N__33499\,
            I => \c0.n7235\
        );

    \I__5011\ : InMux
    port map (
            O => \N__33496\,
            I => \N__33493\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__33493\,
            I => \N__33490\
        );

    \I__5009\ : Span4Mux_v
    port map (
            O => \N__33490\,
            I => \N__33487\
        );

    \I__5008\ : Span4Mux_v
    port map (
            O => \N__33487\,
            I => \N__33484\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__33484\,
            I => \c0.n2_adj_3147\
        );

    \I__5006\ : SRMux
    port map (
            O => \N__33481\,
            I => \N__33478\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__33478\,
            I => \N__33475\
        );

    \I__5004\ : Span4Mux_h
    port map (
            O => \N__33475\,
            I => \N__33472\
        );

    \I__5003\ : Span4Mux_v
    port map (
            O => \N__33472\,
            I => \N__33469\
        );

    \I__5002\ : Odrv4
    port map (
            O => \N__33469\,
            I => \c0.n6_adj_3151\
        );

    \I__5001\ : InMux
    port map (
            O => \N__33466\,
            I => \N__33463\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__33463\,
            I => \N__33459\
        );

    \I__4999\ : CascadeMux
    port map (
            O => \N__33462\,
            I => \N__33455\
        );

    \I__4998\ : Span12Mux_v
    port map (
            O => \N__33459\,
            I => \N__33452\
        );

    \I__4997\ : InMux
    port map (
            O => \N__33458\,
            I => \N__33449\
        );

    \I__4996\ : InMux
    port map (
            O => \N__33455\,
            I => \N__33446\
        );

    \I__4995\ : Odrv12
    port map (
            O => \N__33452\,
            I => encoder0_position_21
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__33449\,
            I => encoder0_position_21
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__33446\,
            I => encoder0_position_21
        );

    \I__4992\ : InMux
    port map (
            O => \N__33439\,
            I => \N__33436\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__33436\,
            I => \N__33433\
        );

    \I__4990\ : Odrv4
    port map (
            O => \N__33433\,
            I => \c0.n21470\
        );

    \I__4989\ : CascadeMux
    port map (
            O => \N__33430\,
            I => \N__33427\
        );

    \I__4988\ : InMux
    port map (
            O => \N__33427\,
            I => \N__33424\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__33424\,
            I => \N__33421\
        );

    \I__4986\ : Span4Mux_v
    port map (
            O => \N__33421\,
            I => \N__33418\
        );

    \I__4985\ : Span4Mux_h
    port map (
            O => \N__33418\,
            I => \N__33415\
        );

    \I__4984\ : Odrv4
    port map (
            O => \N__33415\,
            I => \c0.n21542\
        );

    \I__4983\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33409\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__33409\,
            I => \N__33406\
        );

    \I__4981\ : Span4Mux_h
    port map (
            O => \N__33406\,
            I => \N__33403\
        );

    \I__4980\ : Odrv4
    port map (
            O => \N__33403\,
            I => n2316
        );

    \I__4979\ : SRMux
    port map (
            O => \N__33400\,
            I => \N__33397\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__33397\,
            I => \N__33394\
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__33394\,
            I => \c0.n6_adj_3156\
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__33391\,
            I => \N__33388\
        );

    \I__4975\ : InMux
    port map (
            O => \N__33388\,
            I => \N__33385\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__33385\,
            I => \N__33380\
        );

    \I__4973\ : InMux
    port map (
            O => \N__33384\,
            I => \N__33375\
        );

    \I__4972\ : InMux
    port map (
            O => \N__33383\,
            I => \N__33375\
        );

    \I__4971\ : Span4Mux_h
    port map (
            O => \N__33380\,
            I => \N__33372\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__33375\,
            I => encoder1_position_29
        );

    \I__4969\ : Odrv4
    port map (
            O => \N__33372\,
            I => encoder1_position_29
        );

    \I__4968\ : InMux
    port map (
            O => \N__33367\,
            I => \N__33363\
        );

    \I__4967\ : InMux
    port map (
            O => \N__33366\,
            I => \N__33360\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__33363\,
            I => data_out_frame_10_5
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__33360\,
            I => data_out_frame_10_5
        );

    \I__4964\ : InMux
    port map (
            O => \N__33355\,
            I => \N__33351\
        );

    \I__4963\ : CascadeMux
    port map (
            O => \N__33354\,
            I => \N__33347\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__33351\,
            I => \N__33344\
        );

    \I__4961\ : InMux
    port map (
            O => \N__33350\,
            I => \N__33341\
        );

    \I__4960\ : InMux
    port map (
            O => \N__33347\,
            I => \N__33338\
        );

    \I__4959\ : Span4Mux_h
    port map (
            O => \N__33344\,
            I => \N__33335\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__33341\,
            I => \N__33330\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__33338\,
            I => \N__33330\
        );

    \I__4956\ : Odrv4
    port map (
            O => \N__33335\,
            I => encoder0_position_29
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__33330\,
            I => encoder0_position_29
        );

    \I__4954\ : InMux
    port map (
            O => \N__33325\,
            I => \N__33322\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__33322\,
            I => \N__33318\
        );

    \I__4952\ : InMux
    port map (
            O => \N__33321\,
            I => \N__33315\
        );

    \I__4951\ : Span4Mux_h
    port map (
            O => \N__33318\,
            I => \N__33312\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__33315\,
            I => \c0.data_out_frame_7_0\
        );

    \I__4949\ : Odrv4
    port map (
            O => \N__33312\,
            I => \c0.data_out_frame_7_0\
        );

    \I__4948\ : InMux
    port map (
            O => \N__33307\,
            I => \N__33304\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__33304\,
            I => \N__33301\
        );

    \I__4946\ : Span4Mux_v
    port map (
            O => \N__33301\,
            I => \N__33298\
        );

    \I__4945\ : Odrv4
    port map (
            O => \N__33298\,
            I => \c0.n17150\
        );

    \I__4944\ : InMux
    port map (
            O => \N__33295\,
            I => \N__33291\
        );

    \I__4943\ : CascadeMux
    port map (
            O => \N__33294\,
            I => \N__33287\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__33291\,
            I => \N__33284\
        );

    \I__4941\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33281\
        );

    \I__4940\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33278\
        );

    \I__4939\ : Span4Mux_v
    port map (
            O => \N__33284\,
            I => \N__33275\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__33281\,
            I => \N__33270\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__33278\,
            I => \N__33270\
        );

    \I__4936\ : Odrv4
    port map (
            O => \N__33275\,
            I => encoder1_position_18
        );

    \I__4935\ : Odrv4
    port map (
            O => \N__33270\,
            I => encoder1_position_18
        );

    \I__4934\ : InMux
    port map (
            O => \N__33265\,
            I => \N__33262\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__33262\,
            I => \N__33259\
        );

    \I__4932\ : Span4Mux_h
    port map (
            O => \N__33259\,
            I => \N__33254\
        );

    \I__4931\ : CascadeMux
    port map (
            O => \N__33258\,
            I => \N__33251\
        );

    \I__4930\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33248\
        );

    \I__4929\ : Span4Mux_h
    port map (
            O => \N__33254\,
            I => \N__33245\
        );

    \I__4928\ : InMux
    port map (
            O => \N__33251\,
            I => \N__33242\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__33248\,
            I => encoder0_position_11
        );

    \I__4926\ : Odrv4
    port map (
            O => \N__33245\,
            I => encoder0_position_11
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__33242\,
            I => encoder0_position_11
        );

    \I__4924\ : InMux
    port map (
            O => \N__33235\,
            I => \N__33232\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__33232\,
            I => \N__33228\
        );

    \I__4922\ : InMux
    port map (
            O => \N__33231\,
            I => \N__33225\
        );

    \I__4921\ : Span4Mux_h
    port map (
            O => \N__33228\,
            I => \N__33222\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__33225\,
            I => data_out_frame_10_7
        );

    \I__4919\ : Odrv4
    port map (
            O => \N__33222\,
            I => data_out_frame_10_7
        );

    \I__4918\ : InMux
    port map (
            O => \N__33217\,
            I => \N__33214\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__33214\,
            I => \N__33211\
        );

    \I__4916\ : Span4Mux_v
    port map (
            O => \N__33211\,
            I => \N__33208\
        );

    \I__4915\ : Odrv4
    port map (
            O => \N__33208\,
            I => \c0.n21623\
        );

    \I__4914\ : InMux
    port map (
            O => \N__33205\,
            I => \N__33201\
        );

    \I__4913\ : InMux
    port map (
            O => \N__33204\,
            I => \N__33198\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__33201\,
            I => \N__33195\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__33198\,
            I => data_out_frame_9_3
        );

    \I__4910\ : Odrv12
    port map (
            O => \N__33195\,
            I => data_out_frame_9_3
        );

    \I__4909\ : InMux
    port map (
            O => \N__33190\,
            I => \N__33187\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__33187\,
            I => \N__33184\
        );

    \I__4907\ : Span4Mux_h
    port map (
            O => \N__33184\,
            I => \N__33181\
        );

    \I__4906\ : Odrv4
    port map (
            O => \N__33181\,
            I => \c0.n21641\
        );

    \I__4905\ : CascadeMux
    port map (
            O => \N__33178\,
            I => \N__33174\
        );

    \I__4904\ : CascadeMux
    port map (
            O => \N__33177\,
            I => \N__33171\
        );

    \I__4903\ : InMux
    port map (
            O => \N__33174\,
            I => \N__33166\
        );

    \I__4902\ : InMux
    port map (
            O => \N__33171\,
            I => \N__33166\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__33166\,
            I => data_out_frame_8_3
        );

    \I__4900\ : InMux
    port map (
            O => \N__33163\,
            I => \N__33160\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__33160\,
            I => \N__33157\
        );

    \I__4898\ : Span4Mux_h
    port map (
            O => \N__33157\,
            I => \N__33154\
        );

    \I__4897\ : Span4Mux_v
    port map (
            O => \N__33154\,
            I => \N__33151\
        );

    \I__4896\ : Odrv4
    port map (
            O => \N__33151\,
            I => \c0.n21644\
        );

    \I__4895\ : CascadeMux
    port map (
            O => \N__33148\,
            I => \N__33145\
        );

    \I__4894\ : InMux
    port map (
            O => \N__33145\,
            I => \N__33142\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__33142\,
            I => \N__33138\
        );

    \I__4892\ : InMux
    port map (
            O => \N__33141\,
            I => \N__33135\
        );

    \I__4891\ : Span4Mux_v
    port map (
            O => \N__33138\,
            I => \N__33132\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__33135\,
            I => data_out_frame_11_5
        );

    \I__4889\ : Odrv4
    port map (
            O => \N__33132\,
            I => data_out_frame_11_5
        );

    \I__4888\ : InMux
    port map (
            O => \N__33127\,
            I => \N__33123\
        );

    \I__4887\ : InMux
    port map (
            O => \N__33126\,
            I => \N__33120\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__33123\,
            I => \N__33117\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__33120\,
            I => data_out_frame_8_5
        );

    \I__4884\ : Odrv12
    port map (
            O => \N__33117\,
            I => data_out_frame_8_5
        );

    \I__4883\ : CascadeMux
    port map (
            O => \N__33112\,
            I => \c0.n21635_cascade_\
        );

    \I__4882\ : InMux
    port map (
            O => \N__33109\,
            I => \N__33106\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__33106\,
            I => \N__33103\
        );

    \I__4880\ : Span4Mux_h
    port map (
            O => \N__33103\,
            I => \N__33099\
        );

    \I__4879\ : InMux
    port map (
            O => \N__33102\,
            I => \N__33096\
        );

    \I__4878\ : Span4Mux_h
    port map (
            O => \N__33099\,
            I => \N__33093\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__33096\,
            I => data_out_frame_9_5
        );

    \I__4876\ : Odrv4
    port map (
            O => \N__33093\,
            I => data_out_frame_9_5
        );

    \I__4875\ : CascadeMux
    port map (
            O => \N__33088\,
            I => \N__33084\
        );

    \I__4874\ : InMux
    port map (
            O => \N__33087\,
            I => \N__33081\
        );

    \I__4873\ : InMux
    port map (
            O => \N__33084\,
            I => \N__33078\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__33081\,
            I => data_out_frame_5_3
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__33078\,
            I => data_out_frame_5_3
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__33073\,
            I => \N__33070\
        );

    \I__4869\ : InMux
    port map (
            O => \N__33070\,
            I => \N__33067\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__33067\,
            I => \N__33064\
        );

    \I__4867\ : Span4Mux_h
    port map (
            O => \N__33064\,
            I => \N__33060\
        );

    \I__4866\ : InMux
    port map (
            O => \N__33063\,
            I => \N__33057\
        );

    \I__4865\ : Span4Mux_v
    port map (
            O => \N__33060\,
            I => \N__33054\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__33057\,
            I => data_out_frame_28_4
        );

    \I__4863\ : Odrv4
    port map (
            O => \N__33054\,
            I => data_out_frame_28_4
        );

    \I__4862\ : InMux
    port map (
            O => \N__33049\,
            I => \N__33046\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__33046\,
            I => \N__33043\
        );

    \I__4860\ : Span4Mux_v
    port map (
            O => \N__33043\,
            I => \N__33040\
        );

    \I__4859\ : Odrv4
    port map (
            O => \N__33040\,
            I => n2342
        );

    \I__4858\ : CascadeMux
    port map (
            O => \N__33037\,
            I => \N__33033\
        );

    \I__4857\ : InMux
    port map (
            O => \N__33036\,
            I => \N__33030\
        );

    \I__4856\ : InMux
    port map (
            O => \N__33033\,
            I => \N__33027\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__33030\,
            I => \N__33024\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__33027\,
            I => \N__33020\
        );

    \I__4853\ : Span4Mux_v
    port map (
            O => \N__33024\,
            I => \N__33017\
        );

    \I__4852\ : InMux
    port map (
            O => \N__33023\,
            I => \N__33014\
        );

    \I__4851\ : Span4Mux_h
    port map (
            O => \N__33020\,
            I => \N__33011\
        );

    \I__4850\ : Odrv4
    port map (
            O => \N__33017\,
            I => encoder1_position_3
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__33014\,
            I => encoder1_position_3
        );

    \I__4848\ : Odrv4
    port map (
            O => \N__33011\,
            I => encoder1_position_3
        );

    \I__4847\ : InMux
    port map (
            O => \N__33004\,
            I => \N__32999\
        );

    \I__4846\ : CascadeMux
    port map (
            O => \N__33003\,
            I => \N__32996\
        );

    \I__4845\ : InMux
    port map (
            O => \N__33002\,
            I => \N__32993\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__32999\,
            I => \N__32990\
        );

    \I__4843\ : InMux
    port map (
            O => \N__32996\,
            I => \N__32987\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__32993\,
            I => encoder0_position_19
        );

    \I__4841\ : Odrv12
    port map (
            O => \N__32990\,
            I => encoder0_position_19
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__32987\,
            I => encoder0_position_19
        );

    \I__4839\ : CascadeMux
    port map (
            O => \N__32980\,
            I => \c0.n6_adj_3379_cascade_\
        );

    \I__4838\ : InMux
    port map (
            O => \N__32977\,
            I => \N__32974\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__32974\,
            I => \N__32971\
        );

    \I__4836\ : Span4Mux_h
    port map (
            O => \N__32971\,
            I => \N__32968\
        );

    \I__4835\ : Odrv4
    port map (
            O => \N__32968\,
            I => n2324
        );

    \I__4834\ : CascadeMux
    port map (
            O => \N__32965\,
            I => \N__32961\
        );

    \I__4833\ : InMux
    port map (
            O => \N__32964\,
            I => \N__32958\
        );

    \I__4832\ : InMux
    port map (
            O => \N__32961\,
            I => \N__32954\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__32958\,
            I => \N__32951\
        );

    \I__4830\ : InMux
    port map (
            O => \N__32957\,
            I => \N__32948\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__32954\,
            I => \N__32945\
        );

    \I__4828\ : Odrv4
    port map (
            O => \N__32951\,
            I => encoder1_position_21
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__32948\,
            I => encoder1_position_21
        );

    \I__4826\ : Odrv4
    port map (
            O => \N__32945\,
            I => encoder1_position_21
        );

    \I__4825\ : InMux
    port map (
            O => \N__32938\,
            I => \N__32935\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__32935\,
            I => \N__32932\
        );

    \I__4823\ : Span4Mux_h
    port map (
            O => \N__32932\,
            I => \N__32929\
        );

    \I__4822\ : Span4Mux_h
    port map (
            O => \N__32929\,
            I => \N__32926\
        );

    \I__4821\ : Odrv4
    port map (
            O => \N__32926\,
            I => \c0.n21559\
        );

    \I__4820\ : InMux
    port map (
            O => \N__32923\,
            I => \N__32920\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__32920\,
            I => \N__32917\
        );

    \I__4818\ : Span4Mux_h
    port map (
            O => \N__32917\,
            I => \N__32914\
        );

    \I__4817\ : Odrv4
    port map (
            O => \N__32914\,
            I => \c0.n5_adj_3102\
        );

    \I__4816\ : InMux
    port map (
            O => \N__32911\,
            I => \N__32908\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__32908\,
            I => \N__32905\
        );

    \I__4814\ : Span4Mux_v
    port map (
            O => \N__32905\,
            I => \N__32902\
        );

    \I__4813\ : Span4Mux_v
    port map (
            O => \N__32902\,
            I => \N__32899\
        );

    \I__4812\ : Odrv4
    port map (
            O => \N__32899\,
            I => n2322
        );

    \I__4811\ : InMux
    port map (
            O => \N__32896\,
            I => \N__32893\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__32893\,
            I => \N__32890\
        );

    \I__4809\ : Span4Mux_h
    port map (
            O => \N__32890\,
            I => \N__32886\
        );

    \I__4808\ : CascadeMux
    port map (
            O => \N__32889\,
            I => \N__32882\
        );

    \I__4807\ : Span4Mux_h
    port map (
            O => \N__32886\,
            I => \N__32879\
        );

    \I__4806\ : InMux
    port map (
            O => \N__32885\,
            I => \N__32876\
        );

    \I__4805\ : InMux
    port map (
            O => \N__32882\,
            I => \N__32873\
        );

    \I__4804\ : Odrv4
    port map (
            O => \N__32879\,
            I => encoder0_position_24
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__32876\,
            I => encoder0_position_24
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__32873\,
            I => encoder0_position_24
        );

    \I__4801\ : InMux
    port map (
            O => \N__32866\,
            I => \N__32863\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__32863\,
            I => \N__32860\
        );

    \I__4799\ : Odrv4
    port map (
            O => \N__32860\,
            I => n2340
        );

    \I__4798\ : InMux
    port map (
            O => \N__32857\,
            I => \N__32854\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__32854\,
            I => \N__32850\
        );

    \I__4796\ : CascadeMux
    port map (
            O => \N__32853\,
            I => \N__32847\
        );

    \I__4795\ : Span4Mux_h
    port map (
            O => \N__32850\,
            I => \N__32844\
        );

    \I__4794\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32840\
        );

    \I__4793\ : Sp12to4
    port map (
            O => \N__32844\,
            I => \N__32837\
        );

    \I__4792\ : InMux
    port map (
            O => \N__32843\,
            I => \N__32834\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__32840\,
            I => \N__32831\
        );

    \I__4790\ : Odrv12
    port map (
            O => \N__32837\,
            I => encoder1_position_5
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__32834\,
            I => encoder1_position_5
        );

    \I__4788\ : Odrv4
    port map (
            O => \N__32831\,
            I => encoder1_position_5
        );

    \I__4787\ : CascadeMux
    port map (
            O => \N__32824\,
            I => \N__32821\
        );

    \I__4786\ : InMux
    port map (
            O => \N__32821\,
            I => \N__32818\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__32818\,
            I => \N__32815\
        );

    \I__4784\ : Span4Mux_h
    port map (
            O => \N__32815\,
            I => \N__32812\
        );

    \I__4783\ : Span4Mux_h
    port map (
            O => \N__32812\,
            I => \N__32809\
        );

    \I__4782\ : Odrv4
    port map (
            O => \N__32809\,
            I => \c0.n21647\
        );

    \I__4781\ : InMux
    port map (
            O => \N__32806\,
            I => \N__32803\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__32803\,
            I => \N__32800\
        );

    \I__4779\ : Span4Mux_v
    port map (
            O => \N__32800\,
            I => \N__32795\
        );

    \I__4778\ : InMux
    port map (
            O => \N__32799\,
            I => \N__32792\
        );

    \I__4777\ : InMux
    port map (
            O => \N__32798\,
            I => \N__32789\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__32795\,
            I => encoder1_position_26
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__32792\,
            I => encoder1_position_26
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__32789\,
            I => encoder1_position_26
        );

    \I__4773\ : InMux
    port map (
            O => \N__32782\,
            I => \N__32776\
        );

    \I__4772\ : InMux
    port map (
            O => \N__32781\,
            I => \N__32776\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__32776\,
            I => data_out_frame_10_2
        );

    \I__4770\ : SRMux
    port map (
            O => \N__32773\,
            I => \N__32770\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__32770\,
            I => \N__32767\
        );

    \I__4768\ : Odrv4
    port map (
            O => \N__32767\,
            I => \c0.n6_adj_3154\
        );

    \I__4767\ : InMux
    port map (
            O => \N__32764\,
            I => \N__32760\
        );

    \I__4766\ : InMux
    port map (
            O => \N__32763\,
            I => \N__32757\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__32760\,
            I => \N__32754\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__32757\,
            I => data_out_frame_6_0
        );

    \I__4763\ : Odrv4
    port map (
            O => \N__32754\,
            I => data_out_frame_6_0
        );

    \I__4762\ : InMux
    port map (
            O => \N__32749\,
            I => \N__32746\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__32746\,
            I => \N__32743\
        );

    \I__4760\ : Span4Mux_h
    port map (
            O => \N__32743\,
            I => \N__32740\
        );

    \I__4759\ : Odrv4
    port map (
            O => \N__32740\,
            I => \c0.n6_adj_3321\
        );

    \I__4758\ : InMux
    port map (
            O => \N__32737\,
            I => \N__32734\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__32734\,
            I => \N__32731\
        );

    \I__4756\ : Span4Mux_h
    port map (
            O => \N__32731\,
            I => \N__32728\
        );

    \I__4755\ : Odrv4
    port map (
            O => \N__32728\,
            I => n2344
        );

    \I__4754\ : InMux
    port map (
            O => \N__32725\,
            I => \N__32688\
        );

    \I__4753\ : InMux
    port map (
            O => \N__32724\,
            I => \N__32688\
        );

    \I__4752\ : InMux
    port map (
            O => \N__32723\,
            I => \N__32688\
        );

    \I__4751\ : InMux
    port map (
            O => \N__32722\,
            I => \N__32679\
        );

    \I__4750\ : InMux
    port map (
            O => \N__32721\,
            I => \N__32679\
        );

    \I__4749\ : InMux
    port map (
            O => \N__32720\,
            I => \N__32679\
        );

    \I__4748\ : InMux
    port map (
            O => \N__32719\,
            I => \N__32679\
        );

    \I__4747\ : InMux
    port map (
            O => \N__32718\,
            I => \N__32672\
        );

    \I__4746\ : InMux
    port map (
            O => \N__32717\,
            I => \N__32672\
        );

    \I__4745\ : InMux
    port map (
            O => \N__32716\,
            I => \N__32672\
        );

    \I__4744\ : InMux
    port map (
            O => \N__32715\,
            I => \N__32663\
        );

    \I__4743\ : InMux
    port map (
            O => \N__32714\,
            I => \N__32663\
        );

    \I__4742\ : InMux
    port map (
            O => \N__32713\,
            I => \N__32663\
        );

    \I__4741\ : InMux
    port map (
            O => \N__32712\,
            I => \N__32663\
        );

    \I__4740\ : InMux
    port map (
            O => \N__32711\,
            I => \N__32656\
        );

    \I__4739\ : InMux
    port map (
            O => \N__32710\,
            I => \N__32656\
        );

    \I__4738\ : InMux
    port map (
            O => \N__32709\,
            I => \N__32656\
        );

    \I__4737\ : InMux
    port map (
            O => \N__32708\,
            I => \N__32647\
        );

    \I__4736\ : InMux
    port map (
            O => \N__32707\,
            I => \N__32647\
        );

    \I__4735\ : InMux
    port map (
            O => \N__32706\,
            I => \N__32647\
        );

    \I__4734\ : InMux
    port map (
            O => \N__32705\,
            I => \N__32647\
        );

    \I__4733\ : CascadeMux
    port map (
            O => \N__32704\,
            I => \N__32615\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__32703\,
            I => \N__32610\
        );

    \I__4731\ : CascadeMux
    port map (
            O => \N__32702\,
            I => \N__32606\
        );

    \I__4730\ : CascadeMux
    port map (
            O => \N__32701\,
            I => \N__32602\
        );

    \I__4729\ : CascadeMux
    port map (
            O => \N__32700\,
            I => \N__32597\
        );

    \I__4728\ : CascadeMux
    port map (
            O => \N__32699\,
            I => \N__32593\
        );

    \I__4727\ : CascadeMux
    port map (
            O => \N__32698\,
            I => \N__32589\
        );

    \I__4726\ : CascadeMux
    port map (
            O => \N__32697\,
            I => \N__32575\
        );

    \I__4725\ : CascadeMux
    port map (
            O => \N__32696\,
            I => \N__32571\
        );

    \I__4724\ : CascadeMux
    port map (
            O => \N__32695\,
            I => \N__32567\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__32688\,
            I => \N__32550\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__32679\,
            I => \N__32550\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__32672\,
            I => \N__32550\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__32663\,
            I => \N__32550\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__32656\,
            I => \N__32550\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__32647\,
            I => \N__32550\
        );

    \I__4717\ : InMux
    port map (
            O => \N__32646\,
            I => \N__32543\
        );

    \I__4716\ : InMux
    port map (
            O => \N__32645\,
            I => \N__32543\
        );

    \I__4715\ : InMux
    port map (
            O => \N__32644\,
            I => \N__32543\
        );

    \I__4714\ : InMux
    port map (
            O => \N__32643\,
            I => \N__32534\
        );

    \I__4713\ : InMux
    port map (
            O => \N__32642\,
            I => \N__32534\
        );

    \I__4712\ : InMux
    port map (
            O => \N__32641\,
            I => \N__32534\
        );

    \I__4711\ : InMux
    port map (
            O => \N__32640\,
            I => \N__32534\
        );

    \I__4710\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32527\
        );

    \I__4709\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32527\
        );

    \I__4708\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32527\
        );

    \I__4707\ : InMux
    port map (
            O => \N__32636\,
            I => \N__32518\
        );

    \I__4706\ : InMux
    port map (
            O => \N__32635\,
            I => \N__32518\
        );

    \I__4705\ : InMux
    port map (
            O => \N__32634\,
            I => \N__32518\
        );

    \I__4704\ : InMux
    port map (
            O => \N__32633\,
            I => \N__32518\
        );

    \I__4703\ : InMux
    port map (
            O => \N__32632\,
            I => \N__32511\
        );

    \I__4702\ : InMux
    port map (
            O => \N__32631\,
            I => \N__32511\
        );

    \I__4701\ : InMux
    port map (
            O => \N__32630\,
            I => \N__32511\
        );

    \I__4700\ : InMux
    port map (
            O => \N__32629\,
            I => \N__32502\
        );

    \I__4699\ : InMux
    port map (
            O => \N__32628\,
            I => \N__32502\
        );

    \I__4698\ : InMux
    port map (
            O => \N__32627\,
            I => \N__32502\
        );

    \I__4697\ : InMux
    port map (
            O => \N__32626\,
            I => \N__32502\
        );

    \I__4696\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32495\
        );

    \I__4695\ : InMux
    port map (
            O => \N__32624\,
            I => \N__32495\
        );

    \I__4694\ : InMux
    port map (
            O => \N__32623\,
            I => \N__32495\
        );

    \I__4693\ : InMux
    port map (
            O => \N__32622\,
            I => \N__32486\
        );

    \I__4692\ : InMux
    port map (
            O => \N__32621\,
            I => \N__32486\
        );

    \I__4691\ : InMux
    port map (
            O => \N__32620\,
            I => \N__32486\
        );

    \I__4690\ : InMux
    port map (
            O => \N__32619\,
            I => \N__32486\
        );

    \I__4689\ : InMux
    port map (
            O => \N__32618\,
            I => \N__32451\
        );

    \I__4688\ : InMux
    port map (
            O => \N__32615\,
            I => \N__32451\
        );

    \I__4687\ : InMux
    port map (
            O => \N__32614\,
            I => \N__32451\
        );

    \I__4686\ : InMux
    port map (
            O => \N__32613\,
            I => \N__32436\
        );

    \I__4685\ : InMux
    port map (
            O => \N__32610\,
            I => \N__32436\
        );

    \I__4684\ : InMux
    port map (
            O => \N__32609\,
            I => \N__32436\
        );

    \I__4683\ : InMux
    port map (
            O => \N__32606\,
            I => \N__32436\
        );

    \I__4682\ : InMux
    port map (
            O => \N__32605\,
            I => \N__32436\
        );

    \I__4681\ : InMux
    port map (
            O => \N__32602\,
            I => \N__32436\
        );

    \I__4680\ : InMux
    port map (
            O => \N__32601\,
            I => \N__32436\
        );

    \I__4679\ : InMux
    port map (
            O => \N__32600\,
            I => \N__32421\
        );

    \I__4678\ : InMux
    port map (
            O => \N__32597\,
            I => \N__32421\
        );

    \I__4677\ : InMux
    port map (
            O => \N__32596\,
            I => \N__32421\
        );

    \I__4676\ : InMux
    port map (
            O => \N__32593\,
            I => \N__32421\
        );

    \I__4675\ : InMux
    port map (
            O => \N__32592\,
            I => \N__32421\
        );

    \I__4674\ : InMux
    port map (
            O => \N__32589\,
            I => \N__32421\
        );

    \I__4673\ : InMux
    port map (
            O => \N__32588\,
            I => \N__32421\
        );

    \I__4672\ : CascadeMux
    port map (
            O => \N__32587\,
            I => \N__32417\
        );

    \I__4671\ : CascadeMux
    port map (
            O => \N__32586\,
            I => \N__32413\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__32585\,
            I => \N__32409\
        );

    \I__4669\ : CascadeMux
    port map (
            O => \N__32584\,
            I => \N__32404\
        );

    \I__4668\ : CascadeMux
    port map (
            O => \N__32583\,
            I => \N__32400\
        );

    \I__4667\ : CascadeMux
    port map (
            O => \N__32582\,
            I => \N__32396\
        );

    \I__4666\ : CascadeMux
    port map (
            O => \N__32581\,
            I => \N__32391\
        );

    \I__4665\ : CascadeMux
    port map (
            O => \N__32580\,
            I => \N__32387\
        );

    \I__4664\ : CascadeMux
    port map (
            O => \N__32579\,
            I => \N__32383\
        );

    \I__4663\ : InMux
    port map (
            O => \N__32578\,
            I => \N__32361\
        );

    \I__4662\ : InMux
    port map (
            O => \N__32575\,
            I => \N__32361\
        );

    \I__4661\ : InMux
    port map (
            O => \N__32574\,
            I => \N__32361\
        );

    \I__4660\ : InMux
    port map (
            O => \N__32571\,
            I => \N__32361\
        );

    \I__4659\ : InMux
    port map (
            O => \N__32570\,
            I => \N__32361\
        );

    \I__4658\ : InMux
    port map (
            O => \N__32567\,
            I => \N__32361\
        );

    \I__4657\ : InMux
    port map (
            O => \N__32566\,
            I => \N__32361\
        );

    \I__4656\ : CascadeMux
    port map (
            O => \N__32565\,
            I => \N__32357\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__32564\,
            I => \N__32353\
        );

    \I__4654\ : CascadeMux
    port map (
            O => \N__32563\,
            I => \N__32349\
        );

    \I__4653\ : Span4Mux_v
    port map (
            O => \N__32550\,
            I => \N__32329\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__32543\,
            I => \N__32329\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__32534\,
            I => \N__32329\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__32527\,
            I => \N__32329\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__32518\,
            I => \N__32329\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__32511\,
            I => \N__32329\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__32502\,
            I => \N__32329\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__32495\,
            I => \N__32329\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__32486\,
            I => \N__32329\
        );

    \I__4644\ : InMux
    port map (
            O => \N__32485\,
            I => \N__32322\
        );

    \I__4643\ : InMux
    port map (
            O => \N__32484\,
            I => \N__32322\
        );

    \I__4642\ : InMux
    port map (
            O => \N__32483\,
            I => \N__32322\
        );

    \I__4641\ : InMux
    port map (
            O => \N__32482\,
            I => \N__32313\
        );

    \I__4640\ : InMux
    port map (
            O => \N__32481\,
            I => \N__32313\
        );

    \I__4639\ : InMux
    port map (
            O => \N__32480\,
            I => \N__32313\
        );

    \I__4638\ : InMux
    port map (
            O => \N__32479\,
            I => \N__32313\
        );

    \I__4637\ : InMux
    port map (
            O => \N__32478\,
            I => \N__32306\
        );

    \I__4636\ : InMux
    port map (
            O => \N__32477\,
            I => \N__32306\
        );

    \I__4635\ : InMux
    port map (
            O => \N__32476\,
            I => \N__32306\
        );

    \I__4634\ : InMux
    port map (
            O => \N__32475\,
            I => \N__32297\
        );

    \I__4633\ : InMux
    port map (
            O => \N__32474\,
            I => \N__32297\
        );

    \I__4632\ : InMux
    port map (
            O => \N__32473\,
            I => \N__32297\
        );

    \I__4631\ : InMux
    port map (
            O => \N__32472\,
            I => \N__32297\
        );

    \I__4630\ : InMux
    port map (
            O => \N__32471\,
            I => \N__32290\
        );

    \I__4629\ : InMux
    port map (
            O => \N__32470\,
            I => \N__32290\
        );

    \I__4628\ : InMux
    port map (
            O => \N__32469\,
            I => \N__32290\
        );

    \I__4627\ : InMux
    port map (
            O => \N__32468\,
            I => \N__32281\
        );

    \I__4626\ : InMux
    port map (
            O => \N__32467\,
            I => \N__32281\
        );

    \I__4625\ : InMux
    port map (
            O => \N__32466\,
            I => \N__32281\
        );

    \I__4624\ : InMux
    port map (
            O => \N__32465\,
            I => \N__32281\
        );

    \I__4623\ : InMux
    port map (
            O => \N__32464\,
            I => \N__32274\
        );

    \I__4622\ : InMux
    port map (
            O => \N__32463\,
            I => \N__32274\
        );

    \I__4621\ : InMux
    port map (
            O => \N__32462\,
            I => \N__32274\
        );

    \I__4620\ : InMux
    port map (
            O => \N__32461\,
            I => \N__32265\
        );

    \I__4619\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32265\
        );

    \I__4618\ : InMux
    port map (
            O => \N__32459\,
            I => \N__32265\
        );

    \I__4617\ : InMux
    port map (
            O => \N__32458\,
            I => \N__32265\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__32451\,
            I => \N__32251\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__32436\,
            I => \N__32251\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__32421\,
            I => \N__32251\
        );

    \I__4613\ : InMux
    port map (
            O => \N__32420\,
            I => \N__32236\
        );

    \I__4612\ : InMux
    port map (
            O => \N__32417\,
            I => \N__32236\
        );

    \I__4611\ : InMux
    port map (
            O => \N__32416\,
            I => \N__32236\
        );

    \I__4610\ : InMux
    port map (
            O => \N__32413\,
            I => \N__32236\
        );

    \I__4609\ : InMux
    port map (
            O => \N__32412\,
            I => \N__32236\
        );

    \I__4608\ : InMux
    port map (
            O => \N__32409\,
            I => \N__32236\
        );

    \I__4607\ : InMux
    port map (
            O => \N__32408\,
            I => \N__32236\
        );

    \I__4606\ : InMux
    port map (
            O => \N__32407\,
            I => \N__32221\
        );

    \I__4605\ : InMux
    port map (
            O => \N__32404\,
            I => \N__32221\
        );

    \I__4604\ : InMux
    port map (
            O => \N__32403\,
            I => \N__32221\
        );

    \I__4603\ : InMux
    port map (
            O => \N__32400\,
            I => \N__32221\
        );

    \I__4602\ : InMux
    port map (
            O => \N__32399\,
            I => \N__32221\
        );

    \I__4601\ : InMux
    port map (
            O => \N__32396\,
            I => \N__32221\
        );

    \I__4600\ : InMux
    port map (
            O => \N__32395\,
            I => \N__32221\
        );

    \I__4599\ : InMux
    port map (
            O => \N__32394\,
            I => \N__32206\
        );

    \I__4598\ : InMux
    port map (
            O => \N__32391\,
            I => \N__32206\
        );

    \I__4597\ : InMux
    port map (
            O => \N__32390\,
            I => \N__32206\
        );

    \I__4596\ : InMux
    port map (
            O => \N__32387\,
            I => \N__32206\
        );

    \I__4595\ : InMux
    port map (
            O => \N__32386\,
            I => \N__32206\
        );

    \I__4594\ : InMux
    port map (
            O => \N__32383\,
            I => \N__32206\
        );

    \I__4593\ : InMux
    port map (
            O => \N__32382\,
            I => \N__32206\
        );

    \I__4592\ : CascadeMux
    port map (
            O => \N__32381\,
            I => \N__32202\
        );

    \I__4591\ : CascadeMux
    port map (
            O => \N__32380\,
            I => \N__32198\
        );

    \I__4590\ : CascadeMux
    port map (
            O => \N__32379\,
            I => \N__32194\
        );

    \I__4589\ : CascadeMux
    port map (
            O => \N__32378\,
            I => \N__32189\
        );

    \I__4588\ : CascadeMux
    port map (
            O => \N__32377\,
            I => \N__32185\
        );

    \I__4587\ : CascadeMux
    port map (
            O => \N__32376\,
            I => \N__32181\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__32361\,
            I => \N__32177\
        );

    \I__4585\ : InMux
    port map (
            O => \N__32360\,
            I => \N__32162\
        );

    \I__4584\ : InMux
    port map (
            O => \N__32357\,
            I => \N__32162\
        );

    \I__4583\ : InMux
    port map (
            O => \N__32356\,
            I => \N__32162\
        );

    \I__4582\ : InMux
    port map (
            O => \N__32353\,
            I => \N__32162\
        );

    \I__4581\ : InMux
    port map (
            O => \N__32352\,
            I => \N__32162\
        );

    \I__4580\ : InMux
    port map (
            O => \N__32349\,
            I => \N__32162\
        );

    \I__4579\ : InMux
    port map (
            O => \N__32348\,
            I => \N__32162\
        );

    \I__4578\ : Span4Mux_v
    port map (
            O => \N__32329\,
            I => \N__32129\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__32322\,
            I => \N__32129\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__32313\,
            I => \N__32129\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__32306\,
            I => \N__32129\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__32297\,
            I => \N__32129\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__32290\,
            I => \N__32129\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__32281\,
            I => \N__32129\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__32274\,
            I => \N__32129\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__32265\,
            I => \N__32129\
        );

    \I__4569\ : InMux
    port map (
            O => \N__32264\,
            I => \N__32122\
        );

    \I__4568\ : InMux
    port map (
            O => \N__32263\,
            I => \N__32122\
        );

    \I__4567\ : InMux
    port map (
            O => \N__32262\,
            I => \N__32122\
        );

    \I__4566\ : InMux
    port map (
            O => \N__32261\,
            I => \N__32113\
        );

    \I__4565\ : InMux
    port map (
            O => \N__32260\,
            I => \N__32113\
        );

    \I__4564\ : InMux
    port map (
            O => \N__32259\,
            I => \N__32113\
        );

    \I__4563\ : InMux
    port map (
            O => \N__32258\,
            I => \N__32113\
        );

    \I__4562\ : Span4Mux_v
    port map (
            O => \N__32251\,
            I => \N__32104\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__32236\,
            I => \N__32104\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__32221\,
            I => \N__32104\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__32206\,
            I => \N__32104\
        );

    \I__4558\ : InMux
    port map (
            O => \N__32205\,
            I => \N__32089\
        );

    \I__4557\ : InMux
    port map (
            O => \N__32202\,
            I => \N__32089\
        );

    \I__4556\ : InMux
    port map (
            O => \N__32201\,
            I => \N__32089\
        );

    \I__4555\ : InMux
    port map (
            O => \N__32198\,
            I => \N__32089\
        );

    \I__4554\ : InMux
    port map (
            O => \N__32197\,
            I => \N__32089\
        );

    \I__4553\ : InMux
    port map (
            O => \N__32194\,
            I => \N__32089\
        );

    \I__4552\ : InMux
    port map (
            O => \N__32193\,
            I => \N__32089\
        );

    \I__4551\ : InMux
    port map (
            O => \N__32192\,
            I => \N__32074\
        );

    \I__4550\ : InMux
    port map (
            O => \N__32189\,
            I => \N__32074\
        );

    \I__4549\ : InMux
    port map (
            O => \N__32188\,
            I => \N__32074\
        );

    \I__4548\ : InMux
    port map (
            O => \N__32185\,
            I => \N__32074\
        );

    \I__4547\ : InMux
    port map (
            O => \N__32184\,
            I => \N__32074\
        );

    \I__4546\ : InMux
    port map (
            O => \N__32181\,
            I => \N__32074\
        );

    \I__4545\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32074\
        );

    \I__4544\ : Span4Mux_v
    port map (
            O => \N__32177\,
            I => \N__32066\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__32162\,
            I => \N__32066\
        );

    \I__4542\ : InMux
    port map (
            O => \N__32161\,
            I => \N__32059\
        );

    \I__4541\ : InMux
    port map (
            O => \N__32160\,
            I => \N__32059\
        );

    \I__4540\ : InMux
    port map (
            O => \N__32159\,
            I => \N__32059\
        );

    \I__4539\ : InMux
    port map (
            O => \N__32158\,
            I => \N__32050\
        );

    \I__4538\ : InMux
    port map (
            O => \N__32157\,
            I => \N__32050\
        );

    \I__4537\ : InMux
    port map (
            O => \N__32156\,
            I => \N__32050\
        );

    \I__4536\ : InMux
    port map (
            O => \N__32155\,
            I => \N__32050\
        );

    \I__4535\ : InMux
    port map (
            O => \N__32154\,
            I => \N__32043\
        );

    \I__4534\ : InMux
    port map (
            O => \N__32153\,
            I => \N__32043\
        );

    \I__4533\ : InMux
    port map (
            O => \N__32152\,
            I => \N__32043\
        );

    \I__4532\ : InMux
    port map (
            O => \N__32151\,
            I => \N__32034\
        );

    \I__4531\ : InMux
    port map (
            O => \N__32150\,
            I => \N__32034\
        );

    \I__4530\ : InMux
    port map (
            O => \N__32149\,
            I => \N__32034\
        );

    \I__4529\ : InMux
    port map (
            O => \N__32148\,
            I => \N__32034\
        );

    \I__4528\ : Span4Mux_v
    port map (
            O => \N__32129\,
            I => \N__32027\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__32122\,
            I => \N__32027\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__32113\,
            I => \N__32027\
        );

    \I__4525\ : Span4Mux_v
    port map (
            O => \N__32104\,
            I => \N__32020\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__32089\,
            I => \N__32020\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__32074\,
            I => \N__32020\
        );

    \I__4522\ : CascadeMux
    port map (
            O => \N__32073\,
            I => \N__32009\
        );

    \I__4521\ : CascadeMux
    port map (
            O => \N__32072\,
            I => \N__32005\
        );

    \I__4520\ : CascadeMux
    port map (
            O => \N__32071\,
            I => \N__32001\
        );

    \I__4519\ : Span4Mux_v
    port map (
            O => \N__32066\,
            I => \N__31982\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__32059\,
            I => \N__31982\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__32050\,
            I => \N__31982\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__32043\,
            I => \N__31982\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__32034\,
            I => \N__31982\
        );

    \I__4514\ : Span4Mux_v
    port map (
            O => \N__32027\,
            I => \N__31977\
        );

    \I__4513\ : Span4Mux_v
    port map (
            O => \N__32020\,
            I => \N__31977\
        );

    \I__4512\ : InMux
    port map (
            O => \N__32019\,
            I => \N__31970\
        );

    \I__4511\ : InMux
    port map (
            O => \N__32018\,
            I => \N__31970\
        );

    \I__4510\ : InMux
    port map (
            O => \N__32017\,
            I => \N__31970\
        );

    \I__4509\ : InMux
    port map (
            O => \N__32016\,
            I => \N__31961\
        );

    \I__4508\ : InMux
    port map (
            O => \N__32015\,
            I => \N__31961\
        );

    \I__4507\ : InMux
    port map (
            O => \N__32014\,
            I => \N__31961\
        );

    \I__4506\ : InMux
    port map (
            O => \N__32013\,
            I => \N__31961\
        );

    \I__4505\ : InMux
    port map (
            O => \N__32012\,
            I => \N__31946\
        );

    \I__4504\ : InMux
    port map (
            O => \N__32009\,
            I => \N__31946\
        );

    \I__4503\ : InMux
    port map (
            O => \N__32008\,
            I => \N__31946\
        );

    \I__4502\ : InMux
    port map (
            O => \N__32005\,
            I => \N__31946\
        );

    \I__4501\ : InMux
    port map (
            O => \N__32004\,
            I => \N__31946\
        );

    \I__4500\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31946\
        );

    \I__4499\ : InMux
    port map (
            O => \N__32000\,
            I => \N__31946\
        );

    \I__4498\ : InMux
    port map (
            O => \N__31999\,
            I => \N__31939\
        );

    \I__4497\ : InMux
    port map (
            O => \N__31998\,
            I => \N__31939\
        );

    \I__4496\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31939\
        );

    \I__4495\ : InMux
    port map (
            O => \N__31996\,
            I => \N__31930\
        );

    \I__4494\ : InMux
    port map (
            O => \N__31995\,
            I => \N__31930\
        );

    \I__4493\ : InMux
    port map (
            O => \N__31994\,
            I => \N__31930\
        );

    \I__4492\ : InMux
    port map (
            O => \N__31993\,
            I => \N__31930\
        );

    \I__4491\ : Odrv4
    port map (
            O => \N__31982\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__31977\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__31970\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__31961\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__31946\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__31939\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__31930\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4484\ : InMux
    port map (
            O => \N__31915\,
            I => \bfn_14_32_0_\
        );

    \I__4483\ : InMux
    port map (
            O => \N__31912\,
            I => \N__31909\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__31909\,
            I => \N__31906\
        );

    \I__4481\ : Span12Mux_h
    port map (
            O => \N__31906\,
            I => \N__31903\
        );

    \I__4480\ : Span12Mux_v
    port map (
            O => \N__31903\,
            I => \N__31900\
        );

    \I__4479\ : Odrv12
    port map (
            O => \N__31900\,
            I => n20764
        );

    \I__4478\ : InMux
    port map (
            O => \N__31897\,
            I => \N__31894\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__31894\,
            I => \N__31891\
        );

    \I__4476\ : Span4Mux_v
    port map (
            O => \N__31891\,
            I => \N__31888\
        );

    \I__4475\ : Odrv4
    port map (
            O => \N__31888\,
            I => n16
        );

    \I__4474\ : SRMux
    port map (
            O => \N__31885\,
            I => \N__31882\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__31882\,
            I => \N__31879\
        );

    \I__4472\ : Span4Mux_h
    port map (
            O => \N__31879\,
            I => \N__31876\
        );

    \I__4471\ : Odrv4
    port map (
            O => \N__31876\,
            I => \c0.n6_adj_3155\
        );

    \I__4470\ : InMux
    port map (
            O => \N__31873\,
            I => \bfn_14_31_0_\
        );

    \I__4469\ : InMux
    port map (
            O => \N__31870\,
            I => \bfn_14_29_0_\
        );

    \I__4468\ : InMux
    port map (
            O => \N__31867\,
            I => \bfn_14_30_0_\
        );

    \I__4467\ : InMux
    port map (
            O => \N__31864\,
            I => \bfn_14_28_0_\
        );

    \I__4466\ : InMux
    port map (
            O => \N__31861\,
            I => \bfn_14_27_0_\
        );

    \I__4465\ : InMux
    port map (
            O => \N__31858\,
            I => \bfn_14_26_0_\
        );

    \I__4464\ : InMux
    port map (
            O => \N__31855\,
            I => \bfn_14_25_0_\
        );

    \I__4463\ : InMux
    port map (
            O => \N__31852\,
            I => \bfn_14_24_0_\
        );

    \I__4462\ : InMux
    port map (
            O => \N__31849\,
            I => \bfn_14_23_0_\
        );

    \I__4461\ : SRMux
    port map (
            O => \N__31846\,
            I => \N__31843\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__31843\,
            I => \N__31840\
        );

    \I__4459\ : Span4Mux_h
    port map (
            O => \N__31840\,
            I => \N__31837\
        );

    \I__4458\ : Odrv4
    port map (
            O => \N__31837\,
            I => \c0.n6_adj_3178\
        );

    \I__4457\ : SRMux
    port map (
            O => \N__31834\,
            I => \N__31831\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__31831\,
            I => \c0.n6_adj_3182\
        );

    \I__4455\ : InMux
    port map (
            O => \N__31828\,
            I => \bfn_14_22_0_\
        );

    \I__4454\ : SRMux
    port map (
            O => \N__31825\,
            I => \N__31822\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__31822\,
            I => \N__31819\
        );

    \I__4452\ : Odrv4
    port map (
            O => \N__31819\,
            I => \c0.n6_adj_3180\
        );

    \I__4451\ : InMux
    port map (
            O => \N__31816\,
            I => \bfn_14_20_0_\
        );

    \I__4450\ : SRMux
    port map (
            O => \N__31813\,
            I => \N__31810\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__31810\,
            I => \N__31807\
        );

    \I__4448\ : Sp12to4
    port map (
            O => \N__31807\,
            I => \N__31804\
        );

    \I__4447\ : Odrv12
    port map (
            O => \N__31804\,
            I => \c0.n6_adj_3184\
        );

    \I__4446\ : InMux
    port map (
            O => \N__31801\,
            I => \bfn_14_21_0_\
        );

    \I__4445\ : InMux
    port map (
            O => \N__31798\,
            I => \bfn_14_19_0_\
        );

    \I__4444\ : SRMux
    port map (
            O => \N__31795\,
            I => \N__31792\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__31792\,
            I => \N__31789\
        );

    \I__4442\ : Odrv4
    port map (
            O => \N__31789\,
            I => \c0.n6_adj_3186\
        );

    \I__4441\ : InMux
    port map (
            O => \N__31786\,
            I => \bfn_14_18_0_\
        );

    \I__4440\ : SRMux
    port map (
            O => \N__31783\,
            I => \N__31780\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__31780\,
            I => \N__31777\
        );

    \I__4438\ : Span4Mux_v
    port map (
            O => \N__31777\,
            I => \N__31774\
        );

    \I__4437\ : Odrv4
    port map (
            O => \N__31774\,
            I => \c0.n6_adj_3188\
        );

    \I__4436\ : InMux
    port map (
            O => \N__31771\,
            I => \bfn_14_17_0_\
        );

    \I__4435\ : InMux
    port map (
            O => \N__31768\,
            I => \bfn_14_16_0_\
        );

    \I__4434\ : InMux
    port map (
            O => \N__31765\,
            I => \bfn_14_15_0_\
        );

    \I__4433\ : InMux
    port map (
            O => \N__31762\,
            I => \bfn_14_14_0_\
        );

    \I__4432\ : SRMux
    port map (
            O => \N__31759\,
            I => \N__31756\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__31756\,
            I => \N__31753\
        );

    \I__4430\ : Span4Mux_v
    port map (
            O => \N__31753\,
            I => \N__31750\
        );

    \I__4429\ : Odrv4
    port map (
            O => \N__31750\,
            I => \c0.n6_adj_3162\
        );

    \I__4428\ : InMux
    port map (
            O => \N__31747\,
            I => \bfn_14_13_0_\
        );

    \I__4427\ : InMux
    port map (
            O => \N__31744\,
            I => \bfn_14_11_0_\
        );

    \I__4426\ : InMux
    port map (
            O => \N__31741\,
            I => \bfn_14_12_0_\
        );

    \I__4425\ : InMux
    port map (
            O => \N__31738\,
            I => \bfn_14_10_0_\
        );

    \I__4424\ : InMux
    port map (
            O => \N__31735\,
            I => \bfn_14_9_0_\
        );

    \I__4423\ : InMux
    port map (
            O => \N__31732\,
            I => \bfn_14_8_0_\
        );

    \I__4422\ : InMux
    port map (
            O => \N__31729\,
            I => \bfn_14_7_0_\
        );

    \I__4421\ : InMux
    port map (
            O => \N__31726\,
            I => \c0.n17177\
        );

    \I__4420\ : InMux
    port map (
            O => \N__31723\,
            I => \N__31720\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__31720\,
            I => \c0.n2_adj_3145\
        );

    \I__4418\ : InMux
    port map (
            O => \N__31717\,
            I => \c0.n17178\
        );

    \I__4417\ : InMux
    port map (
            O => \N__31714\,
            I => \c0.n17179\
        );

    \I__4416\ : InMux
    port map (
            O => \N__31711\,
            I => \bfn_14_6_0_\
        );

    \I__4415\ : InMux
    port map (
            O => \N__31708\,
            I => \N__31705\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__31705\,
            I => \N__31702\
        );

    \I__4413\ : Odrv4
    port map (
            O => \N__31702\,
            I => \c0.n19638\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__31699\,
            I => \c0.n6_adj_3515_cascade_\
        );

    \I__4411\ : InMux
    port map (
            O => \N__31696\,
            I => \N__31693\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__31693\,
            I => \c0.n5_adj_3516\
        );

    \I__4409\ : CascadeMux
    port map (
            O => \N__31690\,
            I => \N__31685\
        );

    \I__4408\ : InMux
    port map (
            O => \N__31689\,
            I => \N__31682\
        );

    \I__4407\ : InMux
    port map (
            O => \N__31688\,
            I => \N__31677\
        );

    \I__4406\ : InMux
    port map (
            O => \N__31685\,
            I => \N__31677\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__31682\,
            I => \c0.FRAME_MATCHER_state_5\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__31677\,
            I => \c0.FRAME_MATCHER_state_5\
        );

    \I__4403\ : SRMux
    port map (
            O => \N__31672\,
            I => \N__31669\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__31669\,
            I => \c0.n18681\
        );

    \I__4401\ : CascadeMux
    port map (
            O => \N__31666\,
            I => \N__31663\
        );

    \I__4400\ : InMux
    port map (
            O => \N__31663\,
            I => \N__31659\
        );

    \I__4399\ : InMux
    port map (
            O => \N__31662\,
            I => \N__31655\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__31659\,
            I => \N__31652\
        );

    \I__4397\ : InMux
    port map (
            O => \N__31658\,
            I => \N__31649\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__31655\,
            I => \N__31646\
        );

    \I__4395\ : Span4Mux_h
    port map (
            O => \N__31652\,
            I => \N__31643\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__31649\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__4393\ : Odrv4
    port map (
            O => \N__31646\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__31643\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__4391\ : SRMux
    port map (
            O => \N__31636\,
            I => \N__31633\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__31633\,
            I => \N__31630\
        );

    \I__4389\ : Odrv4
    port map (
            O => \N__31630\,
            I => \c0.n18657\
        );

    \I__4388\ : InMux
    port map (
            O => \N__31627\,
            I => \N__31622\
        );

    \I__4387\ : InMux
    port map (
            O => \N__31626\,
            I => \N__31619\
        );

    \I__4386\ : InMux
    port map (
            O => \N__31625\,
            I => \N__31616\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__31622\,
            I => \N__31613\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__31619\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__31616\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__4382\ : Odrv4
    port map (
            O => \N__31613\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__4381\ : SRMux
    port map (
            O => \N__31606\,
            I => \N__31603\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__31603\,
            I => \N__31600\
        );

    \I__4379\ : Odrv4
    port map (
            O => \N__31600\,
            I => \c0.n18629\
        );

    \I__4378\ : InMux
    port map (
            O => \N__31597\,
            I => \c0.n17176\
        );

    \I__4377\ : InMux
    port map (
            O => \N__31594\,
            I => \N__31591\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__31591\,
            I => \c0.n2_adj_3144\
        );

    \I__4375\ : CascadeMux
    port map (
            O => \N__31588\,
            I => \c0.n19638_cascade_\
        );

    \I__4374\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31582\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__31582\,
            I => \c0.FRAME_MATCHER_state_31_N_1864_2\
        );

    \I__4372\ : CascadeMux
    port map (
            O => \N__31579\,
            I => \c0.n6_adj_3521_cascade_\
        );

    \I__4371\ : CascadeMux
    port map (
            O => \N__31576\,
            I => \N__31572\
        );

    \I__4370\ : InMux
    port map (
            O => \N__31575\,
            I => \N__31568\
        );

    \I__4369\ : InMux
    port map (
            O => \N__31572\,
            I => \N__31565\
        );

    \I__4368\ : InMux
    port map (
            O => \N__31571\,
            I => \N__31562\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__31568\,
            I => \N__31559\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__31565\,
            I => \N__31556\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__31562\,
            I => \N__31553\
        );

    \I__4364\ : Span4Mux_h
    port map (
            O => \N__31559\,
            I => \N__31550\
        );

    \I__4363\ : Odrv12
    port map (
            O => \N__31556\,
            I => \c0.n936\
        );

    \I__4362\ : Odrv4
    port map (
            O => \N__31553\,
            I => \c0.n936\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__31550\,
            I => \c0.n936\
        );

    \I__4360\ : InMux
    port map (
            O => \N__31543\,
            I => \N__31540\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__31540\,
            I => \c0.n11_adj_3370\
        );

    \I__4358\ : InMux
    port map (
            O => \N__31537\,
            I => \N__31533\
        );

    \I__4357\ : InMux
    port map (
            O => \N__31536\,
            I => \N__31530\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__31533\,
            I => \N__31527\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__31530\,
            I => \N__31524\
        );

    \I__4354\ : Odrv12
    port map (
            O => \N__31527\,
            I => \c0.tx_transmit_N_2443\
        );

    \I__4353\ : Odrv4
    port map (
            O => \N__31524\,
            I => \c0.tx_transmit_N_2443\
        );

    \I__4352\ : InMux
    port map (
            O => \N__31519\,
            I => \N__31516\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__31516\,
            I => \N__31513\
        );

    \I__4350\ : Span4Mux_h
    port map (
            O => \N__31513\,
            I => \N__31510\
        );

    \I__4349\ : Odrv4
    port map (
            O => \N__31510\,
            I => \c0.n21420\
        );

    \I__4348\ : InMux
    port map (
            O => \N__31507\,
            I => \N__31503\
        );

    \I__4347\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31499\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__31503\,
            I => \N__31496\
        );

    \I__4345\ : InMux
    port map (
            O => \N__31502\,
            I => \N__31493\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__31499\,
            I => \N__31488\
        );

    \I__4343\ : Span4Mux_v
    port map (
            O => \N__31496\,
            I => \N__31488\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__31493\,
            I => \N__31485\
        );

    \I__4341\ : Odrv4
    port map (
            O => \N__31488\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__4340\ : Odrv4
    port map (
            O => \N__31485\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__4339\ : SRMux
    port map (
            O => \N__31480\,
            I => \N__31477\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__31477\,
            I => \N__31474\
        );

    \I__4337\ : Span4Mux_h
    port map (
            O => \N__31474\,
            I => \N__31471\
        );

    \I__4336\ : Odrv4
    port map (
            O => \N__31471\,
            I => \c0.n18627\
        );

    \I__4335\ : InMux
    port map (
            O => \N__31468\,
            I => \N__31465\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__31465\,
            I => \N__31462\
        );

    \I__4333\ : Odrv4
    port map (
            O => \N__31462\,
            I => \c0.n19650\
        );

    \I__4332\ : InMux
    port map (
            O => \N__31459\,
            I => \c0.n17349\
        );

    \I__4331\ : InMux
    port map (
            O => \N__31456\,
            I => \c0.n17350\
        );

    \I__4330\ : InMux
    port map (
            O => \N__31453\,
            I => \c0.n17351\
        );

    \I__4329\ : InMux
    port map (
            O => \N__31450\,
            I => \c0.n17352\
        );

    \I__4328\ : SRMux
    port map (
            O => \N__31447\,
            I => \N__31444\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__31444\,
            I => \N__31441\
        );

    \I__4326\ : Span4Mux_v
    port map (
            O => \N__31441\,
            I => \N__31437\
        );

    \I__4325\ : InMux
    port map (
            O => \N__31440\,
            I => \N__31434\
        );

    \I__4324\ : Odrv4
    port map (
            O => \N__31437\,
            I => \c0.n19052\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__31434\,
            I => \c0.n19052\
        );

    \I__4322\ : CascadeMux
    port map (
            O => \N__31429\,
            I => \N__31425\
        );

    \I__4321\ : CascadeMux
    port map (
            O => \N__31428\,
            I => \N__31422\
        );

    \I__4320\ : InMux
    port map (
            O => \N__31425\,
            I => \N__31419\
        );

    \I__4319\ : InMux
    port map (
            O => \N__31422\,
            I => \N__31416\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__31419\,
            I => \N__31413\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__31416\,
            I => \c0.n6_adj_3338\
        );

    \I__4316\ : Odrv4
    port map (
            O => \N__31413\,
            I => \c0.n6_adj_3338\
        );

    \I__4315\ : CEMux
    port map (
            O => \N__31408\,
            I => \N__31405\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__31405\,
            I => \N__31402\
        );

    \I__4313\ : Span4Mux_v
    port map (
            O => \N__31402\,
            I => \N__31399\
        );

    \I__4312\ : Odrv4
    port map (
            O => \N__31399\,
            I => \c0.n12326\
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__31396\,
            I => \c0.n12326_cascade_\
        );

    \I__4310\ : SRMux
    port map (
            O => \N__31393\,
            I => \N__31390\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__31390\,
            I => \N__31387\
        );

    \I__4308\ : Span4Mux_h
    port map (
            O => \N__31387\,
            I => \N__31384\
        );

    \I__4307\ : Odrv4
    port map (
            O => \N__31384\,
            I => \c0.n12758\
        );

    \I__4306\ : CascadeMux
    port map (
            O => \N__31381\,
            I => \c0.n4_adj_3263_cascade_\
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__31378\,
            I => \c0.n936_cascade_\
        );

    \I__4304\ : InMux
    port map (
            O => \N__31375\,
            I => \N__31372\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__31372\,
            I => \c0.n21566\
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__31369\,
            I => \n10_cascade_\
        );

    \I__4301\ : InMux
    port map (
            O => \N__31366\,
            I => \N__31363\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__31363\,
            I => \N__31359\
        );

    \I__4299\ : InMux
    port map (
            O => \N__31362\,
            I => \N__31356\
        );

    \I__4298\ : Odrv4
    port map (
            O => \N__31359\,
            I => \r_Tx_Data_3\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__31356\,
            I => \r_Tx_Data_3\
        );

    \I__4296\ : InMux
    port map (
            O => \N__31351\,
            I => \N__31345\
        );

    \I__4295\ : InMux
    port map (
            O => \N__31350\,
            I => \N__31345\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__31345\,
            I => data_out_frame_12_1
        );

    \I__4293\ : InMux
    port map (
            O => \N__31342\,
            I => \N__31339\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__31339\,
            I => \c0.n11_adj_3104\
        );

    \I__4291\ : InMux
    port map (
            O => \N__31336\,
            I => \N__31333\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__31333\,
            I => \N__31330\
        );

    \I__4289\ : Span4Mux_v
    port map (
            O => \N__31330\,
            I => \N__31327\
        );

    \I__4288\ : Odrv4
    port map (
            O => \N__31327\,
            I => n10_adj_3593
        );

    \I__4287\ : InMux
    port map (
            O => \N__31324\,
            I => \N__31320\
        );

    \I__4286\ : InMux
    port map (
            O => \N__31323\,
            I => \N__31317\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__31320\,
            I => \r_Tx_Data_2\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__31317\,
            I => \r_Tx_Data_2\
        );

    \I__4283\ : InMux
    port map (
            O => \N__31312\,
            I => \c0.n17346\
        );

    \I__4282\ : InMux
    port map (
            O => \N__31309\,
            I => \c0.n17347\
        );

    \I__4281\ : InMux
    port map (
            O => \N__31306\,
            I => \c0.n17348\
        );

    \I__4280\ : CascadeMux
    port map (
            O => \N__31303\,
            I => \N__31299\
        );

    \I__4279\ : CascadeMux
    port map (
            O => \N__31302\,
            I => \N__31296\
        );

    \I__4278\ : InMux
    port map (
            O => \N__31299\,
            I => \N__31290\
        );

    \I__4277\ : InMux
    port map (
            O => \N__31296\,
            I => \N__31290\
        );

    \I__4276\ : CascadeMux
    port map (
            O => \N__31295\,
            I => \N__31287\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__31290\,
            I => \N__31284\
        );

    \I__4274\ : InMux
    port map (
            O => \N__31287\,
            I => \N__31281\
        );

    \I__4273\ : Span4Mux_h
    port map (
            O => \N__31284\,
            I => \N__31278\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__31281\,
            I => tx_active
        );

    \I__4271\ : Odrv4
    port map (
            O => \N__31278\,
            I => tx_active
        );

    \I__4270\ : InMux
    port map (
            O => \N__31273\,
            I => \N__31267\
        );

    \I__4269\ : InMux
    port map (
            O => \N__31272\,
            I => \N__31267\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__31267\,
            I => \c0.n15842\
        );

    \I__4267\ : InMux
    port map (
            O => \N__31264\,
            I => \N__31261\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__31261\,
            I => \N__31258\
        );

    \I__4265\ : Span4Mux_h
    port map (
            O => \N__31258\,
            I => \N__31255\
        );

    \I__4264\ : Odrv4
    port map (
            O => \N__31255\,
            I => \c0.n11_adj_3404\
        );

    \I__4263\ : InMux
    port map (
            O => \N__31252\,
            I => \N__31249\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__31249\,
            I => \c0.n7_adj_3333\
        );

    \I__4261\ : InMux
    port map (
            O => \N__31246\,
            I => \N__31243\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__31243\,
            I => \N__31239\
        );

    \I__4259\ : InMux
    port map (
            O => \N__31242\,
            I => \N__31236\
        );

    \I__4258\ : Span4Mux_v
    port map (
            O => \N__31239\,
            I => \N__31233\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__31236\,
            I => data_out_frame_9_1
        );

    \I__4256\ : Odrv4
    port map (
            O => \N__31233\,
            I => data_out_frame_9_1
        );

    \I__4255\ : InMux
    port map (
            O => \N__31228\,
            I => \N__31225\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__31225\,
            I => \c0.n21605\
        );

    \I__4253\ : CascadeMux
    port map (
            O => \N__31222\,
            I => \N__31219\
        );

    \I__4252\ : InMux
    port map (
            O => \N__31219\,
            I => \N__31215\
        );

    \I__4251\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31212\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__31215\,
            I => \N__31209\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__31212\,
            I => data_out_frame_8_1
        );

    \I__4248\ : Odrv4
    port map (
            O => \N__31209\,
            I => data_out_frame_8_1
        );

    \I__4247\ : CascadeMux
    port map (
            O => \N__31204\,
            I => \c0.n21608_cascade_\
        );

    \I__4246\ : InMux
    port map (
            O => \N__31201\,
            I => \N__31194\
        );

    \I__4245\ : InMux
    port map (
            O => \N__31200\,
            I => \N__31194\
        );

    \I__4244\ : InMux
    port map (
            O => \N__31199\,
            I => \N__31191\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__31194\,
            I => \c0.r_Tx_Data_0\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__31191\,
            I => \c0.r_Tx_Data_0\
        );

    \I__4241\ : InMux
    port map (
            O => \N__31186\,
            I => \N__31183\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__31183\,
            I => \N__31180\
        );

    \I__4239\ : Span4Mux_h
    port map (
            O => \N__31180\,
            I => \N__31177\
        );

    \I__4238\ : Odrv4
    port map (
            O => \N__31177\,
            I => \c0.n21466\
        );

    \I__4237\ : InMux
    port map (
            O => \N__31174\,
            I => \N__31171\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__31171\,
            I => \N__31168\
        );

    \I__4235\ : Span4Mux_v
    port map (
            O => \N__31168\,
            I => \N__31164\
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__31167\,
            I => \N__31160\
        );

    \I__4233\ : Span4Mux_v
    port map (
            O => \N__31164\,
            I => \N__31157\
        );

    \I__4232\ : InMux
    port map (
            O => \N__31163\,
            I => \N__31154\
        );

    \I__4231\ : InMux
    port map (
            O => \N__31160\,
            I => \N__31151\
        );

    \I__4230\ : Odrv4
    port map (
            O => \N__31157\,
            I => encoder1_position_9
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__31154\,
            I => encoder1_position_9
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__31151\,
            I => encoder1_position_9
        );

    \I__4227\ : InMux
    port map (
            O => \N__31144\,
            I => \N__31141\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__31141\,
            I => \N__31137\
        );

    \I__4225\ : CascadeMux
    port map (
            O => \N__31140\,
            I => \N__31134\
        );

    \I__4224\ : Span4Mux_v
    port map (
            O => \N__31137\,
            I => \N__31131\
        );

    \I__4223\ : InMux
    port map (
            O => \N__31134\,
            I => \N__31128\
        );

    \I__4222\ : Span4Mux_v
    port map (
            O => \N__31131\,
            I => \N__31122\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__31128\,
            I => \N__31122\
        );

    \I__4220\ : InMux
    port map (
            O => \N__31127\,
            I => \N__31119\
        );

    \I__4219\ : Span4Mux_h
    port map (
            O => \N__31122\,
            I => \N__31116\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__31119\,
            I => encoder0_position_0
        );

    \I__4217\ : Odrv4
    port map (
            O => \N__31116\,
            I => encoder0_position_0
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__31111\,
            I => \N__31106\
        );

    \I__4215\ : InMux
    port map (
            O => \N__31110\,
            I => \N__31103\
        );

    \I__4214\ : InMux
    port map (
            O => \N__31109\,
            I => \N__31100\
        );

    \I__4213\ : InMux
    port map (
            O => \N__31106\,
            I => \N__31097\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__31103\,
            I => encoder1_position_25
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__31100\,
            I => encoder1_position_25
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__31097\,
            I => encoder1_position_25
        );

    \I__4209\ : CascadeMux
    port map (
            O => \N__31090\,
            I => \N__31087\
        );

    \I__4208\ : InMux
    port map (
            O => \N__31087\,
            I => \N__31083\
        );

    \I__4207\ : InMux
    port map (
            O => \N__31086\,
            I => \N__31080\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__31083\,
            I => \N__31076\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__31080\,
            I => \N__31073\
        );

    \I__4204\ : InMux
    port map (
            O => \N__31079\,
            I => \N__31070\
        );

    \I__4203\ : Span4Mux_h
    port map (
            O => \N__31076\,
            I => \N__31067\
        );

    \I__4202\ : Odrv4
    port map (
            O => \N__31073\,
            I => encoder1_position_2
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__31070\,
            I => encoder1_position_2
        );

    \I__4200\ : Odrv4
    port map (
            O => \N__31067\,
            I => encoder1_position_2
        );

    \I__4199\ : InMux
    port map (
            O => \N__31060\,
            I => \N__31057\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__31057\,
            I => \N__31053\
        );

    \I__4197\ : CascadeMux
    port map (
            O => \N__31056\,
            I => \N__31049\
        );

    \I__4196\ : Span4Mux_v
    port map (
            O => \N__31053\,
            I => \N__31046\
        );

    \I__4195\ : InMux
    port map (
            O => \N__31052\,
            I => \N__31043\
        );

    \I__4194\ : InMux
    port map (
            O => \N__31049\,
            I => \N__31040\
        );

    \I__4193\ : Odrv4
    port map (
            O => \N__31046\,
            I => encoder1_position_17
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__31043\,
            I => encoder1_position_17
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__31040\,
            I => encoder1_position_17
        );

    \I__4190\ : CascadeMux
    port map (
            O => \N__31033\,
            I => \N__31029\
        );

    \I__4189\ : CascadeMux
    port map (
            O => \N__31032\,
            I => \N__31026\
        );

    \I__4188\ : InMux
    port map (
            O => \N__31029\,
            I => \N__31021\
        );

    \I__4187\ : InMux
    port map (
            O => \N__31026\,
            I => \N__31021\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__31021\,
            I => data_out_frame_13_2
        );

    \I__4185\ : InMux
    port map (
            O => \N__31018\,
            I => \N__31014\
        );

    \I__4184\ : InMux
    port map (
            O => \N__31017\,
            I => \N__31011\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__31014\,
            I => data_out_frame_12_2
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__31011\,
            I => data_out_frame_12_2
        );

    \I__4181\ : InMux
    port map (
            O => \N__31006\,
            I => \N__31003\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__31003\,
            I => \N__31000\
        );

    \I__4179\ : Sp12to4
    port map (
            O => \N__31000\,
            I => \N__30997\
        );

    \I__4178\ : Odrv12
    port map (
            O => \N__30997\,
            I => \c0.n11_adj_3108\
        );

    \I__4177\ : InMux
    port map (
            O => \N__30994\,
            I => \N__30990\
        );

    \I__4176\ : InMux
    port map (
            O => \N__30993\,
            I => \N__30987\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__30990\,
            I => data_out_frame_10_1
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__30987\,
            I => data_out_frame_10_1
        );

    \I__4173\ : CascadeMux
    port map (
            O => \N__30982\,
            I => \N__30978\
        );

    \I__4172\ : InMux
    port map (
            O => \N__30981\,
            I => \N__30973\
        );

    \I__4171\ : InMux
    port map (
            O => \N__30978\,
            I => \N__30973\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__30973\,
            I => data_out_frame_11_1
        );

    \I__4169\ : InMux
    port map (
            O => \N__30970\,
            I => \N__30966\
        );

    \I__4168\ : InMux
    port map (
            O => \N__30969\,
            I => \N__30963\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__30966\,
            I => \N__30960\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__30963\,
            I => data_out_frame_13_5
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__30960\,
            I => data_out_frame_13_5
        );

    \I__4164\ : InMux
    port map (
            O => \N__30955\,
            I => \N__30949\
        );

    \I__4163\ : InMux
    port map (
            O => \N__30954\,
            I => \N__30944\
        );

    \I__4162\ : InMux
    port map (
            O => \N__30953\,
            I => \N__30944\
        );

    \I__4161\ : CascadeMux
    port map (
            O => \N__30952\,
            I => \N__30940\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__30949\,
            I => \N__30935\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__30944\,
            I => \N__30935\
        );

    \I__4158\ : InMux
    port map (
            O => \N__30943\,
            I => \N__30932\
        );

    \I__4157\ : InMux
    port map (
            O => \N__30940\,
            I => \N__30929\
        );

    \I__4156\ : Span4Mux_h
    port map (
            O => \N__30935\,
            I => \N__30926\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__30932\,
            I => \c0.r_SM_Main_2_N_2547_0\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__30929\,
            I => \c0.r_SM_Main_2_N_2547_0\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__30926\,
            I => \c0.r_SM_Main_2_N_2547_0\
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__30919\,
            I => \N__30915\
        );

    \I__4151\ : InMux
    port map (
            O => \N__30918\,
            I => \N__30912\
        );

    \I__4150\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30909\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__30912\,
            I => \N__30905\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__30909\,
            I => \N__30902\
        );

    \I__4147\ : InMux
    port map (
            O => \N__30908\,
            I => \N__30899\
        );

    \I__4146\ : Span4Mux_h
    port map (
            O => \N__30905\,
            I => \N__30894\
        );

    \I__4145\ : Span4Mux_h
    port map (
            O => \N__30902\,
            I => \N__30894\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__30899\,
            I => encoder1_position_4
        );

    \I__4143\ : Odrv4
    port map (
            O => \N__30894\,
            I => encoder1_position_4
        );

    \I__4142\ : InMux
    port map (
            O => \N__30889\,
            I => \N__30886\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__30886\,
            I => \N__30882\
        );

    \I__4140\ : InMux
    port map (
            O => \N__30885\,
            I => \N__30879\
        );

    \I__4139\ : Span4Mux_h
    port map (
            O => \N__30882\,
            I => \N__30876\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__30879\,
            I => data_out_frame_13_4
        );

    \I__4137\ : Odrv4
    port map (
            O => \N__30876\,
            I => data_out_frame_13_4
        );

    \I__4136\ : InMux
    port map (
            O => \N__30871\,
            I => \N__30862\
        );

    \I__4135\ : InMux
    port map (
            O => \N__30870\,
            I => \N__30862\
        );

    \I__4134\ : InMux
    port map (
            O => \N__30869\,
            I => \N__30862\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__30862\,
            I => encoder1_position_31
        );

    \I__4132\ : InMux
    port map (
            O => \N__30859\,
            I => \N__30856\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__30856\,
            I => n2320
        );

    \I__4130\ : InMux
    port map (
            O => \N__30853\,
            I => \N__30849\
        );

    \I__4129\ : CascadeMux
    port map (
            O => \N__30852\,
            I => \N__30846\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__30849\,
            I => \N__30843\
        );

    \I__4127\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30840\
        );

    \I__4126\ : Span4Mux_v
    port map (
            O => \N__30843\,
            I => \N__30837\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__30840\,
            I => \r_Tx_Data_5\
        );

    \I__4124\ : Odrv4
    port map (
            O => \N__30837\,
            I => \r_Tx_Data_5\
        );

    \I__4123\ : InMux
    port map (
            O => \N__30832\,
            I => \N__30829\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__30829\,
            I => \N__30825\
        );

    \I__4121\ : InMux
    port map (
            O => \N__30828\,
            I => \N__30822\
        );

    \I__4120\ : Span4Mux_h
    port map (
            O => \N__30825\,
            I => \N__30819\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__30822\,
            I => data_out_frame_9_4
        );

    \I__4118\ : Odrv4
    port map (
            O => \N__30819\,
            I => data_out_frame_9_4
        );

    \I__4117\ : InMux
    port map (
            O => \N__30814\,
            I => \N__30810\
        );

    \I__4116\ : InMux
    port map (
            O => \N__30813\,
            I => \N__30807\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__30810\,
            I => data_out_frame_8_4
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__30807\,
            I => data_out_frame_8_4
        );

    \I__4113\ : InMux
    port map (
            O => \N__30802\,
            I => \N__30799\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__30799\,
            I => \N__30796\
        );

    \I__4111\ : Span4Mux_v
    port map (
            O => \N__30796\,
            I => \N__30793\
        );

    \I__4110\ : Odrv4
    port map (
            O => \N__30793\,
            I => \c0.n21287\
        );

    \I__4109\ : CascadeMux
    port map (
            O => \N__30790\,
            I => \N__30787\
        );

    \I__4108\ : InMux
    port map (
            O => \N__30787\,
            I => \N__30783\
        );

    \I__4107\ : InMux
    port map (
            O => \N__30786\,
            I => \N__30779\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__30783\,
            I => \N__30776\
        );

    \I__4105\ : InMux
    port map (
            O => \N__30782\,
            I => \N__30773\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__30779\,
            I => \N__30768\
        );

    \I__4103\ : Span4Mux_h
    port map (
            O => \N__30776\,
            I => \N__30768\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__30773\,
            I => encoder0_position_9
        );

    \I__4101\ : Odrv4
    port map (
            O => \N__30768\,
            I => encoder0_position_9
        );

    \I__4100\ : InMux
    port map (
            O => \N__30763\,
            I => \N__30759\
        );

    \I__4099\ : CascadeMux
    port map (
            O => \N__30762\,
            I => \N__30756\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__30759\,
            I => \N__30753\
        );

    \I__4097\ : InMux
    port map (
            O => \N__30756\,
            I => \N__30749\
        );

    \I__4096\ : Span4Mux_v
    port map (
            O => \N__30753\,
            I => \N__30746\
        );

    \I__4095\ : InMux
    port map (
            O => \N__30752\,
            I => \N__30743\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__30749\,
            I => encoder1_position_24
        );

    \I__4093\ : Odrv4
    port map (
            O => \N__30746\,
            I => encoder1_position_24
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__30743\,
            I => encoder1_position_24
        );

    \I__4091\ : CascadeMux
    port map (
            O => \N__30736\,
            I => \N__30732\
        );

    \I__4090\ : InMux
    port map (
            O => \N__30735\,
            I => \N__30729\
        );

    \I__4089\ : InMux
    port map (
            O => \N__30732\,
            I => \N__30726\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__30729\,
            I => \c0.data_out_frame_0_4\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__30726\,
            I => \c0.data_out_frame_0_4\
        );

    \I__4086\ : CascadeMux
    port map (
            O => \N__30721\,
            I => \N__30718\
        );

    \I__4085\ : InMux
    port map (
            O => \N__30718\,
            I => \N__30715\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__30715\,
            I => \N__30710\
        );

    \I__4083\ : InMux
    port map (
            O => \N__30714\,
            I => \N__30707\
        );

    \I__4082\ : InMux
    port map (
            O => \N__30713\,
            I => \N__30704\
        );

    \I__4081\ : Span4Mux_h
    port map (
            O => \N__30710\,
            I => \N__30701\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__30707\,
            I => encoder0_position_8
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__30704\,
            I => encoder0_position_8
        );

    \I__4078\ : Odrv4
    port map (
            O => \N__30701\,
            I => encoder0_position_8
        );

    \I__4077\ : InMux
    port map (
            O => \N__30694\,
            I => \N__30691\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__30691\,
            I => n2319
        );

    \I__4075\ : InMux
    port map (
            O => \N__30688\,
            I => \quad_counter1.n17340\
        );

    \I__4074\ : InMux
    port map (
            O => \N__30685\,
            I => \N__30681\
        );

    \I__4073\ : CascadeMux
    port map (
            O => \N__30684\,
            I => \N__30677\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__30681\,
            I => \N__30674\
        );

    \I__4071\ : InMux
    port map (
            O => \N__30680\,
            I => \N__30671\
        );

    \I__4070\ : InMux
    port map (
            O => \N__30677\,
            I => \N__30668\
        );

    \I__4069\ : Odrv12
    port map (
            O => \N__30674\,
            I => encoder1_position_27
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__30671\,
            I => encoder1_position_27
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__30668\,
            I => encoder1_position_27
        );

    \I__4066\ : InMux
    port map (
            O => \N__30661\,
            I => \N__30658\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__30658\,
            I => n2318
        );

    \I__4064\ : InMux
    port map (
            O => \N__30655\,
            I => \quad_counter1.n17341\
        );

    \I__4063\ : InMux
    port map (
            O => \N__30652\,
            I => \quad_counter1.n17342\
        );

    \I__4062\ : InMux
    port map (
            O => \N__30649\,
            I => \quad_counter1.n17343\
        );

    \I__4061\ : InMux
    port map (
            O => \N__30646\,
            I => \N__30643\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__30643\,
            I => \N__30639\
        );

    \I__4059\ : InMux
    port map (
            O => \N__30642\,
            I => \N__30635\
        );

    \I__4058\ : Span4Mux_v
    port map (
            O => \N__30639\,
            I => \N__30632\
        );

    \I__4057\ : InMux
    port map (
            O => \N__30638\,
            I => \N__30629\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__30635\,
            I => \N__30626\
        );

    \I__4055\ : Span4Mux_v
    port map (
            O => \N__30632\,
            I => \N__30619\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__30629\,
            I => \N__30619\
        );

    \I__4053\ : Span4Mux_v
    port map (
            O => \N__30626\,
            I => \N__30619\
        );

    \I__4052\ : Odrv4
    port map (
            O => \N__30619\,
            I => encoder1_position_30
        );

    \I__4051\ : InMux
    port map (
            O => \N__30616\,
            I => \N__30613\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__30613\,
            I => \N__30610\
        );

    \I__4049\ : Span4Mux_h
    port map (
            O => \N__30610\,
            I => \N__30607\
        );

    \I__4048\ : Odrv4
    port map (
            O => \N__30607\,
            I => n2315
        );

    \I__4047\ : InMux
    port map (
            O => \N__30604\,
            I => \quad_counter1.n17344\
        );

    \I__4046\ : CascadeMux
    port map (
            O => \N__30601\,
            I => \N__30594\
        );

    \I__4045\ : CascadeMux
    port map (
            O => \N__30600\,
            I => \N__30590\
        );

    \I__4044\ : CascadeMux
    port map (
            O => \N__30599\,
            I => \N__30586\
        );

    \I__4043\ : CascadeMux
    port map (
            O => \N__30598\,
            I => \N__30582\
        );

    \I__4042\ : InMux
    port map (
            O => \N__30597\,
            I => \N__30561\
        );

    \I__4041\ : InMux
    port map (
            O => \N__30594\,
            I => \N__30544\
        );

    \I__4040\ : InMux
    port map (
            O => \N__30593\,
            I => \N__30544\
        );

    \I__4039\ : InMux
    port map (
            O => \N__30590\,
            I => \N__30544\
        );

    \I__4038\ : InMux
    port map (
            O => \N__30589\,
            I => \N__30544\
        );

    \I__4037\ : InMux
    port map (
            O => \N__30586\,
            I => \N__30544\
        );

    \I__4036\ : InMux
    port map (
            O => \N__30585\,
            I => \N__30544\
        );

    \I__4035\ : InMux
    port map (
            O => \N__30582\,
            I => \N__30544\
        );

    \I__4034\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30544\
        );

    \I__4033\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30535\
        );

    \I__4032\ : InMux
    port map (
            O => \N__30579\,
            I => \N__30535\
        );

    \I__4031\ : InMux
    port map (
            O => \N__30578\,
            I => \N__30535\
        );

    \I__4030\ : InMux
    port map (
            O => \N__30577\,
            I => \N__30535\
        );

    \I__4029\ : InMux
    port map (
            O => \N__30576\,
            I => \N__30526\
        );

    \I__4028\ : InMux
    port map (
            O => \N__30575\,
            I => \N__30526\
        );

    \I__4027\ : InMux
    port map (
            O => \N__30574\,
            I => \N__30526\
        );

    \I__4026\ : InMux
    port map (
            O => \N__30573\,
            I => \N__30526\
        );

    \I__4025\ : InMux
    port map (
            O => \N__30572\,
            I => \N__30517\
        );

    \I__4024\ : InMux
    port map (
            O => \N__30571\,
            I => \N__30517\
        );

    \I__4023\ : InMux
    port map (
            O => \N__30570\,
            I => \N__30517\
        );

    \I__4022\ : InMux
    port map (
            O => \N__30569\,
            I => \N__30517\
        );

    \I__4021\ : InMux
    port map (
            O => \N__30568\,
            I => \N__30508\
        );

    \I__4020\ : InMux
    port map (
            O => \N__30567\,
            I => \N__30508\
        );

    \I__4019\ : InMux
    port map (
            O => \N__30566\,
            I => \N__30508\
        );

    \I__4018\ : InMux
    port map (
            O => \N__30565\,
            I => \N__30508\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__30564\,
            I => \N__30502\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__30561\,
            I => \N__30493\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__30544\,
            I => \N__30493\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__30535\,
            I => \N__30484\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__30526\,
            I => \N__30484\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__30517\,
            I => \N__30484\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__30508\,
            I => \N__30484\
        );

    \I__4010\ : InMux
    port map (
            O => \N__30507\,
            I => \N__30475\
        );

    \I__4009\ : InMux
    port map (
            O => \N__30506\,
            I => \N__30475\
        );

    \I__4008\ : InMux
    port map (
            O => \N__30505\,
            I => \N__30475\
        );

    \I__4007\ : InMux
    port map (
            O => \N__30502\,
            I => \N__30475\
        );

    \I__4006\ : InMux
    port map (
            O => \N__30501\,
            I => \N__30466\
        );

    \I__4005\ : InMux
    port map (
            O => \N__30500\,
            I => \N__30466\
        );

    \I__4004\ : InMux
    port map (
            O => \N__30499\,
            I => \N__30466\
        );

    \I__4003\ : InMux
    port map (
            O => \N__30498\,
            I => \N__30466\
        );

    \I__4002\ : Odrv12
    port map (
            O => \N__30493\,
            I => \quad_counter1.n2301\
        );

    \I__4001\ : Odrv4
    port map (
            O => \N__30484\,
            I => \quad_counter1.n2301\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__30475\,
            I => \quad_counter1.n2301\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__30466\,
            I => \quad_counter1.n2301\
        );

    \I__3998\ : InMux
    port map (
            O => \N__30457\,
            I => \bfn_13_13_0_\
        );

    \I__3997\ : InMux
    port map (
            O => \N__30454\,
            I => \N__30451\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__30451\,
            I => n2314
        );

    \I__3995\ : InMux
    port map (
            O => \N__30448\,
            I => \N__30445\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__30445\,
            I => \N__30442\
        );

    \I__3993\ : Odrv12
    port map (
            O => \N__30442\,
            I => n2345
        );

    \I__3992\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30435\
        );

    \I__3991\ : InMux
    port map (
            O => \N__30438\,
            I => \N__30432\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__30435\,
            I => data_out_frame_12_5
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__30432\,
            I => data_out_frame_12_5
        );

    \I__3988\ : InMux
    port map (
            O => \N__30427\,
            I => \N__30424\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__30424\,
            I => \N__30421\
        );

    \I__3986\ : Odrv4
    port map (
            O => \N__30421\,
            I => n2327
        );

    \I__3985\ : InMux
    port map (
            O => \N__30418\,
            I => \quad_counter1.n17332\
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__30415\,
            I => \N__30412\
        );

    \I__3983\ : InMux
    port map (
            O => \N__30412\,
            I => \N__30408\
        );

    \I__3982\ : InMux
    port map (
            O => \N__30411\,
            I => \N__30404\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__30408\,
            I => \N__30401\
        );

    \I__3980\ : InMux
    port map (
            O => \N__30407\,
            I => \N__30398\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__30404\,
            I => \N__30393\
        );

    \I__3978\ : Span4Mux_h
    port map (
            O => \N__30401\,
            I => \N__30393\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__30398\,
            I => encoder1_position_19
        );

    \I__3976\ : Odrv4
    port map (
            O => \N__30393\,
            I => encoder1_position_19
        );

    \I__3975\ : InMux
    port map (
            O => \N__30388\,
            I => \N__30385\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__30385\,
            I => \N__30382\
        );

    \I__3973\ : Span4Mux_v
    port map (
            O => \N__30382\,
            I => \N__30379\
        );

    \I__3972\ : Odrv4
    port map (
            O => \N__30379\,
            I => n2326
        );

    \I__3971\ : InMux
    port map (
            O => \N__30376\,
            I => \quad_counter1.n17333\
        );

    \I__3970\ : InMux
    port map (
            O => \N__30373\,
            I => \N__30369\
        );

    \I__3969\ : CascadeMux
    port map (
            O => \N__30372\,
            I => \N__30365\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__30369\,
            I => \N__30362\
        );

    \I__3967\ : InMux
    port map (
            O => \N__30368\,
            I => \N__30359\
        );

    \I__3966\ : InMux
    port map (
            O => \N__30365\,
            I => \N__30356\
        );

    \I__3965\ : Odrv4
    port map (
            O => \N__30362\,
            I => encoder1_position_20
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__30359\,
            I => encoder1_position_20
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__30356\,
            I => encoder1_position_20
        );

    \I__3962\ : InMux
    port map (
            O => \N__30349\,
            I => \N__30346\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__30346\,
            I => n2325
        );

    \I__3960\ : InMux
    port map (
            O => \N__30343\,
            I => \quad_counter1.n17334\
        );

    \I__3959\ : InMux
    port map (
            O => \N__30340\,
            I => \quad_counter1.n17335\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__30337\,
            I => \N__30332\
        );

    \I__3957\ : InMux
    port map (
            O => \N__30336\,
            I => \N__30329\
        );

    \I__3956\ : InMux
    port map (
            O => \N__30335\,
            I => \N__30326\
        );

    \I__3955\ : InMux
    port map (
            O => \N__30332\,
            I => \N__30323\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__30329\,
            I => encoder1_position_22
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__30326\,
            I => encoder1_position_22
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__30323\,
            I => encoder1_position_22
        );

    \I__3951\ : InMux
    port map (
            O => \N__30316\,
            I => \N__30313\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__30313\,
            I => n2323
        );

    \I__3949\ : InMux
    port map (
            O => \N__30310\,
            I => \quad_counter1.n17336\
        );

    \I__3948\ : InMux
    port map (
            O => \N__30307\,
            I => \bfn_13_12_0_\
        );

    \I__3947\ : InMux
    port map (
            O => \N__30304\,
            I => \N__30301\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__30301\,
            I => n2321
        );

    \I__3945\ : InMux
    port map (
            O => \N__30298\,
            I => \quad_counter1.n17338\
        );

    \I__3944\ : InMux
    port map (
            O => \N__30295\,
            I => \quad_counter1.n17339\
        );

    \I__3943\ : InMux
    port map (
            O => \N__30292\,
            I => \N__30288\
        );

    \I__3942\ : CascadeMux
    port map (
            O => \N__30291\,
            I => \N__30284\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__30288\,
            I => \N__30281\
        );

    \I__3940\ : InMux
    port map (
            O => \N__30287\,
            I => \N__30278\
        );

    \I__3939\ : InMux
    port map (
            O => \N__30284\,
            I => \N__30275\
        );

    \I__3938\ : Odrv12
    port map (
            O => \N__30281\,
            I => encoder1_position_10
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__30278\,
            I => encoder1_position_10
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__30275\,
            I => encoder1_position_10
        );

    \I__3935\ : InMux
    port map (
            O => \N__30268\,
            I => \N__30265\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__30265\,
            I => n2335
        );

    \I__3933\ : InMux
    port map (
            O => \N__30262\,
            I => \quad_counter1.n17324\
        );

    \I__3932\ : InMux
    port map (
            O => \N__30259\,
            I => \N__30256\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__30256\,
            I => \N__30252\
        );

    \I__3930\ : CascadeMux
    port map (
            O => \N__30255\,
            I => \N__30248\
        );

    \I__3929\ : Span4Mux_v
    port map (
            O => \N__30252\,
            I => \N__30245\
        );

    \I__3928\ : InMux
    port map (
            O => \N__30251\,
            I => \N__30242\
        );

    \I__3927\ : InMux
    port map (
            O => \N__30248\,
            I => \N__30239\
        );

    \I__3926\ : Odrv4
    port map (
            O => \N__30245\,
            I => encoder1_position_11
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__30242\,
            I => encoder1_position_11
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__30239\,
            I => encoder1_position_11
        );

    \I__3923\ : InMux
    port map (
            O => \N__30232\,
            I => \N__30229\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__30229\,
            I => n2334
        );

    \I__3921\ : InMux
    port map (
            O => \N__30226\,
            I => \quad_counter1.n17325\
        );

    \I__3920\ : InMux
    port map (
            O => \N__30223\,
            I => \quad_counter1.n17326\
        );

    \I__3919\ : InMux
    port map (
            O => \N__30220\,
            I => \N__30215\
        );

    \I__3918\ : CascadeMux
    port map (
            O => \N__30219\,
            I => \N__30212\
        );

    \I__3917\ : InMux
    port map (
            O => \N__30218\,
            I => \N__30209\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__30215\,
            I => \N__30206\
        );

    \I__3915\ : InMux
    port map (
            O => \N__30212\,
            I => \N__30203\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__30209\,
            I => encoder1_position_13
        );

    \I__3913\ : Odrv4
    port map (
            O => \N__30206\,
            I => encoder1_position_13
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__30203\,
            I => encoder1_position_13
        );

    \I__3911\ : InMux
    port map (
            O => \N__30196\,
            I => \N__30193\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__30193\,
            I => n2332
        );

    \I__3909\ : InMux
    port map (
            O => \N__30190\,
            I => \quad_counter1.n17327\
        );

    \I__3908\ : InMux
    port map (
            O => \N__30187\,
            I => \N__30182\
        );

    \I__3907\ : CascadeMux
    port map (
            O => \N__30186\,
            I => \N__30179\
        );

    \I__3906\ : InMux
    port map (
            O => \N__30185\,
            I => \N__30176\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__30182\,
            I => \N__30173\
        );

    \I__3904\ : InMux
    port map (
            O => \N__30179\,
            I => \N__30170\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__30176\,
            I => encoder1_position_14
        );

    \I__3902\ : Odrv4
    port map (
            O => \N__30173\,
            I => encoder1_position_14
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__30170\,
            I => encoder1_position_14
        );

    \I__3900\ : InMux
    port map (
            O => \N__30163\,
            I => \N__30160\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__30160\,
            I => n2331
        );

    \I__3898\ : InMux
    port map (
            O => \N__30157\,
            I => \quad_counter1.n17328\
        );

    \I__3897\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30150\
        );

    \I__3896\ : CascadeMux
    port map (
            O => \N__30153\,
            I => \N__30146\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__30150\,
            I => \N__30143\
        );

    \I__3894\ : InMux
    port map (
            O => \N__30149\,
            I => \N__30140\
        );

    \I__3893\ : InMux
    port map (
            O => \N__30146\,
            I => \N__30137\
        );

    \I__3892\ : Odrv12
    port map (
            O => \N__30143\,
            I => encoder1_position_15
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__30140\,
            I => encoder1_position_15
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__30137\,
            I => encoder1_position_15
        );

    \I__3889\ : InMux
    port map (
            O => \N__30130\,
            I => \N__30127\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__30127\,
            I => n2330
        );

    \I__3887\ : InMux
    port map (
            O => \N__30124\,
            I => \bfn_13_11_0_\
        );

    \I__3886\ : InMux
    port map (
            O => \N__30121\,
            I => \N__30118\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__30118\,
            I => \N__30113\
        );

    \I__3884\ : CascadeMux
    port map (
            O => \N__30117\,
            I => \N__30110\
        );

    \I__3883\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30107\
        );

    \I__3882\ : Span4Mux_h
    port map (
            O => \N__30113\,
            I => \N__30104\
        );

    \I__3881\ : InMux
    port map (
            O => \N__30110\,
            I => \N__30101\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__30107\,
            I => encoder1_position_16
        );

    \I__3879\ : Odrv4
    port map (
            O => \N__30104\,
            I => encoder1_position_16
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__30101\,
            I => encoder1_position_16
        );

    \I__3877\ : InMux
    port map (
            O => \N__30094\,
            I => \N__30091\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__30091\,
            I => n2329
        );

    \I__3875\ : InMux
    port map (
            O => \N__30088\,
            I => \quad_counter1.n17330\
        );

    \I__3874\ : InMux
    port map (
            O => \N__30085\,
            I => \N__30082\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__30082\,
            I => n2328
        );

    \I__3872\ : InMux
    port map (
            O => \N__30079\,
            I => \quad_counter1.n17331\
        );

    \I__3871\ : InMux
    port map (
            O => \N__30076\,
            I => \quad_counter1.n17315\
        );

    \I__3870\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30070\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__30070\,
            I => \N__30067\
        );

    \I__3868\ : Span4Mux_v
    port map (
            O => \N__30067\,
            I => \N__30064\
        );

    \I__3867\ : Odrv4
    port map (
            O => \N__30064\,
            I => n2343
        );

    \I__3866\ : InMux
    port map (
            O => \N__30061\,
            I => \quad_counter1.n17316\
        );

    \I__3865\ : InMux
    port map (
            O => \N__30058\,
            I => \quad_counter1.n17317\
        );

    \I__3864\ : InMux
    port map (
            O => \N__30055\,
            I => \N__30052\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__30052\,
            I => \N__30049\
        );

    \I__3862\ : Span4Mux_h
    port map (
            O => \N__30049\,
            I => \N__30046\
        );

    \I__3861\ : Odrv4
    port map (
            O => \N__30046\,
            I => n2341
        );

    \I__3860\ : InMux
    port map (
            O => \N__30043\,
            I => \quad_counter1.n17318\
        );

    \I__3859\ : InMux
    port map (
            O => \N__30040\,
            I => \quad_counter1.n17319\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__30037\,
            I => \N__30034\
        );

    \I__3857\ : InMux
    port map (
            O => \N__30034\,
            I => \N__30030\
        );

    \I__3856\ : InMux
    port map (
            O => \N__30033\,
            I => \N__30026\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__30030\,
            I => \N__30023\
        );

    \I__3854\ : InMux
    port map (
            O => \N__30029\,
            I => \N__30020\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__30026\,
            I => \N__30017\
        );

    \I__3852\ : Span4Mux_h
    port map (
            O => \N__30023\,
            I => \N__30014\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__30020\,
            I => encoder1_position_6
        );

    \I__3850\ : Odrv12
    port map (
            O => \N__30017\,
            I => encoder1_position_6
        );

    \I__3849\ : Odrv4
    port map (
            O => \N__30014\,
            I => encoder1_position_6
        );

    \I__3848\ : InMux
    port map (
            O => \N__30007\,
            I => \N__30004\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__30004\,
            I => \N__30001\
        );

    \I__3846\ : Span4Mux_v
    port map (
            O => \N__30001\,
            I => \N__29998\
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__29998\,
            I => n2339
        );

    \I__3844\ : InMux
    port map (
            O => \N__29995\,
            I => \quad_counter1.n17320\
        );

    \I__3843\ : CascadeMux
    port map (
            O => \N__29992\,
            I => \N__29988\
        );

    \I__3842\ : InMux
    port map (
            O => \N__29991\,
            I => \N__29985\
        );

    \I__3841\ : InMux
    port map (
            O => \N__29988\,
            I => \N__29982\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__29985\,
            I => \N__29979\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__29982\,
            I => \N__29975\
        );

    \I__3838\ : Span4Mux_v
    port map (
            O => \N__29979\,
            I => \N__29972\
        );

    \I__3837\ : InMux
    port map (
            O => \N__29978\,
            I => \N__29969\
        );

    \I__3836\ : Span4Mux_h
    port map (
            O => \N__29975\,
            I => \N__29966\
        );

    \I__3835\ : Odrv4
    port map (
            O => \N__29972\,
            I => encoder1_position_7
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__29969\,
            I => encoder1_position_7
        );

    \I__3833\ : Odrv4
    port map (
            O => \N__29966\,
            I => encoder1_position_7
        );

    \I__3832\ : InMux
    port map (
            O => \N__29959\,
            I => \N__29956\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__29956\,
            I => \N__29953\
        );

    \I__3830\ : Span4Mux_h
    port map (
            O => \N__29953\,
            I => \N__29950\
        );

    \I__3829\ : Odrv4
    port map (
            O => \N__29950\,
            I => n2338
        );

    \I__3828\ : InMux
    port map (
            O => \N__29947\,
            I => \bfn_13_10_0_\
        );

    \I__3827\ : InMux
    port map (
            O => \N__29944\,
            I => \N__29941\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__29941\,
            I => \N__29938\
        );

    \I__3825\ : Span4Mux_h
    port map (
            O => \N__29938\,
            I => \N__29935\
        );

    \I__3824\ : Odrv4
    port map (
            O => \N__29935\,
            I => n2337
        );

    \I__3823\ : InMux
    port map (
            O => \N__29932\,
            I => \quad_counter1.n17322\
        );

    \I__3822\ : InMux
    port map (
            O => \N__29929\,
            I => \N__29926\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__29926\,
            I => n2336
        );

    \I__3820\ : InMux
    port map (
            O => \N__29923\,
            I => \quad_counter1.n17323\
        );

    \I__3819\ : InMux
    port map (
            O => \N__29920\,
            I => \N__29917\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__29917\,
            I => \quad_counter1.A_delayed\
        );

    \I__3817\ : InMux
    port map (
            O => \N__29914\,
            I => \N__29910\
        );

    \I__3816\ : InMux
    port map (
            O => \N__29913\,
            I => \N__29907\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__29910\,
            I => \N__29904\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__29907\,
            I => \N__29900\
        );

    \I__3813\ : Span4Mux_h
    port map (
            O => \N__29904\,
            I => \N__29897\
        );

    \I__3812\ : InMux
    port map (
            O => \N__29903\,
            I => \N__29894\
        );

    \I__3811\ : Span4Mux_h
    port map (
            O => \N__29900\,
            I => \N__29891\
        );

    \I__3810\ : Odrv4
    port map (
            O => \N__29897\,
            I => \B_filtered_adj_3582\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__29894\,
            I => \B_filtered_adj_3582\
        );

    \I__3808\ : Odrv4
    port map (
            O => \N__29891\,
            I => \B_filtered_adj_3582\
        );

    \I__3807\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29879\
        );

    \I__3806\ : InMux
    port map (
            O => \N__29883\,
            I => \N__29874\
        );

    \I__3805\ : InMux
    port map (
            O => \N__29882\,
            I => \N__29874\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__29879\,
            I => \quad_counter1.B_delayed\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__29874\,
            I => \quad_counter1.B_delayed\
        );

    \I__3802\ : CascadeMux
    port map (
            O => \N__29869\,
            I => \N__29863\
        );

    \I__3801\ : InMux
    port map (
            O => \N__29868\,
            I => \N__29858\
        );

    \I__3800\ : InMux
    port map (
            O => \N__29867\,
            I => \N__29858\
        );

    \I__3799\ : InMux
    port map (
            O => \N__29866\,
            I => \N__29852\
        );

    \I__3798\ : InMux
    port map (
            O => \N__29863\,
            I => \N__29852\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__29858\,
            I => \N__29849\
        );

    \I__3796\ : InMux
    port map (
            O => \N__29857\,
            I => \N__29846\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__29852\,
            I => \N__29843\
        );

    \I__3794\ : Span4Mux_h
    port map (
            O => \N__29849\,
            I => \N__29840\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__29846\,
            I => \A_filtered_adj_3581\
        );

    \I__3792\ : Odrv4
    port map (
            O => \N__29843\,
            I => \A_filtered_adj_3581\
        );

    \I__3791\ : Odrv4
    port map (
            O => \N__29840\,
            I => \A_filtered_adj_3581\
        );

    \I__3790\ : InMux
    port map (
            O => \N__29833\,
            I => \N__29830\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__29830\,
            I => \quad_counter1.count_direction\
        );

    \I__3788\ : InMux
    port map (
            O => \N__29827\,
            I => \quad_counter1.n17314\
        );

    \I__3787\ : InMux
    port map (
            O => \N__29824\,
            I => \N__29821\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__29821\,
            I => \N__29818\
        );

    \I__3785\ : Span4Mux_v
    port map (
            O => \N__29818\,
            I => \N__29813\
        );

    \I__3784\ : InMux
    port map (
            O => \N__29817\,
            I => \N__29810\
        );

    \I__3783\ : InMux
    port map (
            O => \N__29816\,
            I => \N__29807\
        );

    \I__3782\ : Span4Mux_h
    port map (
            O => \N__29813\,
            I => \N__29804\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__29810\,
            I => \c0.FRAME_MATCHER_state_27\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__29807\,
            I => \c0.FRAME_MATCHER_state_27\
        );

    \I__3779\ : Odrv4
    port map (
            O => \N__29804\,
            I => \c0.FRAME_MATCHER_state_27\
        );

    \I__3778\ : InMux
    port map (
            O => \N__29797\,
            I => \N__29793\
        );

    \I__3777\ : InMux
    port map (
            O => \N__29796\,
            I => \N__29789\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__29793\,
            I => \N__29786\
        );

    \I__3775\ : InMux
    port map (
            O => \N__29792\,
            I => \N__29783\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__29789\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__3773\ : Odrv4
    port map (
            O => \N__29786\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__29783\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__3771\ : InMux
    port map (
            O => \N__29776\,
            I => \N__29772\
        );

    \I__3770\ : InMux
    port map (
            O => \N__29775\,
            I => \N__29768\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__29772\,
            I => \N__29765\
        );

    \I__3768\ : InMux
    port map (
            O => \N__29771\,
            I => \N__29762\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__29768\,
            I => \N__29759\
        );

    \I__3766\ : Span4Mux_h
    port map (
            O => \N__29765\,
            I => \N__29756\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__29762\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__3764\ : Odrv4
    port map (
            O => \N__29759\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__3763\ : Odrv4
    port map (
            O => \N__29756\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__3762\ : CascadeMux
    port map (
            O => \N__29749\,
            I => \N__29746\
        );

    \I__3761\ : InMux
    port map (
            O => \N__29746\,
            I => \N__29743\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__29743\,
            I => \N__29740\
        );

    \I__3759\ : Odrv4
    port map (
            O => \N__29740\,
            I => \c0.n17_adj_3486\
        );

    \I__3758\ : InMux
    port map (
            O => \N__29737\,
            I => \N__29730\
        );

    \I__3757\ : InMux
    port map (
            O => \N__29736\,
            I => \N__29730\
        );

    \I__3756\ : InMux
    port map (
            O => \N__29735\,
            I => \N__29726\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__29730\,
            I => \N__29723\
        );

    \I__3754\ : InMux
    port map (
            O => \N__29729\,
            I => \N__29720\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__29726\,
            I => \N__29717\
        );

    \I__3752\ : Span4Mux_v
    port map (
            O => \N__29723\,
            I => \N__29714\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__29720\,
            I => \c0.FRAME_MATCHER_state_7\
        );

    \I__3750\ : Odrv4
    port map (
            O => \N__29717\,
            I => \c0.FRAME_MATCHER_state_7\
        );

    \I__3749\ : Odrv4
    port map (
            O => \N__29714\,
            I => \c0.FRAME_MATCHER_state_7\
        );

    \I__3748\ : SRMux
    port map (
            O => \N__29707\,
            I => \N__29704\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__29704\,
            I => \N__29701\
        );

    \I__3746\ : Span4Mux_h
    port map (
            O => \N__29701\,
            I => \N__29698\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__29698\,
            I => \c0.n18677\
        );

    \I__3744\ : CascadeMux
    port map (
            O => \N__29695\,
            I => \N__29691\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__29694\,
            I => \N__29688\
        );

    \I__3742\ : InMux
    port map (
            O => \N__29691\,
            I => \N__29684\
        );

    \I__3741\ : InMux
    port map (
            O => \N__29688\,
            I => \N__29681\
        );

    \I__3740\ : InMux
    port map (
            O => \N__29687\,
            I => \N__29678\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__29684\,
            I => \N__29675\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__29681\,
            I => \N__29672\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__29678\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__3736\ : Odrv12
    port map (
            O => \N__29675\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__3735\ : Odrv4
    port map (
            O => \N__29672\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__3734\ : SRMux
    port map (
            O => \N__29665\,
            I => \N__29662\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__29662\,
            I => \N__29659\
        );

    \I__3732\ : Span4Mux_v
    port map (
            O => \N__29659\,
            I => \N__29656\
        );

    \I__3731\ : Odrv4
    port map (
            O => \N__29656\,
            I => \c0.n18601\
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__29653\,
            I => \c0.n6_adj_3143_cascade_\
        );

    \I__3729\ : InMux
    port map (
            O => \N__29650\,
            I => \N__29647\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__29647\,
            I => \N__29644\
        );

    \I__3727\ : Span4Mux_v
    port map (
            O => \N__29644\,
            I => \N__29641\
        );

    \I__3726\ : Sp12to4
    port map (
            O => \N__29641\,
            I => \N__29638\
        );

    \I__3725\ : Odrv12
    port map (
            O => \N__29638\,
            I => \c0.n4_adj_3227\
        );

    \I__3724\ : CascadeMux
    port map (
            O => \N__29635\,
            I => \N__29632\
        );

    \I__3723\ : InMux
    port map (
            O => \N__29632\,
            I => \N__29629\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__29629\,
            I => \c0.n19045\
        );

    \I__3721\ : InMux
    port map (
            O => \N__29626\,
            I => \N__29619\
        );

    \I__3720\ : InMux
    port map (
            O => \N__29625\,
            I => \N__29619\
        );

    \I__3719\ : InMux
    port map (
            O => \N__29624\,
            I => \N__29615\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__29619\,
            I => \N__29612\
        );

    \I__3717\ : InMux
    port map (
            O => \N__29618\,
            I => \N__29609\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__29615\,
            I => \N__29604\
        );

    \I__3715\ : Span4Mux_v
    port map (
            O => \N__29612\,
            I => \N__29604\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__29609\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__3713\ : Odrv4
    port map (
            O => \N__29604\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__3712\ : InMux
    port map (
            O => \N__29599\,
            I => \N__29595\
        );

    \I__3711\ : InMux
    port map (
            O => \N__29598\,
            I => \N__29592\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__29595\,
            I => \N__29585\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__29592\,
            I => \N__29585\
        );

    \I__3708\ : InMux
    port map (
            O => \N__29591\,
            I => \N__29582\
        );

    \I__3707\ : InMux
    port map (
            O => \N__29590\,
            I => \N__29579\
        );

    \I__3706\ : Span4Mux_h
    port map (
            O => \N__29585\,
            I => \N__29576\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__29582\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__29579\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__3703\ : Odrv4
    port map (
            O => \N__29576\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__3702\ : InMux
    port map (
            O => \N__29569\,
            I => \N__29563\
        );

    \I__3701\ : InMux
    port map (
            O => \N__29568\,
            I => \N__29563\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__29563\,
            I => \c0.n10_adj_3438\
        );

    \I__3699\ : InMux
    port map (
            O => \N__29560\,
            I => \N__29557\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__29557\,
            I => \c0.n19050\
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__29554\,
            I => \N__29550\
        );

    \I__3696\ : InMux
    port map (
            O => \N__29553\,
            I => \N__29545\
        );

    \I__3695\ : InMux
    port map (
            O => \N__29550\,
            I => \N__29540\
        );

    \I__3694\ : InMux
    port map (
            O => \N__29549\,
            I => \N__29540\
        );

    \I__3693\ : InMux
    port map (
            O => \N__29548\,
            I => \N__29537\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__29545\,
            I => \N__29532\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__29540\,
            I => \N__29532\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__29537\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__3689\ : Odrv12
    port map (
            O => \N__29532\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__3688\ : InMux
    port map (
            O => \N__29527\,
            I => \N__29524\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__29524\,
            I => \N__29520\
        );

    \I__3686\ : InMux
    port map (
            O => \N__29523\,
            I => \N__29517\
        );

    \I__3685\ : Span4Mux_h
    port map (
            O => \N__29520\,
            I => \N__29514\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__29517\,
            I => \c0.n63\
        );

    \I__3683\ : Odrv4
    port map (
            O => \N__29514\,
            I => \c0.n63\
        );

    \I__3682\ : InMux
    port map (
            O => \N__29509\,
            I => \N__29506\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__29506\,
            I => \N__29503\
        );

    \I__3680\ : Odrv12
    port map (
            O => \N__29503\,
            I => \c0.rx.r_Rx_Data_R\
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__29500\,
            I => \N__29497\
        );

    \I__3678\ : InMux
    port map (
            O => \N__29497\,
            I => \N__29492\
        );

    \I__3677\ : InMux
    port map (
            O => \N__29496\,
            I => \N__29489\
        );

    \I__3676\ : InMux
    port map (
            O => \N__29495\,
            I => \N__29486\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__29492\,
            I => \N__29483\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__29489\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__29486\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__3672\ : Odrv4
    port map (
            O => \N__29483\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__3671\ : SRMux
    port map (
            O => \N__29476\,
            I => \N__29473\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__29473\,
            I => \c0.n18659\
        );

    \I__3669\ : InMux
    port map (
            O => \N__29470\,
            I => \N__29466\
        );

    \I__3668\ : InMux
    port map (
            O => \N__29469\,
            I => \N__29463\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__29466\,
            I => \N__29460\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__29463\,
            I => \N__29457\
        );

    \I__3665\ : Odrv12
    port map (
            O => \N__29460\,
            I => \c0.n19146\
        );

    \I__3664\ : Odrv4
    port map (
            O => \N__29457\,
            I => \c0.n19146\
        );

    \I__3663\ : InMux
    port map (
            O => \N__29452\,
            I => \N__29447\
        );

    \I__3662\ : InMux
    port map (
            O => \N__29451\,
            I => \N__29442\
        );

    \I__3661\ : InMux
    port map (
            O => \N__29450\,
            I => \N__29442\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__29447\,
            I => \c0.FRAME_MATCHER_state_3\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__29442\,
            I => \c0.FRAME_MATCHER_state_3\
        );

    \I__3658\ : SRMux
    port map (
            O => \N__29437\,
            I => \N__29434\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__29434\,
            I => \N__29431\
        );

    \I__3656\ : Span4Mux_h
    port map (
            O => \N__29431\,
            I => \N__29428\
        );

    \I__3655\ : Odrv4
    port map (
            O => \N__29428\,
            I => \c0.n18633\
        );

    \I__3654\ : InMux
    port map (
            O => \N__29425\,
            I => \N__29420\
        );

    \I__3653\ : InMux
    port map (
            O => \N__29424\,
            I => \N__29417\
        );

    \I__3652\ : InMux
    port map (
            O => \N__29423\,
            I => \N__29414\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__29420\,
            I => \N__29411\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__29417\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__29414\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__3648\ : Odrv4
    port map (
            O => \N__29411\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__3647\ : InMux
    port map (
            O => \N__29404\,
            I => \N__29401\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__29401\,
            I => \N__29398\
        );

    \I__3645\ : Span4Mux_v
    port map (
            O => \N__29398\,
            I => \N__29393\
        );

    \I__3644\ : InMux
    port map (
            O => \N__29397\,
            I => \N__29390\
        );

    \I__3643\ : InMux
    port map (
            O => \N__29396\,
            I => \N__29387\
        );

    \I__3642\ : Span4Mux_h
    port map (
            O => \N__29393\,
            I => \N__29384\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__29390\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__29387\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__3639\ : Odrv4
    port map (
            O => \N__29384\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__3638\ : InMux
    port map (
            O => \N__29377\,
            I => \N__29374\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__29374\,
            I => \c0.n10_adj_3488\
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__29371\,
            I => \c0.n15850_cascade_\
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__29368\,
            I => \c0.n11427_cascade_\
        );

    \I__3634\ : InMux
    port map (
            O => \N__29365\,
            I => \N__29362\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__29362\,
            I => \N__29359\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__29359\,
            I => \c0.n16_adj_3484\
        );

    \I__3631\ : InMux
    port map (
            O => \N__29356\,
            I => \N__29351\
        );

    \I__3630\ : InMux
    port map (
            O => \N__29355\,
            I => \N__29348\
        );

    \I__3629\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29345\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__29351\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__29348\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__29345\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__3625\ : CascadeMux
    port map (
            O => \N__29338\,
            I => \c0.n19045_cascade_\
        );

    \I__3624\ : InMux
    port map (
            O => \N__29335\,
            I => \N__29332\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__29332\,
            I => \c0.n4_adj_3046\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__29329\,
            I => \N__29325\
        );

    \I__3621\ : InMux
    port map (
            O => \N__29328\,
            I => \N__29321\
        );

    \I__3620\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29316\
        );

    \I__3619\ : InMux
    port map (
            O => \N__29324\,
            I => \N__29316\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__29321\,
            I => \N__29313\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__29316\,
            I => \N__29310\
        );

    \I__3616\ : Odrv4
    port map (
            O => \N__29313\,
            I => \c0.n15920\
        );

    \I__3615\ : Odrv4
    port map (
            O => \N__29310\,
            I => \c0.n15920\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__29305\,
            I => \N__29299\
        );

    \I__3613\ : InMux
    port map (
            O => \N__29304\,
            I => \N__29295\
        );

    \I__3612\ : InMux
    port map (
            O => \N__29303\,
            I => \N__29292\
        );

    \I__3611\ : InMux
    port map (
            O => \N__29302\,
            I => \N__29285\
        );

    \I__3610\ : InMux
    port map (
            O => \N__29299\,
            I => \N__29285\
        );

    \I__3609\ : InMux
    port map (
            O => \N__29298\,
            I => \N__29285\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__29295\,
            I => \N__29273\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__29292\,
            I => \N__29273\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__29285\,
            I => \N__29273\
        );

    \I__3605\ : InMux
    port map (
            O => \N__29284\,
            I => \N__29264\
        );

    \I__3604\ : InMux
    port map (
            O => \N__29283\,
            I => \N__29264\
        );

    \I__3603\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29261\
        );

    \I__3602\ : InMux
    port map (
            O => \N__29281\,
            I => \N__29256\
        );

    \I__3601\ : InMux
    port map (
            O => \N__29280\,
            I => \N__29256\
        );

    \I__3600\ : Span4Mux_v
    port map (
            O => \N__29273\,
            I => \N__29253\
        );

    \I__3599\ : InMux
    port map (
            O => \N__29272\,
            I => \N__29244\
        );

    \I__3598\ : InMux
    port map (
            O => \N__29271\,
            I => \N__29244\
        );

    \I__3597\ : InMux
    port map (
            O => \N__29270\,
            I => \N__29244\
        );

    \I__3596\ : InMux
    port map (
            O => \N__29269\,
            I => \N__29244\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__29264\,
            I => \r_SM_Main_1_adj_3592\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__29261\,
            I => \r_SM_Main_1_adj_3592\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__29256\,
            I => \r_SM_Main_1_adj_3592\
        );

    \I__3592\ : Odrv4
    port map (
            O => \N__29253\,
            I => \r_SM_Main_1_adj_3592\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__29244\,
            I => \r_SM_Main_1_adj_3592\
        );

    \I__3590\ : InMux
    port map (
            O => \N__29233\,
            I => \N__29230\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__29230\,
            I => \N__29227\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__29227\,
            I => n4_adj_3580
        );

    \I__3587\ : InMux
    port map (
            O => \N__29224\,
            I => \N__29221\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__29221\,
            I => \N__29218\
        );

    \I__3585\ : Odrv4
    port map (
            O => \N__29218\,
            I => n9_adj_3591
        );

    \I__3584\ : InMux
    port map (
            O => \N__29215\,
            I => \N__29211\
        );

    \I__3583\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29208\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__29211\,
            I => \r_Tx_Data_4\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__29208\,
            I => \r_Tx_Data_4\
        );

    \I__3580\ : CEMux
    port map (
            O => \N__29203\,
            I => \N__29200\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__29200\,
            I => \N__29196\
        );

    \I__3578\ : CEMux
    port map (
            O => \N__29199\,
            I => \N__29193\
        );

    \I__3577\ : Span4Mux_v
    port map (
            O => \N__29196\,
            I => \N__29190\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__29193\,
            I => \N__29187\
        );

    \I__3575\ : Span4Mux_h
    port map (
            O => \N__29190\,
            I => \N__29183\
        );

    \I__3574\ : Sp12to4
    port map (
            O => \N__29187\,
            I => \N__29180\
        );

    \I__3573\ : InMux
    port map (
            O => \N__29186\,
            I => \N__29177\
        );

    \I__3572\ : Odrv4
    port map (
            O => \N__29183\,
            I => \c0.n12512\
        );

    \I__3571\ : Odrv12
    port map (
            O => \N__29180\,
            I => \c0.n12512\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__29177\,
            I => \c0.n12512\
        );

    \I__3569\ : CascadeMux
    port map (
            O => \N__29170\,
            I => \N__29165\
        );

    \I__3568\ : InMux
    port map (
            O => \N__29169\,
            I => \N__29149\
        );

    \I__3567\ : InMux
    port map (
            O => \N__29168\,
            I => \N__29149\
        );

    \I__3566\ : InMux
    port map (
            O => \N__29165\,
            I => \N__29149\
        );

    \I__3565\ : InMux
    port map (
            O => \N__29164\,
            I => \N__29149\
        );

    \I__3564\ : CascadeMux
    port map (
            O => \N__29163\,
            I => \N__29146\
        );

    \I__3563\ : InMux
    port map (
            O => \N__29162\,
            I => \N__29139\
        );

    \I__3562\ : InMux
    port map (
            O => \N__29161\,
            I => \N__29134\
        );

    \I__3561\ : InMux
    port map (
            O => \N__29160\,
            I => \N__29134\
        );

    \I__3560\ : InMux
    port map (
            O => \N__29159\,
            I => \N__29129\
        );

    \I__3559\ : InMux
    port map (
            O => \N__29158\,
            I => \N__29129\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__29149\,
            I => \N__29126\
        );

    \I__3557\ : InMux
    port map (
            O => \N__29146\,
            I => \N__29121\
        );

    \I__3556\ : InMux
    port map (
            O => \N__29145\,
            I => \N__29121\
        );

    \I__3555\ : InMux
    port map (
            O => \N__29144\,
            I => \N__29118\
        );

    \I__3554\ : InMux
    port map (
            O => \N__29143\,
            I => \N__29113\
        );

    \I__3553\ : InMux
    port map (
            O => \N__29142\,
            I => \N__29113\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__29139\,
            I => \N__29108\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__29134\,
            I => \N__29108\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__29129\,
            I => \N__29105\
        );

    \I__3549\ : Span4Mux_v
    port map (
            O => \N__29126\,
            I => \N__29102\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__29121\,
            I => \c0.r_SM_Main_0\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__29118\,
            I => \c0.r_SM_Main_0\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__29113\,
            I => \c0.r_SM_Main_0\
        );

    \I__3545\ : Odrv4
    port map (
            O => \N__29108\,
            I => \c0.r_SM_Main_0\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__29105\,
            I => \c0.r_SM_Main_0\
        );

    \I__3543\ : Odrv4
    port map (
            O => \N__29102\,
            I => \c0.r_SM_Main_0\
        );

    \I__3542\ : InMux
    port map (
            O => \N__29089\,
            I => \N__29086\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__29086\,
            I => \c0.n19023\
        );

    \I__3540\ : SRMux
    port map (
            O => \N__29083\,
            I => \N__29080\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__29080\,
            I => \N__29077\
        );

    \I__3538\ : Sp12to4
    port map (
            O => \N__29077\,
            I => \N__29074\
        );

    \I__3537\ : Odrv12
    port map (
            O => \N__29074\,
            I => \c0.n18609\
        );

    \I__3536\ : InMux
    port map (
            O => \N__29071\,
            I => \N__29068\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__29068\,
            I => \N__29065\
        );

    \I__3534\ : Span4Mux_h
    port map (
            O => \N__29065\,
            I => \N__29062\
        );

    \I__3533\ : Odrv4
    port map (
            O => \N__29062\,
            I => \c0.n21456\
        );

    \I__3532\ : InMux
    port map (
            O => \N__29059\,
            I => \N__29052\
        );

    \I__3531\ : InMux
    port map (
            O => \N__29058\,
            I => \N__29043\
        );

    \I__3530\ : InMux
    port map (
            O => \N__29057\,
            I => \N__29043\
        );

    \I__3529\ : InMux
    port map (
            O => \N__29056\,
            I => \N__29043\
        );

    \I__3528\ : InMux
    port map (
            O => \N__29055\,
            I => \N__29043\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__29052\,
            I => \c0.r_Bit_Index_1\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__29043\,
            I => \c0.r_Bit_Index_1\
        );

    \I__3525\ : InMux
    port map (
            O => \N__29038\,
            I => \N__29035\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__29035\,
            I => \c0.n21614\
        );

    \I__3523\ : InMux
    port map (
            O => \N__29032\,
            I => \N__29029\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__29029\,
            I => \N__29026\
        );

    \I__3521\ : Odrv4
    port map (
            O => \N__29026\,
            I => \c0.n32\
        );

    \I__3520\ : CascadeMux
    port map (
            O => \N__29023\,
            I => \c0.n2_adj_3556_cascade_\
        );

    \I__3519\ : InMux
    port map (
            O => \N__29020\,
            I => \N__29017\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__29017\,
            I => \c0.n7_adj_3557\
        );

    \I__3517\ : InMux
    port map (
            O => \N__29014\,
            I => \N__29011\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__29011\,
            I => \c0.n21329\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__29008\,
            I => \c0.n19001_cascade_\
        );

    \I__3514\ : InMux
    port map (
            O => \N__29005\,
            I => \N__29002\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__29002\,
            I => \N__28999\
        );

    \I__3512\ : Span4Mux_v
    port map (
            O => \N__28999\,
            I => \N__28996\
        );

    \I__3511\ : Odrv4
    port map (
            O => \N__28996\,
            I => \c0.n30_adj_3559\
        );

    \I__3510\ : CascadeMux
    port map (
            O => \N__28993\,
            I => \N__28989\
        );

    \I__3509\ : InMux
    port map (
            O => \N__28992\,
            I => \N__28985\
        );

    \I__3508\ : InMux
    port map (
            O => \N__28989\,
            I => \N__28980\
        );

    \I__3507\ : InMux
    port map (
            O => \N__28988\,
            I => \N__28980\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__28985\,
            I => \c0.n12498\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__28980\,
            I => \c0.n12498\
        );

    \I__3504\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28972\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__28972\,
            I => \c0.n21577\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__28969\,
            I => \n21578_cascade_\
        );

    \I__3501\ : InMux
    port map (
            O => \N__28966\,
            I => \N__28963\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__28963\,
            I => n21656
        );

    \I__3499\ : InMux
    port map (
            O => \N__28960\,
            I => \N__28956\
        );

    \I__3498\ : InMux
    port map (
            O => \N__28959\,
            I => \N__28953\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__28956\,
            I => \N__28950\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__28953\,
            I => data_out_frame_13_7
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__28950\,
            I => data_out_frame_13_7
        );

    \I__3494\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28942\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__28942\,
            I => \c0.n21467\
        );

    \I__3492\ : InMux
    port map (
            O => \N__28939\,
            I => \N__28936\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__28936\,
            I => \N__28933\
        );

    \I__3490\ : Span4Mux_h
    port map (
            O => \N__28933\,
            I => \N__28930\
        );

    \I__3489\ : Odrv4
    port map (
            O => \N__28930\,
            I => \c0.tx.n21330\
        );

    \I__3488\ : InMux
    port map (
            O => \N__28927\,
            I => \N__28924\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__28924\,
            I => n9_adj_3588
        );

    \I__3486\ : InMux
    port map (
            O => \N__28921\,
            I => \N__28915\
        );

    \I__3485\ : InMux
    port map (
            O => \N__28920\,
            I => \N__28915\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__28915\,
            I => \r_Tx_Data_6\
        );

    \I__3483\ : CascadeMux
    port map (
            O => \N__28912\,
            I => \c0.n9753_cascade_\
        );

    \I__3482\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28905\
        );

    \I__3481\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28902\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__28905\,
            I => \N__28899\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__28902\,
            I => data_out_frame_12_3
        );

    \I__3478\ : Odrv4
    port map (
            O => \N__28899\,
            I => data_out_frame_12_3
        );

    \I__3477\ : CascadeMux
    port map (
            O => \N__28894\,
            I => \N__28891\
        );

    \I__3476\ : InMux
    port map (
            O => \N__28891\,
            I => \N__28885\
        );

    \I__3475\ : InMux
    port map (
            O => \N__28890\,
            I => \N__28885\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__28885\,
            I => data_out_frame_13_3
        );

    \I__3473\ : InMux
    port map (
            O => \N__28882\,
            I => \N__28878\
        );

    \I__3472\ : InMux
    port map (
            O => \N__28881\,
            I => \N__28875\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__28878\,
            I => data_out_frame_12_7
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__28875\,
            I => data_out_frame_12_7
        );

    \I__3469\ : CascadeMux
    port map (
            O => \N__28870\,
            I => \N__28866\
        );

    \I__3468\ : InMux
    port map (
            O => \N__28869\,
            I => \N__28863\
        );

    \I__3467\ : InMux
    port map (
            O => \N__28866\,
            I => \N__28860\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__28863\,
            I => data_out_frame_11_3
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__28860\,
            I => data_out_frame_11_3
        );

    \I__3464\ : InMux
    port map (
            O => \N__28855\,
            I => \N__28849\
        );

    \I__3463\ : InMux
    port map (
            O => \N__28854\,
            I => \N__28849\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__28849\,
            I => data_out_frame_10_3
        );

    \I__3461\ : InMux
    port map (
            O => \N__28846\,
            I => \N__28843\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__28843\,
            I => \N__28839\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__28842\,
            I => \N__28835\
        );

    \I__3458\ : Span4Mux_h
    port map (
            O => \N__28839\,
            I => \N__28832\
        );

    \I__3457\ : InMux
    port map (
            O => \N__28838\,
            I => \N__28829\
        );

    \I__3456\ : InMux
    port map (
            O => \N__28835\,
            I => \N__28826\
        );

    \I__3455\ : Span4Mux_v
    port map (
            O => \N__28832\,
            I => \N__28819\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__28829\,
            I => \N__28819\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__28826\,
            I => \N__28819\
        );

    \I__3452\ : Odrv4
    port map (
            O => \N__28819\,
            I => encoder0_position_12
        );

    \I__3451\ : InMux
    port map (
            O => \N__28816\,
            I => \N__28812\
        );

    \I__3450\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28809\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__28812\,
            I => data_out_frame_13_6
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__28809\,
            I => data_out_frame_13_6
        );

    \I__3447\ : InMux
    port map (
            O => \N__28804\,
            I => \N__28801\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__28801\,
            I => \c0.n21301\
        );

    \I__3445\ : InMux
    port map (
            O => \N__28798\,
            I => \N__28795\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__28795\,
            I => \N__28792\
        );

    \I__3443\ : Odrv4
    port map (
            O => \N__28792\,
            I => \c0.n21653\
        );

    \I__3442\ : InMux
    port map (
            O => \N__28789\,
            I => \N__28786\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__28786\,
            I => \N__28783\
        );

    \I__3440\ : Span4Mux_h
    port map (
            O => \N__28783\,
            I => \N__28780\
        );

    \I__3439\ : Odrv4
    port map (
            O => \N__28780\,
            I => \c0.n21305\
        );

    \I__3438\ : InMux
    port map (
            O => \N__28777\,
            I => \N__28774\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__28774\,
            I => \c0.n21570\
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__28771\,
            I => \c0.n21307_cascade_\
        );

    \I__3435\ : InMux
    port map (
            O => \N__28768\,
            I => \N__28764\
        );

    \I__3434\ : InMux
    port map (
            O => \N__28767\,
            I => \N__28761\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__28764\,
            I => \N__28758\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__28761\,
            I => data_out_frame_11_4
        );

    \I__3431\ : Odrv4
    port map (
            O => \N__28758\,
            I => data_out_frame_11_4
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__28753\,
            I => \N__28750\
        );

    \I__3429\ : InMux
    port map (
            O => \N__28750\,
            I => \N__28747\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__28747\,
            I => \N__28744\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__28744\,
            I => \c0.n5_adj_3033\
        );

    \I__3426\ : InMux
    port map (
            O => \N__28741\,
            I => \N__28737\
        );

    \I__3425\ : InMux
    port map (
            O => \N__28740\,
            I => \N__28734\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__28737\,
            I => \N__28731\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__28734\,
            I => data_out_frame_12_6
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__28731\,
            I => data_out_frame_12_6
        );

    \I__3421\ : InMux
    port map (
            O => \N__28726\,
            I => \N__28722\
        );

    \I__3420\ : InMux
    port map (
            O => \N__28725\,
            I => \N__28718\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__28722\,
            I => \N__28715\
        );

    \I__3418\ : InMux
    port map (
            O => \N__28721\,
            I => \N__28712\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__28718\,
            I => encoder0_position_17
        );

    \I__3416\ : Odrv4
    port map (
            O => \N__28715\,
            I => encoder0_position_17
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__28712\,
            I => encoder0_position_17
        );

    \I__3414\ : InMux
    port map (
            O => \N__28705\,
            I => \N__28701\
        );

    \I__3413\ : InMux
    port map (
            O => \N__28704\,
            I => \N__28698\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__28701\,
            I => data_out_frame_7_1
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__28698\,
            I => data_out_frame_7_1
        );

    \I__3410\ : InMux
    port map (
            O => \N__28693\,
            I => \N__28690\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__28690\,
            I => \c0.n6_adj_3324\
        );

    \I__3408\ : InMux
    port map (
            O => \N__28687\,
            I => \N__28684\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__28684\,
            I => \N__28681\
        );

    \I__3406\ : Odrv4
    port map (
            O => \N__28681\,
            I => n2250
        );

    \I__3405\ : InMux
    port map (
            O => \N__28678\,
            I => \N__28675\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__28675\,
            I => \N__28670\
        );

    \I__3403\ : CascadeMux
    port map (
            O => \N__28674\,
            I => \N__28667\
        );

    \I__3402\ : InMux
    port map (
            O => \N__28673\,
            I => \N__28664\
        );

    \I__3401\ : Span4Mux_v
    port map (
            O => \N__28670\,
            I => \N__28661\
        );

    \I__3400\ : InMux
    port map (
            O => \N__28667\,
            I => \N__28658\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__28664\,
            I => encoder0_position_13
        );

    \I__3398\ : Odrv4
    port map (
            O => \N__28661\,
            I => encoder0_position_13
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__28658\,
            I => encoder0_position_13
        );

    \I__3396\ : CascadeMux
    port map (
            O => \N__28651\,
            I => \N__28648\
        );

    \I__3395\ : InMux
    port map (
            O => \N__28648\,
            I => \N__28645\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__28645\,
            I => \N__28641\
        );

    \I__3393\ : InMux
    port map (
            O => \N__28644\,
            I => \N__28638\
        );

    \I__3392\ : Span4Mux_h
    port map (
            O => \N__28641\,
            I => \N__28635\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__28638\,
            I => data_out_frame_11_6
        );

    \I__3390\ : Odrv4
    port map (
            O => \N__28635\,
            I => data_out_frame_11_6
        );

    \I__3389\ : InMux
    port map (
            O => \N__28630\,
            I => \N__28627\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__28627\,
            I => \N__28624\
        );

    \I__3387\ : Span4Mux_v
    port map (
            O => \N__28624\,
            I => \N__28621\
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__28621\,
            I => n2271
        );

    \I__3385\ : InMux
    port map (
            O => \N__28618\,
            I => \N__28615\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__28615\,
            I => \c0.n21650\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__28612\,
            I => \c0.n21564_cascade_\
        );

    \I__3382\ : InMux
    port map (
            O => \N__28609\,
            I => \N__28606\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__28606\,
            I => \N__28603\
        );

    \I__3380\ : Span4Mux_h
    port map (
            O => \N__28603\,
            I => \N__28600\
        );

    \I__3379\ : Odrv4
    port map (
            O => \N__28600\,
            I => n2270
        );

    \I__3378\ : CascadeMux
    port map (
            O => \N__28597\,
            I => \N__28593\
        );

    \I__3377\ : InMux
    port map (
            O => \N__28596\,
            I => \N__28590\
        );

    \I__3376\ : InMux
    port map (
            O => \N__28593\,
            I => \N__28587\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__28590\,
            I => \quad_counter1.a_delay_counter_11\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__28587\,
            I => \quad_counter1.a_delay_counter_11\
        );

    \I__3373\ : InMux
    port map (
            O => \N__28582\,
            I => \quad_counter1.n17262\
        );

    \I__3372\ : InMux
    port map (
            O => \N__28579\,
            I => \N__28575\
        );

    \I__3371\ : InMux
    port map (
            O => \N__28578\,
            I => \N__28572\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__28575\,
            I => \quad_counter1.a_delay_counter_12\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__28572\,
            I => \quad_counter1.a_delay_counter_12\
        );

    \I__3368\ : InMux
    port map (
            O => \N__28567\,
            I => \quad_counter1.n17263\
        );

    \I__3367\ : InMux
    port map (
            O => \N__28564\,
            I => \N__28560\
        );

    \I__3366\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28557\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__28560\,
            I => \quad_counter1.a_delay_counter_13\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__28557\,
            I => \quad_counter1.a_delay_counter_13\
        );

    \I__3363\ : InMux
    port map (
            O => \N__28552\,
            I => \quad_counter1.n17264\
        );

    \I__3362\ : InMux
    port map (
            O => \N__28549\,
            I => \N__28545\
        );

    \I__3361\ : InMux
    port map (
            O => \N__28548\,
            I => \N__28542\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__28545\,
            I => \quad_counter1.a_delay_counter_14\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__28542\,
            I => \quad_counter1.a_delay_counter_14\
        );

    \I__3358\ : InMux
    port map (
            O => \N__28537\,
            I => \quad_counter1.n17265\
        );

    \I__3357\ : InMux
    port map (
            O => \N__28534\,
            I => \quad_counter1.n17266\
        );

    \I__3356\ : InMux
    port map (
            O => \N__28531\,
            I => \N__28527\
        );

    \I__3355\ : InMux
    port map (
            O => \N__28530\,
            I => \N__28524\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__28527\,
            I => \quad_counter1.a_delay_counter_15\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__28524\,
            I => \quad_counter1.a_delay_counter_15\
        );

    \I__3352\ : CEMux
    port map (
            O => \N__28519\,
            I => \N__28516\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__28516\,
            I => \N__28512\
        );

    \I__3350\ : CEMux
    port map (
            O => \N__28515\,
            I => \N__28509\
        );

    \I__3349\ : Span4Mux_h
    port map (
            O => \N__28512\,
            I => \N__28505\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__28509\,
            I => \N__28502\
        );

    \I__3347\ : InMux
    port map (
            O => \N__28508\,
            I => \N__28499\
        );

    \I__3346\ : Odrv4
    port map (
            O => \N__28505\,
            I => n12477
        );

    \I__3345\ : Odrv4
    port map (
            O => \N__28502\,
            I => n12477
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__28499\,
            I => n12477
        );

    \I__3343\ : SRMux
    port map (
            O => \N__28492\,
            I => \N__28488\
        );

    \I__3342\ : SRMux
    port map (
            O => \N__28491\,
            I => \N__28485\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__28488\,
            I => \N__28482\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__28485\,
            I => \N__28479\
        );

    \I__3339\ : Odrv12
    port map (
            O => \N__28482\,
            I => \a_delay_counter_15__N_2916_adj_3589\
        );

    \I__3338\ : Odrv4
    port map (
            O => \N__28479\,
            I => \a_delay_counter_15__N_2916_adj_3589\
        );

    \I__3337\ : InMux
    port map (
            O => \N__28474\,
            I => \N__28470\
        );

    \I__3336\ : InMux
    port map (
            O => \N__28473\,
            I => \N__28467\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__28470\,
            I => \N__28464\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__28467\,
            I => data_out_frame_9_2
        );

    \I__3333\ : Odrv4
    port map (
            O => \N__28464\,
            I => data_out_frame_9_2
        );

    \I__3332\ : InMux
    port map (
            O => \N__28459\,
            I => \N__28455\
        );

    \I__3331\ : InMux
    port map (
            O => \N__28458\,
            I => \N__28452\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__28455\,
            I => data_out_frame_8_2
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__28452\,
            I => data_out_frame_8_2
        );

    \I__3328\ : InMux
    port map (
            O => \N__28447\,
            I => \quad_counter1.n17253\
        );

    \I__3327\ : InMux
    port map (
            O => \N__28444\,
            I => \N__28440\
        );

    \I__3326\ : InMux
    port map (
            O => \N__28443\,
            I => \N__28437\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__28440\,
            I => \quad_counter1.a_delay_counter_3\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__28437\,
            I => \quad_counter1.a_delay_counter_3\
        );

    \I__3323\ : InMux
    port map (
            O => \N__28432\,
            I => \quad_counter1.n17254\
        );

    \I__3322\ : InMux
    port map (
            O => \N__28429\,
            I => \N__28425\
        );

    \I__3321\ : InMux
    port map (
            O => \N__28428\,
            I => \N__28422\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__28425\,
            I => \quad_counter1.a_delay_counter_4\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__28422\,
            I => \quad_counter1.a_delay_counter_4\
        );

    \I__3318\ : InMux
    port map (
            O => \N__28417\,
            I => \quad_counter1.n17255\
        );

    \I__3317\ : InMux
    port map (
            O => \N__28414\,
            I => \N__28410\
        );

    \I__3316\ : InMux
    port map (
            O => \N__28413\,
            I => \N__28407\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__28410\,
            I => \quad_counter1.a_delay_counter_5\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__28407\,
            I => \quad_counter1.a_delay_counter_5\
        );

    \I__3313\ : InMux
    port map (
            O => \N__28402\,
            I => \quad_counter1.n17256\
        );

    \I__3312\ : InMux
    port map (
            O => \N__28399\,
            I => \N__28395\
        );

    \I__3311\ : InMux
    port map (
            O => \N__28398\,
            I => \N__28392\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__28395\,
            I => \quad_counter1.a_delay_counter_6\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__28392\,
            I => \quad_counter1.a_delay_counter_6\
        );

    \I__3308\ : InMux
    port map (
            O => \N__28387\,
            I => \quad_counter1.n17257\
        );

    \I__3307\ : InMux
    port map (
            O => \N__28384\,
            I => \N__28380\
        );

    \I__3306\ : InMux
    port map (
            O => \N__28383\,
            I => \N__28377\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__28380\,
            I => \quad_counter1.a_delay_counter_7\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__28377\,
            I => \quad_counter1.a_delay_counter_7\
        );

    \I__3303\ : InMux
    port map (
            O => \N__28372\,
            I => \quad_counter1.n17258\
        );

    \I__3302\ : CascadeMux
    port map (
            O => \N__28369\,
            I => \N__28365\
        );

    \I__3301\ : InMux
    port map (
            O => \N__28368\,
            I => \N__28362\
        );

    \I__3300\ : InMux
    port map (
            O => \N__28365\,
            I => \N__28359\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__28362\,
            I => \quad_counter1.a_delay_counter_8\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__28359\,
            I => \quad_counter1.a_delay_counter_8\
        );

    \I__3297\ : InMux
    port map (
            O => \N__28354\,
            I => \bfn_12_9_0_\
        );

    \I__3296\ : InMux
    port map (
            O => \N__28351\,
            I => \N__28347\
        );

    \I__3295\ : InMux
    port map (
            O => \N__28350\,
            I => \N__28344\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__28347\,
            I => \N__28341\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__28344\,
            I => \quad_counter1.a_delay_counter_9\
        );

    \I__3292\ : Odrv4
    port map (
            O => \N__28341\,
            I => \quad_counter1.a_delay_counter_9\
        );

    \I__3291\ : InMux
    port map (
            O => \N__28336\,
            I => \quad_counter1.n17260\
        );

    \I__3290\ : InMux
    port map (
            O => \N__28333\,
            I => \N__28329\
        );

    \I__3289\ : InMux
    port map (
            O => \N__28332\,
            I => \N__28326\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__28329\,
            I => \quad_counter1.a_delay_counter_10\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__28326\,
            I => \quad_counter1.a_delay_counter_10\
        );

    \I__3286\ : InMux
    port map (
            O => \N__28321\,
            I => \quad_counter1.n17261\
        );

    \I__3285\ : InMux
    port map (
            O => \N__28318\,
            I => \N__28314\
        );

    \I__3284\ : InMux
    port map (
            O => \N__28317\,
            I => \N__28311\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__28314\,
            I => \quad_counter1.b_delay_counter_13\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__28311\,
            I => \quad_counter1.b_delay_counter_13\
        );

    \I__3281\ : InMux
    port map (
            O => \N__28306\,
            I => \quad_counter1.n17249\
        );

    \I__3280\ : InMux
    port map (
            O => \N__28303\,
            I => \N__28299\
        );

    \I__3279\ : InMux
    port map (
            O => \N__28302\,
            I => \N__28296\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__28299\,
            I => \quad_counter1.b_delay_counter_14\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__28296\,
            I => \quad_counter1.b_delay_counter_14\
        );

    \I__3276\ : InMux
    port map (
            O => \N__28291\,
            I => \quad_counter1.n17250\
        );

    \I__3275\ : InMux
    port map (
            O => \N__28288\,
            I => \quad_counter1.n17251\
        );

    \I__3274\ : InMux
    port map (
            O => \N__28285\,
            I => \N__28281\
        );

    \I__3273\ : InMux
    port map (
            O => \N__28284\,
            I => \N__28278\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__28281\,
            I => \quad_counter1.b_delay_counter_15\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__28278\,
            I => \quad_counter1.b_delay_counter_15\
        );

    \I__3270\ : CEMux
    port map (
            O => \N__28273\,
            I => \N__28270\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__28270\,
            I => \N__28267\
        );

    \I__3268\ : Span4Mux_v
    port map (
            O => \N__28267\,
            I => \N__28263\
        );

    \I__3267\ : CEMux
    port map (
            O => \N__28266\,
            I => \N__28260\
        );

    \I__3266\ : Span4Mux_s2_v
    port map (
            O => \N__28263\,
            I => \N__28255\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__28260\,
            I => \N__28255\
        );

    \I__3264\ : Span4Mux_v
    port map (
            O => \N__28255\,
            I => \N__28252\
        );

    \I__3263\ : Span4Mux_s2_v
    port map (
            O => \N__28252\,
            I => \N__28249\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__28249\,
            I => n12417
        );

    \I__3261\ : SRMux
    port map (
            O => \N__28246\,
            I => \N__28241\
        );

    \I__3260\ : InMux
    port map (
            O => \N__28245\,
            I => \N__28238\
        );

    \I__3259\ : SRMux
    port map (
            O => \N__28244\,
            I => \N__28235\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__28241\,
            I => \N__28232\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__28238\,
            I => \N__28228\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__28235\,
            I => \N__28223\
        );

    \I__3255\ : Span4Mux_v
    port map (
            O => \N__28232\,
            I => \N__28223\
        );

    \I__3254\ : InMux
    port map (
            O => \N__28231\,
            I => \N__28220\
        );

    \I__3253\ : Odrv4
    port map (
            O => \N__28228\,
            I => \b_delay_counter_15__N_2933\
        );

    \I__3252\ : Odrv4
    port map (
            O => \N__28223\,
            I => \b_delay_counter_15__N_2933\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__28220\,
            I => \b_delay_counter_15__N_2933\
        );

    \I__3250\ : InMux
    port map (
            O => \N__28213\,
            I => \N__28207\
        );

    \I__3249\ : InMux
    port map (
            O => \N__28212\,
            I => \N__28207\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__28207\,
            I => \N__28202\
        );

    \I__3247\ : InMux
    port map (
            O => \N__28206\,
            I => \N__28199\
        );

    \I__3246\ : InMux
    port map (
            O => \N__28205\,
            I => \N__28196\
        );

    \I__3245\ : Span4Mux_v
    port map (
            O => \N__28202\,
            I => \N__28191\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__28199\,
            I => \N__28191\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__28196\,
            I => \N__28188\
        );

    \I__3242\ : IoSpan4Mux
    port map (
            O => \N__28191\,
            I => \N__28185\
        );

    \I__3241\ : Span12Mux_h
    port map (
            O => \N__28188\,
            I => \N__28182\
        );

    \I__3240\ : IoSpan4Mux
    port map (
            O => \N__28185\,
            I => \N__28179\
        );

    \I__3239\ : Odrv12
    port map (
            O => \N__28182\,
            I => \PIN_12_c\
        );

    \I__3238\ : Odrv4
    port map (
            O => \N__28179\,
            I => \PIN_12_c\
        );

    \I__3237\ : CascadeMux
    port map (
            O => \N__28174\,
            I => \N__28171\
        );

    \I__3236\ : InMux
    port map (
            O => \N__28171\,
            I => \N__28164\
        );

    \I__3235\ : InMux
    port map (
            O => \N__28170\,
            I => \N__28164\
        );

    \I__3234\ : InMux
    port map (
            O => \N__28169\,
            I => \N__28161\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__28164\,
            I => \N__28156\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__28161\,
            I => \N__28156\
        );

    \I__3231\ : Span4Mux_h
    port map (
            O => \N__28156\,
            I => \N__28153\
        );

    \I__3230\ : Odrv4
    port map (
            O => \N__28153\,
            I => \quadA_delayed_adj_3584\
        );

    \I__3229\ : CascadeMux
    port map (
            O => \N__28150\,
            I => \a_delay_counter_15__N_2916_adj_3589_cascade_\
        );

    \I__3228\ : InMux
    port map (
            O => \N__28147\,
            I => \N__28144\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__28144\,
            I => \quad_counter1.n20\
        );

    \I__3226\ : InMux
    port map (
            O => \N__28141\,
            I => \N__28136\
        );

    \I__3225\ : InMux
    port map (
            O => \N__28140\,
            I => \N__28131\
        );

    \I__3224\ : InMux
    port map (
            O => \N__28139\,
            I => \N__28131\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__28136\,
            I => a_delay_counter_0_adj_3583
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__28131\,
            I => a_delay_counter_0_adj_3583
        );

    \I__3221\ : InMux
    port map (
            O => \N__28126\,
            I => \N__28123\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__28123\,
            I => n39_adj_3587
        );

    \I__3219\ : InMux
    port map (
            O => \N__28120\,
            I => \bfn_12_8_0_\
        );

    \I__3218\ : InMux
    port map (
            O => \N__28117\,
            I => \N__28113\
        );

    \I__3217\ : InMux
    port map (
            O => \N__28116\,
            I => \N__28110\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__28113\,
            I => \quad_counter1.a_delay_counter_1\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__28110\,
            I => \quad_counter1.a_delay_counter_1\
        );

    \I__3214\ : InMux
    port map (
            O => \N__28105\,
            I => \quad_counter1.n17252\
        );

    \I__3213\ : InMux
    port map (
            O => \N__28102\,
            I => \N__28098\
        );

    \I__3212\ : InMux
    port map (
            O => \N__28101\,
            I => \N__28095\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__28098\,
            I => \quad_counter1.a_delay_counter_2\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__28095\,
            I => \quad_counter1.a_delay_counter_2\
        );

    \I__3209\ : InMux
    port map (
            O => \N__28090\,
            I => \N__28086\
        );

    \I__3208\ : InMux
    port map (
            O => \N__28089\,
            I => \N__28083\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__28086\,
            I => \quad_counter1.b_delay_counter_5\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__28083\,
            I => \quad_counter1.b_delay_counter_5\
        );

    \I__3205\ : InMux
    port map (
            O => \N__28078\,
            I => \quad_counter1.n17241\
        );

    \I__3204\ : CascadeMux
    port map (
            O => \N__28075\,
            I => \N__28071\
        );

    \I__3203\ : InMux
    port map (
            O => \N__28074\,
            I => \N__28068\
        );

    \I__3202\ : InMux
    port map (
            O => \N__28071\,
            I => \N__28065\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__28068\,
            I => \quad_counter1.b_delay_counter_6\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__28065\,
            I => \quad_counter1.b_delay_counter_6\
        );

    \I__3199\ : InMux
    port map (
            O => \N__28060\,
            I => \quad_counter1.n17242\
        );

    \I__3198\ : InMux
    port map (
            O => \N__28057\,
            I => \N__28053\
        );

    \I__3197\ : InMux
    port map (
            O => \N__28056\,
            I => \N__28050\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__28053\,
            I => \quad_counter1.b_delay_counter_7\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__28050\,
            I => \quad_counter1.b_delay_counter_7\
        );

    \I__3194\ : InMux
    port map (
            O => \N__28045\,
            I => \quad_counter1.n17243\
        );

    \I__3193\ : InMux
    port map (
            O => \N__28042\,
            I => \N__28038\
        );

    \I__3192\ : InMux
    port map (
            O => \N__28041\,
            I => \N__28035\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__28038\,
            I => \quad_counter1.b_delay_counter_8\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__28035\,
            I => \quad_counter1.b_delay_counter_8\
        );

    \I__3189\ : InMux
    port map (
            O => \N__28030\,
            I => \bfn_12_6_0_\
        );

    \I__3188\ : InMux
    port map (
            O => \N__28027\,
            I => \N__28023\
        );

    \I__3187\ : InMux
    port map (
            O => \N__28026\,
            I => \N__28020\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__28023\,
            I => \quad_counter1.b_delay_counter_9\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__28020\,
            I => \quad_counter1.b_delay_counter_9\
        );

    \I__3184\ : InMux
    port map (
            O => \N__28015\,
            I => \quad_counter1.n17245\
        );

    \I__3183\ : InMux
    port map (
            O => \N__28012\,
            I => \N__28008\
        );

    \I__3182\ : InMux
    port map (
            O => \N__28011\,
            I => \N__28005\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__28008\,
            I => \quad_counter1.b_delay_counter_10\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__28005\,
            I => \quad_counter1.b_delay_counter_10\
        );

    \I__3179\ : InMux
    port map (
            O => \N__28000\,
            I => \quad_counter1.n17246\
        );

    \I__3178\ : InMux
    port map (
            O => \N__27997\,
            I => \N__27993\
        );

    \I__3177\ : InMux
    port map (
            O => \N__27996\,
            I => \N__27990\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__27993\,
            I => \quad_counter1.b_delay_counter_11\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__27990\,
            I => \quad_counter1.b_delay_counter_11\
        );

    \I__3174\ : InMux
    port map (
            O => \N__27985\,
            I => \quad_counter1.n17247\
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__27982\,
            I => \N__27978\
        );

    \I__3172\ : InMux
    port map (
            O => \N__27981\,
            I => \N__27975\
        );

    \I__3171\ : InMux
    port map (
            O => \N__27978\,
            I => \N__27972\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__27975\,
            I => \quad_counter1.b_delay_counter_12\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__27972\,
            I => \quad_counter1.b_delay_counter_12\
        );

    \I__3168\ : InMux
    port map (
            O => \N__27967\,
            I => \quad_counter1.n17248\
        );

    \I__3167\ : SRMux
    port map (
            O => \N__27964\,
            I => \N__27961\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__27961\,
            I => \N__27958\
        );

    \I__3165\ : Span4Mux_h
    port map (
            O => \N__27958\,
            I => \N__27955\
        );

    \I__3164\ : Odrv4
    port map (
            O => \N__27955\,
            I => \c0.n18651\
        );

    \I__3163\ : SRMux
    port map (
            O => \N__27952\,
            I => \N__27949\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__27949\,
            I => \N__27946\
        );

    \I__3161\ : Span4Mux_h
    port map (
            O => \N__27946\,
            I => \N__27943\
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__27943\,
            I => \c0.n18625\
        );

    \I__3159\ : SRMux
    port map (
            O => \N__27940\,
            I => \N__27937\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__27937\,
            I => \N__27934\
        );

    \I__3157\ : Span4Mux_h
    port map (
            O => \N__27934\,
            I => \N__27931\
        );

    \I__3156\ : Odrv4
    port map (
            O => \N__27931\,
            I => \c0.n18641\
        );

    \I__3155\ : InMux
    port map (
            O => \N__27928\,
            I => \N__27923\
        );

    \I__3154\ : InMux
    port map (
            O => \N__27927\,
            I => \N__27918\
        );

    \I__3153\ : InMux
    port map (
            O => \N__27926\,
            I => \N__27918\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__27923\,
            I => b_delay_counter_0
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__27918\,
            I => b_delay_counter_0
        );

    \I__3150\ : InMux
    port map (
            O => \N__27913\,
            I => \N__27910\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__27910\,
            I => n187
        );

    \I__3148\ : InMux
    port map (
            O => \N__27907\,
            I => \bfn_12_5_0_\
        );

    \I__3147\ : CascadeMux
    port map (
            O => \N__27904\,
            I => \N__27900\
        );

    \I__3146\ : InMux
    port map (
            O => \N__27903\,
            I => \N__27897\
        );

    \I__3145\ : InMux
    port map (
            O => \N__27900\,
            I => \N__27894\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__27897\,
            I => \quad_counter1.b_delay_counter_1\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__27894\,
            I => \quad_counter1.b_delay_counter_1\
        );

    \I__3142\ : InMux
    port map (
            O => \N__27889\,
            I => \quad_counter1.n17237\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__27886\,
            I => \N__27882\
        );

    \I__3140\ : InMux
    port map (
            O => \N__27885\,
            I => \N__27879\
        );

    \I__3139\ : InMux
    port map (
            O => \N__27882\,
            I => \N__27876\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__27879\,
            I => \quad_counter1.b_delay_counter_2\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__27876\,
            I => \quad_counter1.b_delay_counter_2\
        );

    \I__3136\ : InMux
    port map (
            O => \N__27871\,
            I => \quad_counter1.n17238\
        );

    \I__3135\ : InMux
    port map (
            O => \N__27868\,
            I => \N__27864\
        );

    \I__3134\ : InMux
    port map (
            O => \N__27867\,
            I => \N__27861\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__27864\,
            I => \quad_counter1.b_delay_counter_3\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__27861\,
            I => \quad_counter1.b_delay_counter_3\
        );

    \I__3131\ : InMux
    port map (
            O => \N__27856\,
            I => \quad_counter1.n17239\
        );

    \I__3130\ : InMux
    port map (
            O => \N__27853\,
            I => \N__27849\
        );

    \I__3129\ : InMux
    port map (
            O => \N__27852\,
            I => \N__27846\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__27849\,
            I => \quad_counter1.b_delay_counter_4\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__27846\,
            I => \quad_counter1.b_delay_counter_4\
        );

    \I__3126\ : InMux
    port map (
            O => \N__27841\,
            I => \quad_counter1.n17240\
        );

    \I__3125\ : SRMux
    port map (
            O => \N__27838\,
            I => \N__27835\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__27835\,
            I => \N__27832\
        );

    \I__3123\ : Span4Mux_v
    port map (
            O => \N__27832\,
            I => \N__27829\
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__27829\,
            I => \c0.n18637\
        );

    \I__3121\ : InMux
    port map (
            O => \N__27826\,
            I => \N__27817\
        );

    \I__3120\ : InMux
    port map (
            O => \N__27825\,
            I => \N__27817\
        );

    \I__3119\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27817\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__27817\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__3117\ : SRMux
    port map (
            O => \N__27814\,
            I => \N__27811\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__27811\,
            I => \N__27808\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__27808\,
            I => \c0.n18635\
        );

    \I__3114\ : InMux
    port map (
            O => \N__27805\,
            I => \N__27799\
        );

    \I__3113\ : InMux
    port map (
            O => \N__27804\,
            I => \N__27799\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__27799\,
            I => \N__27795\
        );

    \I__3111\ : InMux
    port map (
            O => \N__27798\,
            I => \N__27792\
        );

    \I__3110\ : Span4Mux_v
    port map (
            O => \N__27795\,
            I => \N__27789\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__27792\,
            I => \c0.FRAME_MATCHER_state_26\
        );

    \I__3108\ : Odrv4
    port map (
            O => \N__27789\,
            I => \c0.FRAME_MATCHER_state_26\
        );

    \I__3107\ : SRMux
    port map (
            O => \N__27784\,
            I => \N__27781\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__27781\,
            I => \N__27778\
        );

    \I__3105\ : Span4Mux_h
    port map (
            O => \N__27778\,
            I => \N__27775\
        );

    \I__3104\ : Odrv4
    port map (
            O => \N__27775\,
            I => \c0.n18623\
        );

    \I__3103\ : InMux
    port map (
            O => \N__27772\,
            I => \N__27767\
        );

    \I__3102\ : InMux
    port map (
            O => \N__27771\,
            I => \N__27764\
        );

    \I__3101\ : InMux
    port map (
            O => \N__27770\,
            I => \N__27761\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__27767\,
            I => \N__27756\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__27764\,
            I => \N__27756\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__27761\,
            I => \c0.FRAME_MATCHER_state_13\
        );

    \I__3097\ : Odrv4
    port map (
            O => \N__27756\,
            I => \c0.FRAME_MATCHER_state_13\
        );

    \I__3096\ : SRMux
    port map (
            O => \N__27751\,
            I => \N__27748\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__27748\,
            I => \N__27745\
        );

    \I__3094\ : Span4Mux_h
    port map (
            O => \N__27745\,
            I => \N__27742\
        );

    \I__3093\ : Odrv4
    port map (
            O => \N__27742\,
            I => \c0.n18665\
        );

    \I__3092\ : InMux
    port map (
            O => \N__27739\,
            I => \N__27734\
        );

    \I__3091\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27731\
        );

    \I__3090\ : InMux
    port map (
            O => \N__27737\,
            I => \N__27728\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__27734\,
            I => \N__27723\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__27731\,
            I => \N__27723\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__27728\,
            I => \c0.FRAME_MATCHER_state_23\
        );

    \I__3086\ : Odrv12
    port map (
            O => \N__27723\,
            I => \c0.FRAME_MATCHER_state_23\
        );

    \I__3085\ : InMux
    port map (
            O => \N__27718\,
            I => \N__27714\
        );

    \I__3084\ : CascadeMux
    port map (
            O => \N__27717\,
            I => \N__27711\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__27714\,
            I => \N__27707\
        );

    \I__3082\ : InMux
    port map (
            O => \N__27711\,
            I => \N__27702\
        );

    \I__3081\ : InMux
    port map (
            O => \N__27710\,
            I => \N__27702\
        );

    \I__3080\ : Odrv4
    port map (
            O => \N__27707\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__27702\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__3078\ : InMux
    port map (
            O => \N__27697\,
            I => \N__27694\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__27694\,
            I => \c0.tx.n4\
        );

    \I__3076\ : CascadeMux
    port map (
            O => \N__27691\,
            I => \c0.tx.n21179_cascade_\
        );

    \I__3075\ : InMux
    port map (
            O => \N__27688\,
            I => \N__27682\
        );

    \I__3074\ : InMux
    port map (
            O => \N__27687\,
            I => \N__27682\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__27682\,
            I => \N__27675\
        );

    \I__3072\ : InMux
    port map (
            O => \N__27681\,
            I => \N__27672\
        );

    \I__3071\ : InMux
    port map (
            O => \N__27680\,
            I => \N__27665\
        );

    \I__3070\ : InMux
    port map (
            O => \N__27679\,
            I => \N__27665\
        );

    \I__3069\ : InMux
    port map (
            O => \N__27678\,
            I => \N__27665\
        );

    \I__3068\ : Span4Mux_h
    port map (
            O => \N__27675\,
            I => \N__27662\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__27672\,
            I => \c0.r_Clock_Count_8\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__27665\,
            I => \c0.r_Clock_Count_8\
        );

    \I__3065\ : Odrv4
    port map (
            O => \N__27662\,
            I => \c0.r_Clock_Count_8\
        );

    \I__3064\ : SRMux
    port map (
            O => \N__27655\,
            I => \N__27652\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__27652\,
            I => \N__27648\
        );

    \I__3062\ : SRMux
    port map (
            O => \N__27651\,
            I => \N__27645\
        );

    \I__3061\ : Span4Mux_h
    port map (
            O => \N__27648\,
            I => \N__27642\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__27645\,
            I => \N__27639\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__27642\,
            I => \c0.tx.n12759\
        );

    \I__3058\ : Odrv4
    port map (
            O => \N__27639\,
            I => \c0.tx.n12759\
        );

    \I__3057\ : InMux
    port map (
            O => \N__27634\,
            I => \N__27629\
        );

    \I__3056\ : InMux
    port map (
            O => \N__27633\,
            I => \N__27626\
        );

    \I__3055\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27623\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__27629\,
            I => \N__27620\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__27626\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__27623\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__3051\ : Odrv12
    port map (
            O => \N__27620\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__3050\ : CascadeMux
    port map (
            O => \N__27613\,
            I => \N__27608\
        );

    \I__3049\ : InMux
    port map (
            O => \N__27612\,
            I => \N__27605\
        );

    \I__3048\ : InMux
    port map (
            O => \N__27611\,
            I => \N__27602\
        );

    \I__3047\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27599\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__27605\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__27602\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__27599\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__3043\ : InMux
    port map (
            O => \N__27592\,
            I => \N__27583\
        );

    \I__3042\ : InMux
    port map (
            O => \N__27591\,
            I => \N__27583\
        );

    \I__3041\ : InMux
    port map (
            O => \N__27590\,
            I => \N__27583\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__27583\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__3039\ : SRMux
    port map (
            O => \N__27580\,
            I => \N__27577\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__27577\,
            I => \N__27574\
        );

    \I__3037\ : Span4Mux_h
    port map (
            O => \N__27574\,
            I => \N__27571\
        );

    \I__3036\ : Odrv4
    port map (
            O => \N__27571\,
            I => \c0.n18669\
        );

    \I__3035\ : SRMux
    port map (
            O => \N__27568\,
            I => \N__27565\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__27565\,
            I => \N__27562\
        );

    \I__3033\ : Odrv4
    port map (
            O => \N__27562\,
            I => \c0.n18679\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__27559\,
            I => \c0.n21506_cascade_\
        );

    \I__3031\ : InMux
    port map (
            O => \N__27556\,
            I => \N__27552\
        );

    \I__3030\ : InMux
    port map (
            O => \N__27555\,
            I => \N__27549\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__27552\,
            I => \c0.n55\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__27549\,
            I => \c0.n55\
        );

    \I__3027\ : CascadeMux
    port map (
            O => \N__27544\,
            I => \N__27539\
        );

    \I__3026\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27536\
        );

    \I__3025\ : InMux
    port map (
            O => \N__27542\,
            I => \N__27531\
        );

    \I__3024\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27531\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__27536\,
            I => \c0.r_Bit_Index_2\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__27531\,
            I => \c0.r_Bit_Index_2\
        );

    \I__3021\ : CascadeMux
    port map (
            O => \N__27526\,
            I => \c0.n21414_cascade_\
        );

    \I__3020\ : InMux
    port map (
            O => \N__27523\,
            I => \N__27520\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__27520\,
            I => \c0.n11\
        );

    \I__3018\ : InMux
    port map (
            O => \N__27517\,
            I => \N__27511\
        );

    \I__3017\ : InMux
    port map (
            O => \N__27516\,
            I => \N__27508\
        );

    \I__3016\ : InMux
    port map (
            O => \N__27515\,
            I => \N__27503\
        );

    \I__3015\ : InMux
    port map (
            O => \N__27514\,
            I => \N__27503\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__27511\,
            I => \c0.n15938\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__27508\,
            I => \c0.n15938\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__27503\,
            I => \c0.n15938\
        );

    \I__3011\ : InMux
    port map (
            O => \N__27496\,
            I => \N__27493\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__27493\,
            I => \c0.tx.n8\
        );

    \I__3009\ : CascadeMux
    port map (
            O => \N__27490\,
            I => \c0.n55_cascade_\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__27487\,
            I => \c0.n14301_cascade_\
        );

    \I__3007\ : InMux
    port map (
            O => \N__27484\,
            I => \N__27481\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__27481\,
            I => \c0.n15942\
        );

    \I__3005\ : InMux
    port map (
            O => \N__27478\,
            I => \N__27475\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__27475\,
            I => n6866
        );

    \I__3003\ : InMux
    port map (
            O => \N__27472\,
            I => \N__27468\
        );

    \I__3002\ : InMux
    port map (
            O => \N__27471\,
            I => \N__27465\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__27468\,
            I => data_out_frame_10_4
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__27465\,
            I => data_out_frame_10_4
        );

    \I__2999\ : InMux
    port map (
            O => \N__27460\,
            I => \N__27457\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__27457\,
            I => \c0.n21288\
        );

    \I__2997\ : InMux
    port map (
            O => \N__27454\,
            I => \N__27451\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__27451\,
            I => \N__27448\
        );

    \I__2995\ : Span4Mux_v
    port map (
            O => \N__27448\,
            I => \N__27445\
        );

    \I__2994\ : Odrv4
    port map (
            O => \N__27445\,
            I => n2273
        );

    \I__2993\ : CascadeMux
    port map (
            O => \N__27442\,
            I => \N__27439\
        );

    \I__2992\ : InMux
    port map (
            O => \N__27439\,
            I => \N__27436\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__27436\,
            I => \N__27432\
        );

    \I__2990\ : InMux
    port map (
            O => \N__27435\,
            I => \N__27428\
        );

    \I__2989\ : Span4Mux_h
    port map (
            O => \N__27432\,
            I => \N__27425\
        );

    \I__2988\ : InMux
    port map (
            O => \N__27431\,
            I => \N__27422\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__27428\,
            I => \N__27417\
        );

    \I__2986\ : Span4Mux_v
    port map (
            O => \N__27425\,
            I => \N__27417\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__27422\,
            I => encoder0_position_6
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__27417\,
            I => encoder0_position_6
        );

    \I__2983\ : InMux
    port map (
            O => \N__27412\,
            I => \N__27409\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__27409\,
            I => \c0.n21517\
        );

    \I__2981\ : CascadeMux
    port map (
            O => \N__27406\,
            I => \c0.n21626_cascade_\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__27403\,
            I => \N__27399\
        );

    \I__2979\ : InMux
    port map (
            O => \N__27402\,
            I => \N__27395\
        );

    \I__2978\ : InMux
    port map (
            O => \N__27399\,
            I => \N__27392\
        );

    \I__2977\ : InMux
    port map (
            O => \N__27398\,
            I => \N__27389\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__27395\,
            I => \N__27386\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__27392\,
            I => \N__27383\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__27389\,
            I => encoder0_position_7
        );

    \I__2973\ : Odrv4
    port map (
            O => \N__27386\,
            I => encoder0_position_7
        );

    \I__2972\ : Odrv4
    port map (
            O => \N__27383\,
            I => encoder0_position_7
        );

    \I__2971\ : InMux
    port map (
            O => \N__27376\,
            I => \N__27370\
        );

    \I__2970\ : InMux
    port map (
            O => \N__27375\,
            I => \N__27370\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__27370\,
            I => data_out_frame_9_7
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__27367\,
            I => \N__27364\
        );

    \I__2967\ : InMux
    port map (
            O => \N__27364\,
            I => \N__27361\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__27361\,
            I => \c0.n11_adj_3472\
        );

    \I__2965\ : InMux
    port map (
            O => \N__27358\,
            I => \N__27355\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__27355\,
            I => \c0.n11_adj_3479\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__27352\,
            I => \c0.n11_adj_3444_cascade_\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__27349\,
            I => \c0.n21289_cascade_\
        );

    \I__2961\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27342\
        );

    \I__2960\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27339\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__27342\,
            I => \N__27336\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__27339\,
            I => data_out_frame_6_1
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__27336\,
            I => data_out_frame_6_1
        );

    \I__2956\ : InMux
    port map (
            O => \N__27331\,
            I => \N__27328\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__27328\,
            I => \N__27323\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__27327\,
            I => \N__27320\
        );

    \I__2953\ : InMux
    port map (
            O => \N__27326\,
            I => \N__27317\
        );

    \I__2952\ : Span4Mux_v
    port map (
            O => \N__27323\,
            I => \N__27314\
        );

    \I__2951\ : InMux
    port map (
            O => \N__27320\,
            I => \N__27311\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__27317\,
            I => encoder0_position_1
        );

    \I__2949\ : Odrv4
    port map (
            O => \N__27314\,
            I => encoder0_position_1
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__27311\,
            I => encoder0_position_1
        );

    \I__2947\ : InMux
    port map (
            O => \N__27304\,
            I => \N__27301\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__27301\,
            I => n2251
        );

    \I__2945\ : InMux
    port map (
            O => \N__27298\,
            I => \N__27294\
        );

    \I__2944\ : CascadeMux
    port map (
            O => \N__27297\,
            I => \N__27290\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__27294\,
            I => \N__27287\
        );

    \I__2942\ : InMux
    port map (
            O => \N__27293\,
            I => \N__27284\
        );

    \I__2941\ : InMux
    port map (
            O => \N__27290\,
            I => \N__27281\
        );

    \I__2940\ : Odrv4
    port map (
            O => \N__27287\,
            I => encoder0_position_28
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__27284\,
            I => encoder0_position_28
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__27281\,
            I => encoder0_position_28
        );

    \I__2937\ : InMux
    port map (
            O => \N__27274\,
            I => \N__27270\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__27273\,
            I => \N__27266\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__27270\,
            I => \N__27263\
        );

    \I__2934\ : InMux
    port map (
            O => \N__27269\,
            I => \N__27260\
        );

    \I__2933\ : InMux
    port map (
            O => \N__27266\,
            I => \N__27257\
        );

    \I__2932\ : Odrv4
    port map (
            O => \N__27263\,
            I => encoder0_position_16
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__27260\,
            I => encoder0_position_16
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__27257\,
            I => encoder0_position_16
        );

    \I__2929\ : InMux
    port map (
            O => \N__27250\,
            I => \N__27246\
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__27249\,
            I => \N__27242\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__27246\,
            I => \N__27239\
        );

    \I__2926\ : InMux
    port map (
            O => \N__27245\,
            I => \N__27236\
        );

    \I__2925\ : InMux
    port map (
            O => \N__27242\,
            I => \N__27233\
        );

    \I__2924\ : Odrv12
    port map (
            O => \N__27239\,
            I => encoder0_position_14
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__27236\,
            I => encoder0_position_14
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__27233\,
            I => encoder0_position_14
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__27226\,
            I => \N__27222\
        );

    \I__2920\ : InMux
    port map (
            O => \N__27225\,
            I => \N__27219\
        );

    \I__2919\ : InMux
    port map (
            O => \N__27222\,
            I => \N__27216\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__27219\,
            I => data_out_frame_8_6
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__27216\,
            I => data_out_frame_8_6
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__27211\,
            I => \N__27208\
        );

    \I__2915\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27204\
        );

    \I__2914\ : InMux
    port map (
            O => \N__27207\,
            I => \N__27200\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__27204\,
            I => \N__27197\
        );

    \I__2912\ : InMux
    port map (
            O => \N__27203\,
            I => \N__27194\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__27200\,
            I => \N__27189\
        );

    \I__2910\ : Span4Mux_h
    port map (
            O => \N__27197\,
            I => \N__27189\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__27194\,
            I => encoder0_position_4
        );

    \I__2908\ : Odrv4
    port map (
            O => \N__27189\,
            I => encoder0_position_4
        );

    \I__2907\ : InMux
    port map (
            O => \N__27184\,
            I => \N__27181\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__27181\,
            I => \c0.n21632\
        );

    \I__2905\ : InMux
    port map (
            O => \N__27178\,
            I => \N__27175\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__27175\,
            I => \N__27172\
        );

    \I__2903\ : Odrv4
    port map (
            O => \N__27172\,
            I => \c0.n21299\
        );

    \I__2902\ : InMux
    port map (
            O => \N__27169\,
            I => \N__27165\
        );

    \I__2901\ : InMux
    port map (
            O => \N__27168\,
            I => \N__27162\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__27165\,
            I => \N__27159\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__27162\,
            I => data_out_frame_8_7
        );

    \I__2898\ : Odrv4
    port map (
            O => \N__27159\,
            I => data_out_frame_8_7
        );

    \I__2897\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27150\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__27153\,
            I => \N__27146\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__27150\,
            I => \N__27143\
        );

    \I__2894\ : InMux
    port map (
            O => \N__27149\,
            I => \N__27140\
        );

    \I__2893\ : InMux
    port map (
            O => \N__27146\,
            I => \N__27137\
        );

    \I__2892\ : Odrv4
    port map (
            O => \N__27143\,
            I => encoder0_position_25
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__27140\,
            I => encoder0_position_25
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__27137\,
            I => encoder0_position_25
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__27130\,
            I => \N__27125\
        );

    \I__2888\ : InMux
    port map (
            O => \N__27129\,
            I => \N__27122\
        );

    \I__2887\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27119\
        );

    \I__2886\ : InMux
    port map (
            O => \N__27125\,
            I => \N__27116\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__27122\,
            I => encoder0_position_10
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__27119\,
            I => encoder0_position_10
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__27116\,
            I => encoder0_position_10
        );

    \I__2882\ : InMux
    port map (
            O => \N__27109\,
            I => \N__27104\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__27108\,
            I => \N__27101\
        );

    \I__2880\ : InMux
    port map (
            O => \N__27107\,
            I => \N__27098\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__27104\,
            I => \N__27095\
        );

    \I__2878\ : InMux
    port map (
            O => \N__27101\,
            I => \N__27092\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__27098\,
            I => encoder0_position_20
        );

    \I__2876\ : Odrv4
    port map (
            O => \N__27095\,
            I => encoder0_position_20
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__27092\,
            I => encoder0_position_20
        );

    \I__2874\ : InMux
    port map (
            O => \N__27085\,
            I => \N__27082\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__27082\,
            I => \N__27078\
        );

    \I__2872\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27075\
        );

    \I__2871\ : Span4Mux_h
    port map (
            O => \N__27078\,
            I => \N__27072\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__27075\,
            I => data_out_frame_7_4
        );

    \I__2869\ : Odrv4
    port map (
            O => \N__27072\,
            I => data_out_frame_7_4
        );

    \I__2868\ : InMux
    port map (
            O => \N__27067\,
            I => \N__27064\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__27064\,
            I => n2253
        );

    \I__2866\ : InMux
    port map (
            O => \N__27061\,
            I => \N__27058\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__27058\,
            I => n2249
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__27055\,
            I => \N__27052\
        );

    \I__2863\ : InMux
    port map (
            O => \N__27052\,
            I => \N__27048\
        );

    \I__2862\ : CascadeMux
    port map (
            O => \N__27051\,
            I => \N__27044\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__27048\,
            I => \N__27041\
        );

    \I__2860\ : InMux
    port map (
            O => \N__27047\,
            I => \N__27038\
        );

    \I__2859\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27035\
        );

    \I__2858\ : Odrv4
    port map (
            O => \N__27041\,
            I => encoder0_position_30
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__27038\,
            I => encoder0_position_30
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__27035\,
            I => encoder0_position_30
        );

    \I__2855\ : InMux
    port map (
            O => \N__27028\,
            I => \N__27025\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__27025\,
            I => n2267
        );

    \I__2853\ : InMux
    port map (
            O => \N__27022\,
            I => \N__27019\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__27019\,
            I => n2266
        );

    \I__2851\ : InMux
    port map (
            O => \N__27016\,
            I => \N__27013\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__27013\,
            I => n2265
        );

    \I__2849\ : InMux
    port map (
            O => \N__27010\,
            I => \N__27007\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__27007\,
            I => n2264
        );

    \I__2847\ : InMux
    port map (
            O => \N__27004\,
            I => \N__27000\
        );

    \I__2846\ : CascadeMux
    port map (
            O => \N__27003\,
            I => \N__26997\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__27000\,
            I => \N__26993\
        );

    \I__2844\ : InMux
    port map (
            O => \N__26997\,
            I => \N__26990\
        );

    \I__2843\ : InMux
    port map (
            O => \N__26996\,
            I => \N__26987\
        );

    \I__2842\ : Span12Mux_v
    port map (
            O => \N__26993\,
            I => \N__26984\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__26990\,
            I => \N__26981\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__26987\,
            I => encoder0_position_15
        );

    \I__2839\ : Odrv12
    port map (
            O => \N__26984\,
            I => encoder0_position_15
        );

    \I__2838\ : Odrv4
    port map (
            O => \N__26981\,
            I => encoder0_position_15
        );

    \I__2837\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26971\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__26971\,
            I => n2263
        );

    \I__2835\ : InMux
    port map (
            O => \N__26968\,
            I => \N__26965\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__26965\,
            I => n2262
        );

    \I__2833\ : InMux
    port map (
            O => \N__26962\,
            I => \N__26959\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__26959\,
            I => \N__26955\
        );

    \I__2831\ : InMux
    port map (
            O => \N__26958\,
            I => \N__26952\
        );

    \I__2830\ : Span4Mux_h
    port map (
            O => \N__26955\,
            I => \N__26949\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__26952\,
            I => data_out_frame_6_4
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__26949\,
            I => data_out_frame_6_4
        );

    \I__2827\ : CascadeMux
    port map (
            O => \N__26944\,
            I => \quad_counter1.n16_cascade_\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__26941\,
            I => \quad_counter1.n24_adj_3578_cascade_\
        );

    \I__2825\ : InMux
    port map (
            O => \N__26938\,
            I => \N__26932\
        );

    \I__2824\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26932\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__26932\,
            I => n11351
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__26929\,
            I => \N__26924\
        );

    \I__2821\ : InMux
    port map (
            O => \N__26928\,
            I => \N__26919\
        );

    \I__2820\ : InMux
    port map (
            O => \N__26927\,
            I => \N__26919\
        );

    \I__2819\ : InMux
    port map (
            O => \N__26924\,
            I => \N__26916\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__26919\,
            I => \N__26911\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__26916\,
            I => \N__26911\
        );

    \I__2816\ : Odrv4
    port map (
            O => \N__26911\,
            I => \B_filtered\
        );

    \I__2815\ : InMux
    port map (
            O => \N__26908\,
            I => \N__26905\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__26905\,
            I => \N__26900\
        );

    \I__2813\ : InMux
    port map (
            O => \N__26904\,
            I => \N__26895\
        );

    \I__2812\ : InMux
    port map (
            O => \N__26903\,
            I => \N__26895\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__26900\,
            I => \quad_counter0.B_delayed\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__26895\,
            I => \quad_counter0.B_delayed\
        );

    \I__2809\ : InMux
    port map (
            O => \N__26890\,
            I => \N__26887\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__26887\,
            I => \quad_counter1.n6\
        );

    \I__2807\ : InMux
    port map (
            O => \N__26884\,
            I => \N__26875\
        );

    \I__2806\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26875\
        );

    \I__2805\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26870\
        );

    \I__2804\ : InMux
    port map (
            O => \N__26881\,
            I => \N__26870\
        );

    \I__2803\ : InMux
    port map (
            O => \N__26880\,
            I => \N__26867\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__26875\,
            I => \N__26864\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__26870\,
            I => \N__26861\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__26867\,
            I => \A_filtered\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__26864\,
            I => \A_filtered\
        );

    \I__2798\ : Odrv4
    port map (
            O => \N__26861\,
            I => \A_filtered\
        );

    \I__2797\ : InMux
    port map (
            O => \N__26854\,
            I => \N__26851\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__26851\,
            I => \quad_counter0.A_delayed\
        );

    \I__2795\ : InMux
    port map (
            O => \N__26848\,
            I => \N__26845\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__26845\,
            I => \quad_counter1.n22\
        );

    \I__2793\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26839\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__26839\,
            I => n2269
        );

    \I__2791\ : InMux
    port map (
            O => \N__26836\,
            I => \N__26833\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__26833\,
            I => n2268
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__26830\,
            I => \n11343_cascade_\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__26827\,
            I => \n12417_cascade_\
        );

    \I__2787\ : InMux
    port map (
            O => \N__26824\,
            I => \N__26821\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__26821\,
            I => \quad_counter1.n28_adj_3574\
        );

    \I__2785\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26810\
        );

    \I__2784\ : InMux
    port map (
            O => \N__26817\,
            I => \N__26810\
        );

    \I__2783\ : InMux
    port map (
            O => \N__26816\,
            I => \N__26805\
        );

    \I__2782\ : InMux
    port map (
            O => \N__26815\,
            I => \N__26805\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__26810\,
            I => \N__26800\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__26805\,
            I => \N__26800\
        );

    \I__2779\ : Span4Mux_v
    port map (
            O => \N__26800\,
            I => \N__26797\
        );

    \I__2778\ : Sp12to4
    port map (
            O => \N__26797\,
            I => \N__26794\
        );

    \I__2777\ : Odrv12
    port map (
            O => \N__26794\,
            I => \PIN_13_c\
        );

    \I__2776\ : CascadeMux
    port map (
            O => \N__26791\,
            I => \N__26788\
        );

    \I__2775\ : InMux
    port map (
            O => \N__26788\,
            I => \N__26785\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__26785\,
            I => n11343
        );

    \I__2773\ : InMux
    port map (
            O => \N__26782\,
            I => \N__26775\
        );

    \I__2772\ : InMux
    port map (
            O => \N__26781\,
            I => \N__26775\
        );

    \I__2771\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26772\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__26775\,
            I => \quadB_delayed_adj_3585\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__26772\,
            I => \quadB_delayed_adj_3585\
        );

    \I__2768\ : InMux
    port map (
            O => \N__26767\,
            I => \N__26764\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__26764\,
            I => \quad_counter1.n26_adj_3575\
        );

    \I__2766\ : InMux
    port map (
            O => \N__26761\,
            I => \N__26758\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__26758\,
            I => \quad_counter1.n27_adj_3576\
        );

    \I__2764\ : SRMux
    port map (
            O => \N__26755\,
            I => \N__26752\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__26752\,
            I => \N__26749\
        );

    \I__2762\ : Odrv4
    port map (
            O => \N__26749\,
            I => \c0.n18671\
        );

    \I__2761\ : SRMux
    port map (
            O => \N__26746\,
            I => \N__26743\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__26743\,
            I => \N__26740\
        );

    \I__2759\ : Span4Mux_h
    port map (
            O => \N__26740\,
            I => \N__26737\
        );

    \I__2758\ : Odrv4
    port map (
            O => \N__26737\,
            I => \c0.n18617\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__26734\,
            I => \quad_counter1.n25_adj_3577_cascade_\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__26731\,
            I => \N__26727\
        );

    \I__2755\ : InMux
    port map (
            O => \N__26730\,
            I => \N__26724\
        );

    \I__2754\ : InMux
    port map (
            O => \N__26727\,
            I => \N__26721\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__26724\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__26721\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__2751\ : InMux
    port map (
            O => \N__26716\,
            I => \c0.tx.n17274\
        );

    \I__2750\ : InMux
    port map (
            O => \N__26713\,
            I => \N__26709\
        );

    \I__2749\ : InMux
    port map (
            O => \N__26712\,
            I => \N__26706\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__26709\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__26706\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__2746\ : InMux
    port map (
            O => \N__26701\,
            I => \c0.tx.n17275\
        );

    \I__2745\ : InMux
    port map (
            O => \N__26698\,
            I => \N__26694\
        );

    \I__2744\ : InMux
    port map (
            O => \N__26697\,
            I => \N__26691\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__26694\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__26691\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__2741\ : InMux
    port map (
            O => \N__26686\,
            I => \c0.tx.n17276\
        );

    \I__2740\ : InMux
    port map (
            O => \N__26683\,
            I => \N__26679\
        );

    \I__2739\ : InMux
    port map (
            O => \N__26682\,
            I => \N__26676\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__26679\,
            I => \c0.tx.r_Clock_Count_4\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__26676\,
            I => \c0.tx.r_Clock_Count_4\
        );

    \I__2736\ : InMux
    port map (
            O => \N__26671\,
            I => \c0.tx.n17277\
        );

    \I__2735\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26664\
        );

    \I__2734\ : InMux
    port map (
            O => \N__26667\,
            I => \N__26661\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__26664\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__26661\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__2731\ : InMux
    port map (
            O => \N__26656\,
            I => \c0.tx.n17278\
        );

    \I__2730\ : InMux
    port map (
            O => \N__26653\,
            I => \N__26649\
        );

    \I__2729\ : InMux
    port map (
            O => \N__26652\,
            I => \N__26646\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__26649\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__26646\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__2726\ : InMux
    port map (
            O => \N__26641\,
            I => \c0.tx.n17279\
        );

    \I__2725\ : InMux
    port map (
            O => \N__26638\,
            I => \N__26634\
        );

    \I__2724\ : InMux
    port map (
            O => \N__26637\,
            I => \N__26631\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__26634\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__26631\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__2721\ : InMux
    port map (
            O => \N__26626\,
            I => \c0.tx.n17280\
        );

    \I__2720\ : InMux
    port map (
            O => \N__26623\,
            I => \bfn_10_19_0_\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__26620\,
            I => \N__26617\
        );

    \I__2718\ : InMux
    port map (
            O => \N__26617\,
            I => \N__26596\
        );

    \I__2717\ : InMux
    port map (
            O => \N__26616\,
            I => \N__26596\
        );

    \I__2716\ : InMux
    port map (
            O => \N__26615\,
            I => \N__26596\
        );

    \I__2715\ : InMux
    port map (
            O => \N__26614\,
            I => \N__26591\
        );

    \I__2714\ : InMux
    port map (
            O => \N__26613\,
            I => \N__26588\
        );

    \I__2713\ : InMux
    port map (
            O => \N__26612\,
            I => \N__26581\
        );

    \I__2712\ : InMux
    port map (
            O => \N__26611\,
            I => \N__26581\
        );

    \I__2711\ : InMux
    port map (
            O => \N__26610\,
            I => \N__26581\
        );

    \I__2710\ : InMux
    port map (
            O => \N__26609\,
            I => \N__26578\
        );

    \I__2709\ : InMux
    port map (
            O => \N__26608\,
            I => \N__26565\
        );

    \I__2708\ : InMux
    port map (
            O => \N__26607\,
            I => \N__26565\
        );

    \I__2707\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26565\
        );

    \I__2706\ : InMux
    port map (
            O => \N__26605\,
            I => \N__26565\
        );

    \I__2705\ : InMux
    port map (
            O => \N__26604\,
            I => \N__26565\
        );

    \I__2704\ : InMux
    port map (
            O => \N__26603\,
            I => \N__26565\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__26596\,
            I => \N__26562\
        );

    \I__2702\ : InMux
    port map (
            O => \N__26595\,
            I => \N__26559\
        );

    \I__2701\ : InMux
    port map (
            O => \N__26594\,
            I => \N__26556\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__26591\,
            I => \N__26551\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__26588\,
            I => \N__26551\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__26581\,
            I => \N__26548\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__26578\,
            I => \N__26543\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__26565\,
            I => \N__26543\
        );

    \I__2695\ : Span4Mux_h
    port map (
            O => \N__26562\,
            I => \N__26536\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__26559\,
            I => \N__26536\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__26556\,
            I => \N__26533\
        );

    \I__2692\ : Sp12to4
    port map (
            O => \N__26551\,
            I => \N__26530\
        );

    \I__2691\ : Span4Mux_v
    port map (
            O => \N__26548\,
            I => \N__26527\
        );

    \I__2690\ : Sp12to4
    port map (
            O => \N__26543\,
            I => \N__26524\
        );

    \I__2689\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26519\
        );

    \I__2688\ : InMux
    port map (
            O => \N__26541\,
            I => \N__26519\
        );

    \I__2687\ : Span4Mux_h
    port map (
            O => \N__26536\,
            I => \N__26516\
        );

    \I__2686\ : Span4Mux_v
    port map (
            O => \N__26533\,
            I => \N__26513\
        );

    \I__2685\ : Span12Mux_v
    port map (
            O => \N__26530\,
            I => \N__26504\
        );

    \I__2684\ : Sp12to4
    port map (
            O => \N__26527\,
            I => \N__26504\
        );

    \I__2683\ : Span12Mux_v
    port map (
            O => \N__26524\,
            I => \N__26504\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__26519\,
            I => \N__26504\
        );

    \I__2681\ : Span4Mux_v
    port map (
            O => \N__26516\,
            I => \N__26499\
        );

    \I__2680\ : Span4Mux_h
    port map (
            O => \N__26513\,
            I => \N__26499\
        );

    \I__2679\ : Odrv12
    port map (
            O => \N__26504\,
            I => \PIN_8_c\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__26499\,
            I => \PIN_8_c\
        );

    \I__2677\ : CascadeMux
    port map (
            O => \N__26494\,
            I => \N__26479\
        );

    \I__2676\ : InMux
    port map (
            O => \N__26493\,
            I => \N__26475\
        );

    \I__2675\ : InMux
    port map (
            O => \N__26492\,
            I => \N__26466\
        );

    \I__2674\ : InMux
    port map (
            O => \N__26491\,
            I => \N__26466\
        );

    \I__2673\ : InMux
    port map (
            O => \N__26490\,
            I => \N__26453\
        );

    \I__2672\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26453\
        );

    \I__2671\ : InMux
    port map (
            O => \N__26488\,
            I => \N__26453\
        );

    \I__2670\ : InMux
    port map (
            O => \N__26487\,
            I => \N__26453\
        );

    \I__2669\ : InMux
    port map (
            O => \N__26486\,
            I => \N__26453\
        );

    \I__2668\ : InMux
    port map (
            O => \N__26485\,
            I => \N__26453\
        );

    \I__2667\ : InMux
    port map (
            O => \N__26484\,
            I => \N__26446\
        );

    \I__2666\ : InMux
    port map (
            O => \N__26483\,
            I => \N__26446\
        );

    \I__2665\ : InMux
    port map (
            O => \N__26482\,
            I => \N__26446\
        );

    \I__2664\ : InMux
    port map (
            O => \N__26479\,
            I => \N__26443\
        );

    \I__2663\ : InMux
    port map (
            O => \N__26478\,
            I => \N__26440\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__26475\,
            I => \N__26437\
        );

    \I__2661\ : InMux
    port map (
            O => \N__26474\,
            I => \N__26430\
        );

    \I__2660\ : InMux
    port map (
            O => \N__26473\,
            I => \N__26430\
        );

    \I__2659\ : InMux
    port map (
            O => \N__26472\,
            I => \N__26430\
        );

    \I__2658\ : InMux
    port map (
            O => \N__26471\,
            I => \N__26427\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__26466\,
            I => \N__26424\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__26453\,
            I => \N__26419\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__26446\,
            I => \N__26419\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__26443\,
            I => \N__26416\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__26440\,
            I => \N__26411\
        );

    \I__2652\ : Span4Mux_h
    port map (
            O => \N__26437\,
            I => \N__26411\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__26430\,
            I => \N__26408\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__26427\,
            I => \N__26405\
        );

    \I__2649\ : Span4Mux_v
    port map (
            O => \N__26424\,
            I => \N__26400\
        );

    \I__2648\ : Span4Mux_v
    port map (
            O => \N__26419\,
            I => \N__26400\
        );

    \I__2647\ : Span12Mux_h
    port map (
            O => \N__26416\,
            I => \N__26397\
        );

    \I__2646\ : Span4Mux_v
    port map (
            O => \N__26411\,
            I => \N__26392\
        );

    \I__2645\ : Span4Mux_h
    port map (
            O => \N__26408\,
            I => \N__26392\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__26405\,
            I => \quadB_delayed\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__26400\,
            I => \quadB_delayed\
        );

    \I__2642\ : Odrv12
    port map (
            O => \N__26397\,
            I => \quadB_delayed\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__26392\,
            I => \quadB_delayed\
        );

    \I__2640\ : InMux
    port map (
            O => \N__26383\,
            I => \N__26380\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__26380\,
            I => \N__26377\
        );

    \I__2638\ : Odrv4
    port map (
            O => \N__26377\,
            I => \quad_counter0.n13187\
        );

    \I__2637\ : InMux
    port map (
            O => \N__26374\,
            I => \N__26370\
        );

    \I__2636\ : InMux
    port map (
            O => \N__26373\,
            I => \N__26367\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__26370\,
            I => \N__26361\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__26367\,
            I => \N__26361\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__26366\,
            I => \N__26358\
        );

    \I__2632\ : Span4Mux_h
    port map (
            O => \N__26361\,
            I => \N__26355\
        );

    \I__2631\ : InMux
    port map (
            O => \N__26358\,
            I => \N__26352\
        );

    \I__2630\ : Odrv4
    port map (
            O => \N__26355\,
            I => \quad_counter0.b_delay_counter_2\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__26352\,
            I => \quad_counter0.b_delay_counter_2\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__26347\,
            I => \c0.n21331_cascade_\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__26344\,
            I => \c0.n17354_cascade_\
        );

    \I__2626\ : InMux
    port map (
            O => \N__26341\,
            I => \N__26338\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__26338\,
            I => \c0.n21521\
        );

    \I__2624\ : CascadeMux
    port map (
            O => \N__26335\,
            I => \c0.tx.n6_cascade_\
        );

    \I__2623\ : CascadeMux
    port map (
            O => \N__26332\,
            I => \c0.n15938_cascade_\
        );

    \I__2622\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26326\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__26326\,
            I => \c0.tx.r_Clock_Count_0\
        );

    \I__2620\ : InMux
    port map (
            O => \N__26323\,
            I => \bfn_10_18_0_\
        );

    \I__2619\ : InMux
    port map (
            O => \N__26320\,
            I => \N__26317\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__26317\,
            I => \quad_counter0.n13269\
        );

    \I__2617\ : InMux
    port map (
            O => \N__26314\,
            I => \N__26309\
        );

    \I__2616\ : InMux
    port map (
            O => \N__26313\,
            I => \N__26306\
        );

    \I__2615\ : InMux
    port map (
            O => \N__26312\,
            I => \N__26303\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__26309\,
            I => \N__26300\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__26306\,
            I => \N__26295\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__26303\,
            I => \N__26295\
        );

    \I__2611\ : Odrv12
    port map (
            O => \N__26300\,
            I => \quad_counter0.b_delay_counter_15\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__26295\,
            I => \quad_counter0.b_delay_counter_15\
        );

    \I__2609\ : InMux
    port map (
            O => \N__26290\,
            I => \N__26287\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__26287\,
            I => \N__26284\
        );

    \I__2607\ : Odrv4
    port map (
            O => \N__26284\,
            I => \quad_counter0.n26_adj_2991\
        );

    \I__2606\ : InMux
    port map (
            O => \N__26281\,
            I => \N__26278\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__26278\,
            I => \N__26275\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__26275\,
            I => \quad_counter0.n27_adj_2992\
        );

    \I__2603\ : CascadeMux
    port map (
            O => \N__26272\,
            I => \N__26269\
        );

    \I__2602\ : InMux
    port map (
            O => \N__26269\,
            I => \N__26266\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__26266\,
            I => \quad_counter0.n28_adj_2990\
        );

    \I__2600\ : InMux
    port map (
            O => \N__26263\,
            I => \N__26260\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__26260\,
            I => \quad_counter0.n25_adj_2993\
        );

    \I__2598\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26254\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__26254\,
            I => \N__26251\
        );

    \I__2596\ : Span12Mux_v
    port map (
            O => \N__26251\,
            I => \N__26248\
        );

    \I__2595\ : Odrv12
    port map (
            O => \N__26248\,
            I => n11347
        );

    \I__2594\ : CascadeMux
    port map (
            O => \N__26245\,
            I => \n11347_cascade_\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__26242\,
            I => \N__26224\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__26241\,
            I => \N__26221\
        );

    \I__2591\ : CascadeMux
    port map (
            O => \N__26240\,
            I => \N__26218\
        );

    \I__2590\ : CascadeMux
    port map (
            O => \N__26239\,
            I => \N__26215\
        );

    \I__2589\ : CascadeMux
    port map (
            O => \N__26238\,
            I => \N__26212\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__26237\,
            I => \N__26209\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__26236\,
            I => \N__26206\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__26235\,
            I => \N__26203\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__26234\,
            I => \N__26200\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__26233\,
            I => \N__26197\
        );

    \I__2583\ : CascadeMux
    port map (
            O => \N__26232\,
            I => \N__26194\
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__26231\,
            I => \N__26191\
        );

    \I__2581\ : CascadeMux
    port map (
            O => \N__26230\,
            I => \N__26188\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__26229\,
            I => \N__26185\
        );

    \I__2579\ : CascadeMux
    port map (
            O => \N__26228\,
            I => \N__26182\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__26227\,
            I => \N__26179\
        );

    \I__2577\ : InMux
    port map (
            O => \N__26224\,
            I => \N__26170\
        );

    \I__2576\ : InMux
    port map (
            O => \N__26221\,
            I => \N__26170\
        );

    \I__2575\ : InMux
    port map (
            O => \N__26218\,
            I => \N__26170\
        );

    \I__2574\ : InMux
    port map (
            O => \N__26215\,
            I => \N__26170\
        );

    \I__2573\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26161\
        );

    \I__2572\ : InMux
    port map (
            O => \N__26209\,
            I => \N__26161\
        );

    \I__2571\ : InMux
    port map (
            O => \N__26206\,
            I => \N__26161\
        );

    \I__2570\ : InMux
    port map (
            O => \N__26203\,
            I => \N__26161\
        );

    \I__2569\ : InMux
    port map (
            O => \N__26200\,
            I => \N__26152\
        );

    \I__2568\ : InMux
    port map (
            O => \N__26197\,
            I => \N__26152\
        );

    \I__2567\ : InMux
    port map (
            O => \N__26194\,
            I => \N__26152\
        );

    \I__2566\ : InMux
    port map (
            O => \N__26191\,
            I => \N__26152\
        );

    \I__2565\ : InMux
    port map (
            O => \N__26188\,
            I => \N__26143\
        );

    \I__2564\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26143\
        );

    \I__2563\ : InMux
    port map (
            O => \N__26182\,
            I => \N__26143\
        );

    \I__2562\ : InMux
    port map (
            O => \N__26179\,
            I => \N__26143\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__26170\,
            I => \quad_counter0.n21603\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__26161\,
            I => \quad_counter0.n21603\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__26152\,
            I => \quad_counter0.n21603\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__26143\,
            I => \quad_counter0.n21603\
        );

    \I__2557\ : InMux
    port map (
            O => \N__26134\,
            I => \N__26128\
        );

    \I__2556\ : InMux
    port map (
            O => \N__26133\,
            I => \N__26128\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__26128\,
            I => data_out_frame_10_6
        );

    \I__2554\ : InMux
    port map (
            O => \N__26125\,
            I => \N__26122\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__26122\,
            I => \c0.n21629\
        );

    \I__2552\ : InMux
    port map (
            O => \N__26119\,
            I => \N__26116\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__26116\,
            I => \N__26113\
        );

    \I__2550\ : Span4Mux_v
    port map (
            O => \N__26113\,
            I => \N__26110\
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__26110\,
            I => n2275
        );

    \I__2548\ : InMux
    port map (
            O => \N__26107\,
            I => \N__26104\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__26104\,
            I => \N__26101\
        );

    \I__2546\ : Odrv12
    port map (
            O => \N__26101\,
            I => n2272
        );

    \I__2545\ : InMux
    port map (
            O => \N__26098\,
            I => \N__26095\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__26095\,
            I => \N__26092\
        );

    \I__2543\ : Odrv12
    port map (
            O => \N__26092\,
            I => n2274
        );

    \I__2542\ : InMux
    port map (
            O => \N__26089\,
            I => \N__26086\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__26086\,
            I => n2248
        );

    \I__2540\ : InMux
    port map (
            O => \N__26083\,
            I => \N__26080\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__26080\,
            I => \N__26077\
        );

    \I__2538\ : Odrv4
    port map (
            O => \N__26077\,
            I => \c0.n5_adj_3471\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__26074\,
            I => \N__26070\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__26073\,
            I => \N__26066\
        );

    \I__2535\ : InMux
    port map (
            O => \N__26070\,
            I => \N__26063\
        );

    \I__2534\ : InMux
    port map (
            O => \N__26069\,
            I => \N__26060\
        );

    \I__2533\ : InMux
    port map (
            O => \N__26066\,
            I => \N__26057\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__26063\,
            I => \N__26054\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__26060\,
            I => encoder0_position_5
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__26057\,
            I => encoder0_position_5
        );

    \I__2529\ : Odrv12
    port map (
            O => \N__26054\,
            I => encoder0_position_5
        );

    \I__2528\ : InMux
    port map (
            O => \N__26047\,
            I => \N__26041\
        );

    \I__2527\ : InMux
    port map (
            O => \N__26046\,
            I => \N__26041\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__26041\,
            I => data_out_frame_9_6
        );

    \I__2525\ : InMux
    port map (
            O => \N__26038\,
            I => \N__26035\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__26035\,
            I => \quad_counter0.n13254\
        );

    \I__2523\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26027\
        );

    \I__2522\ : InMux
    port map (
            O => \N__26031\,
            I => \N__26024\
        );

    \I__2521\ : InMux
    port map (
            O => \N__26030\,
            I => \N__26021\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__26027\,
            I => \N__26018\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__26024\,
            I => \quad_counter0.b_delay_counter_10\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__26021\,
            I => \quad_counter0.b_delay_counter_10\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__26018\,
            I => \quad_counter0.b_delay_counter_10\
        );

    \I__2516\ : InMux
    port map (
            O => \N__26011\,
            I => \N__26008\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__26008\,
            I => n2255
        );

    \I__2514\ : InMux
    port map (
            O => \N__26005\,
            I => \quad_counter0.n17306\
        );

    \I__2513\ : InMux
    port map (
            O => \N__26002\,
            I => \N__25999\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__25999\,
            I => n2254
        );

    \I__2511\ : InMux
    port map (
            O => \N__25996\,
            I => \quad_counter0.n17307\
        );

    \I__2510\ : InMux
    port map (
            O => \N__25993\,
            I => \quad_counter0.n17308\
        );

    \I__2509\ : InMux
    port map (
            O => \N__25990\,
            I => \quad_counter0.n17309\
        );

    \I__2508\ : InMux
    port map (
            O => \N__25987\,
            I => \quad_counter0.n17310\
        );

    \I__2507\ : InMux
    port map (
            O => \N__25984\,
            I => \quad_counter0.n17311\
        );

    \I__2506\ : InMux
    port map (
            O => \N__25981\,
            I => \quad_counter0.n17312\
        );

    \I__2505\ : InMux
    port map (
            O => \N__25978\,
            I => \N__25974\
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__25977\,
            I => \N__25960\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__25974\,
            I => \N__25951\
        );

    \I__2502\ : InMux
    port map (
            O => \N__25973\,
            I => \N__25942\
        );

    \I__2501\ : InMux
    port map (
            O => \N__25972\,
            I => \N__25942\
        );

    \I__2500\ : InMux
    port map (
            O => \N__25971\,
            I => \N__25942\
        );

    \I__2499\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25942\
        );

    \I__2498\ : InMux
    port map (
            O => \N__25969\,
            I => \N__25933\
        );

    \I__2497\ : InMux
    port map (
            O => \N__25968\,
            I => \N__25933\
        );

    \I__2496\ : InMux
    port map (
            O => \N__25967\,
            I => \N__25933\
        );

    \I__2495\ : InMux
    port map (
            O => \N__25966\,
            I => \N__25933\
        );

    \I__2494\ : InMux
    port map (
            O => \N__25965\,
            I => \N__25922\
        );

    \I__2493\ : InMux
    port map (
            O => \N__25964\,
            I => \N__25922\
        );

    \I__2492\ : InMux
    port map (
            O => \N__25963\,
            I => \N__25922\
        );

    \I__2491\ : InMux
    port map (
            O => \N__25960\,
            I => \N__25922\
        );

    \I__2490\ : InMux
    port map (
            O => \N__25959\,
            I => \N__25922\
        );

    \I__2489\ : InMux
    port map (
            O => \N__25958\,
            I => \N__25915\
        );

    \I__2488\ : InMux
    port map (
            O => \N__25957\,
            I => \N__25915\
        );

    \I__2487\ : InMux
    port map (
            O => \N__25956\,
            I => \N__25915\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__25955\,
            I => \N__25902\
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__25954\,
            I => \N__25897\
        );

    \I__2484\ : Span4Mux_v
    port map (
            O => \N__25951\,
            I => \N__25884\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__25942\,
            I => \N__25884\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__25933\,
            I => \N__25884\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__25922\,
            I => \N__25884\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__25915\,
            I => \N__25884\
        );

    \I__2479\ : InMux
    port map (
            O => \N__25914\,
            I => \N__25875\
        );

    \I__2478\ : InMux
    port map (
            O => \N__25913\,
            I => \N__25875\
        );

    \I__2477\ : InMux
    port map (
            O => \N__25912\,
            I => \N__25875\
        );

    \I__2476\ : InMux
    port map (
            O => \N__25911\,
            I => \N__25875\
        );

    \I__2475\ : InMux
    port map (
            O => \N__25910\,
            I => \N__25866\
        );

    \I__2474\ : InMux
    port map (
            O => \N__25909\,
            I => \N__25866\
        );

    \I__2473\ : InMux
    port map (
            O => \N__25908\,
            I => \N__25866\
        );

    \I__2472\ : InMux
    port map (
            O => \N__25907\,
            I => \N__25866\
        );

    \I__2471\ : InMux
    port map (
            O => \N__25906\,
            I => \N__25859\
        );

    \I__2470\ : InMux
    port map (
            O => \N__25905\,
            I => \N__25859\
        );

    \I__2469\ : InMux
    port map (
            O => \N__25902\,
            I => \N__25859\
        );

    \I__2468\ : InMux
    port map (
            O => \N__25901\,
            I => \N__25848\
        );

    \I__2467\ : InMux
    port map (
            O => \N__25900\,
            I => \N__25848\
        );

    \I__2466\ : InMux
    port map (
            O => \N__25897\,
            I => \N__25848\
        );

    \I__2465\ : InMux
    port map (
            O => \N__25896\,
            I => \N__25848\
        );

    \I__2464\ : InMux
    port map (
            O => \N__25895\,
            I => \N__25848\
        );

    \I__2463\ : Odrv4
    port map (
            O => \N__25884\,
            I => \quad_counter0.n2228\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__25875\,
            I => \quad_counter0.n2228\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__25866\,
            I => \quad_counter0.n2228\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__25859\,
            I => \quad_counter0.n2228\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__25848\,
            I => \quad_counter0.n2228\
        );

    \I__2458\ : InMux
    port map (
            O => \N__25837\,
            I => \bfn_10_13_0_\
        );

    \I__2457\ : InMux
    port map (
            O => \N__25834\,
            I => \quad_counter0.n17298\
        );

    \I__2456\ : InMux
    port map (
            O => \N__25831\,
            I => \quad_counter0.n17299\
        );

    \I__2455\ : InMux
    port map (
            O => \N__25828\,
            I => \N__25825\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__25825\,
            I => n2261
        );

    \I__2453\ : InMux
    port map (
            O => \N__25822\,
            I => \quad_counter0.n17300\
        );

    \I__2452\ : InMux
    port map (
            O => \N__25819\,
            I => \N__25816\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__25816\,
            I => n2260
        );

    \I__2450\ : InMux
    port map (
            O => \N__25813\,
            I => \quad_counter0.n17301\
        );

    \I__2449\ : InMux
    port map (
            O => \N__25810\,
            I => \N__25807\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__25807\,
            I => n2259
        );

    \I__2447\ : InMux
    port map (
            O => \N__25804\,
            I => \quad_counter0.n17302\
        );

    \I__2446\ : InMux
    port map (
            O => \N__25801\,
            I => \N__25798\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__25798\,
            I => n2258
        );

    \I__2444\ : InMux
    port map (
            O => \N__25795\,
            I => \quad_counter0.n17303\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__25792\,
            I => \N__25787\
        );

    \I__2442\ : InMux
    port map (
            O => \N__25791\,
            I => \N__25784\
        );

    \I__2441\ : InMux
    port map (
            O => \N__25790\,
            I => \N__25781\
        );

    \I__2440\ : InMux
    port map (
            O => \N__25787\,
            I => \N__25778\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__25784\,
            I => encoder0_position_22
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__25781\,
            I => encoder0_position_22
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__25778\,
            I => encoder0_position_22
        );

    \I__2436\ : InMux
    port map (
            O => \N__25771\,
            I => \N__25768\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__25768\,
            I => n2257
        );

    \I__2434\ : InMux
    port map (
            O => \N__25765\,
            I => \quad_counter0.n17304\
        );

    \I__2433\ : InMux
    port map (
            O => \N__25762\,
            I => \N__25759\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__25759\,
            I => n2256
        );

    \I__2431\ : InMux
    port map (
            O => \N__25756\,
            I => \bfn_10_12_0_\
        );

    \I__2430\ : InMux
    port map (
            O => \N__25753\,
            I => \bfn_10_10_0_\
        );

    \I__2429\ : InMux
    port map (
            O => \N__25750\,
            I => \quad_counter0.n17290\
        );

    \I__2428\ : InMux
    port map (
            O => \N__25747\,
            I => \quad_counter0.n17291\
        );

    \I__2427\ : InMux
    port map (
            O => \N__25744\,
            I => \quad_counter0.n17292\
        );

    \I__2426\ : InMux
    port map (
            O => \N__25741\,
            I => \quad_counter0.n17293\
        );

    \I__2425\ : InMux
    port map (
            O => \N__25738\,
            I => \quad_counter0.n17294\
        );

    \I__2424\ : InMux
    port map (
            O => \N__25735\,
            I => \quad_counter0.n17295\
        );

    \I__2423\ : InMux
    port map (
            O => \N__25732\,
            I => \quad_counter0.n17296\
        );

    \I__2422\ : InMux
    port map (
            O => \N__25729\,
            I => \bfn_10_11_0_\
        );

    \I__2421\ : InMux
    port map (
            O => \N__25726\,
            I => \N__25723\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__25723\,
            I => \quad_counter0.count_direction\
        );

    \I__2419\ : InMux
    port map (
            O => \N__25720\,
            I => \N__25717\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__25717\,
            I => \N__25714\
        );

    \I__2417\ : Odrv12
    port map (
            O => \N__25714\,
            I => n2279
        );

    \I__2416\ : InMux
    port map (
            O => \N__25711\,
            I => \quad_counter0.n17282\
        );

    \I__2415\ : InMux
    port map (
            O => \N__25708\,
            I => \N__25705\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__25705\,
            I => n2278
        );

    \I__2413\ : InMux
    port map (
            O => \N__25702\,
            I => \quad_counter0.n17283\
        );

    \I__2412\ : InMux
    port map (
            O => \N__25699\,
            I => \N__25694\
        );

    \I__2411\ : InMux
    port map (
            O => \N__25698\,
            I => \N__25691\
        );

    \I__2410\ : InMux
    port map (
            O => \N__25697\,
            I => \N__25688\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__25694\,
            I => encoder0_position_2
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__25691\,
            I => encoder0_position_2
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__25688\,
            I => encoder0_position_2
        );

    \I__2406\ : InMux
    port map (
            O => \N__25681\,
            I => \N__25678\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__25678\,
            I => n2277
        );

    \I__2404\ : InMux
    port map (
            O => \N__25675\,
            I => \quad_counter0.n17284\
        );

    \I__2403\ : InMux
    port map (
            O => \N__25672\,
            I => \N__25668\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__25671\,
            I => \N__25665\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__25668\,
            I => \N__25662\
        );

    \I__2400\ : InMux
    port map (
            O => \N__25665\,
            I => \N__25658\
        );

    \I__2399\ : Span4Mux_v
    port map (
            O => \N__25662\,
            I => \N__25655\
        );

    \I__2398\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25652\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__25658\,
            I => \N__25649\
        );

    \I__2396\ : Odrv4
    port map (
            O => \N__25655\,
            I => encoder0_position_3
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__25652\,
            I => encoder0_position_3
        );

    \I__2394\ : Odrv4
    port map (
            O => \N__25649\,
            I => encoder0_position_3
        );

    \I__2393\ : InMux
    port map (
            O => \N__25642\,
            I => \N__25639\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__25639\,
            I => n2276
        );

    \I__2391\ : InMux
    port map (
            O => \N__25636\,
            I => \quad_counter0.n17285\
        );

    \I__2390\ : InMux
    port map (
            O => \N__25633\,
            I => \quad_counter0.n17286\
        );

    \I__2389\ : InMux
    port map (
            O => \N__25630\,
            I => \quad_counter0.n17287\
        );

    \I__2388\ : InMux
    port map (
            O => \N__25627\,
            I => \quad_counter0.n17288\
        );

    \I__2387\ : CEMux
    port map (
            O => \N__25624\,
            I => \N__25621\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__25621\,
            I => \N__25618\
        );

    \I__2385\ : Span4Mux_v
    port map (
            O => \N__25618\,
            I => \N__25613\
        );

    \I__2384\ : CEMux
    port map (
            O => \N__25617\,
            I => \N__25610\
        );

    \I__2383\ : InMux
    port map (
            O => \N__25616\,
            I => \N__25607\
        );

    \I__2382\ : Odrv4
    port map (
            O => \N__25613\,
            I => n12447
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__25610\,
            I => n12447
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__25607\,
            I => n12447
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__25600\,
            I => \N__25595\
        );

    \I__2378\ : InMux
    port map (
            O => \N__25599\,
            I => \N__25585\
        );

    \I__2377\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25585\
        );

    \I__2376\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25585\
        );

    \I__2375\ : InMux
    port map (
            O => \N__25594\,
            I => \N__25585\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__25585\,
            I => \N__25582\
        );

    \I__2373\ : Span4Mux_v
    port map (
            O => \N__25582\,
            I => \N__25579\
        );

    \I__2372\ : Sp12to4
    port map (
            O => \N__25579\,
            I => \N__25576\
        );

    \I__2371\ : Span12Mux_h
    port map (
            O => \N__25576\,
            I => \N__25573\
        );

    \I__2370\ : Span12Mux_v
    port map (
            O => \N__25573\,
            I => \N__25570\
        );

    \I__2369\ : Odrv12
    port map (
            O => \N__25570\,
            I => \PIN_7_c\
        );

    \I__2368\ : InMux
    port map (
            O => \N__25567\,
            I => \N__25558\
        );

    \I__2367\ : InMux
    port map (
            O => \N__25566\,
            I => \N__25558\
        );

    \I__2366\ : InMux
    port map (
            O => \N__25565\,
            I => \N__25558\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__25558\,
            I => \quadA_delayed\
        );

    \I__2364\ : InMux
    port map (
            O => \N__25555\,
            I => \N__25551\
        );

    \I__2363\ : InMux
    port map (
            O => \N__25554\,
            I => \N__25548\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__25551\,
            I => \quad_counter0.a_delay_counter_15\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__25548\,
            I => \quad_counter0.a_delay_counter_15\
        );

    \I__2360\ : InMux
    port map (
            O => \N__25543\,
            I => \N__25539\
        );

    \I__2359\ : InMux
    port map (
            O => \N__25542\,
            I => \N__25536\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__25539\,
            I => \quad_counter0.a_delay_counter_8\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__25536\,
            I => \quad_counter0.a_delay_counter_8\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__25531\,
            I => \N__25527\
        );

    \I__2355\ : InMux
    port map (
            O => \N__25530\,
            I => \N__25524\
        );

    \I__2354\ : InMux
    port map (
            O => \N__25527\,
            I => \N__25521\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__25524\,
            I => \quad_counter0.a_delay_counter_1\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__25521\,
            I => \quad_counter0.a_delay_counter_1\
        );

    \I__2351\ : InMux
    port map (
            O => \N__25516\,
            I => \N__25512\
        );

    \I__2350\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25509\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__25512\,
            I => \quad_counter0.a_delay_counter_6\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__25509\,
            I => \quad_counter0.a_delay_counter_6\
        );

    \I__2347\ : InMux
    port map (
            O => \N__25504\,
            I => \N__25500\
        );

    \I__2346\ : InMux
    port map (
            O => \N__25503\,
            I => \N__25497\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__25500\,
            I => \quad_counter0.a_delay_counter_9\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__25497\,
            I => \quad_counter0.a_delay_counter_9\
        );

    \I__2343\ : InMux
    port map (
            O => \N__25492\,
            I => \N__25488\
        );

    \I__2342\ : InMux
    port map (
            O => \N__25491\,
            I => \N__25485\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__25488\,
            I => \quad_counter0.a_delay_counter_7\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__25485\,
            I => \quad_counter0.a_delay_counter_7\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__25480\,
            I => \quad_counter0.n18_cascade_\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__25477\,
            I => \N__25474\
        );

    \I__2337\ : InMux
    port map (
            O => \N__25474\,
            I => \N__25469\
        );

    \I__2336\ : InMux
    port map (
            O => \N__25473\,
            I => \N__25466\
        );

    \I__2335\ : InMux
    port map (
            O => \N__25472\,
            I => \N__25463\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__25469\,
            I => a_delay_counter_0
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__25466\,
            I => a_delay_counter_0
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__25463\,
            I => a_delay_counter_0
        );

    \I__2331\ : CascadeMux
    port map (
            O => \N__25456\,
            I => \quad_counter0.n20_cascade_\
        );

    \I__2330\ : InMux
    port map (
            O => \N__25453\,
            I => \N__25449\
        );

    \I__2329\ : InMux
    port map (
            O => \N__25452\,
            I => \N__25446\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__25449\,
            I => \quad_counter0.a_delay_counter_2\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__25446\,
            I => \quad_counter0.a_delay_counter_2\
        );

    \I__2326\ : InMux
    port map (
            O => \N__25441\,
            I => \N__25435\
        );

    \I__2325\ : InMux
    port map (
            O => \N__25440\,
            I => \N__25435\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__25435\,
            I => n11349
        );

    \I__2323\ : InMux
    port map (
            O => \N__25432\,
            I => \N__25428\
        );

    \I__2322\ : InMux
    port map (
            O => \N__25431\,
            I => \N__25425\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__25428\,
            I => \quad_counter0.a_delay_counter_5\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__25425\,
            I => \quad_counter0.a_delay_counter_5\
        );

    \I__2319\ : InMux
    port map (
            O => \N__25420\,
            I => \N__25416\
        );

    \I__2318\ : InMux
    port map (
            O => \N__25419\,
            I => \N__25413\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__25416\,
            I => \quad_counter0.a_delay_counter_10\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__25413\,
            I => \quad_counter0.a_delay_counter_10\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__25408\,
            I => \N__25404\
        );

    \I__2314\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25401\
        );

    \I__2313\ : InMux
    port map (
            O => \N__25404\,
            I => \N__25398\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__25401\,
            I => \quad_counter0.a_delay_counter_12\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__25398\,
            I => \quad_counter0.a_delay_counter_12\
        );

    \I__2310\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25389\
        );

    \I__2309\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25386\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__25389\,
            I => \quad_counter0.a_delay_counter_3\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__25386\,
            I => \quad_counter0.a_delay_counter_3\
        );

    \I__2306\ : InMux
    port map (
            O => \N__25381\,
            I => \N__25378\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__25378\,
            I => \quad_counter0.n20954\
        );

    \I__2304\ : InMux
    port map (
            O => \N__25375\,
            I => \N__25371\
        );

    \I__2303\ : InMux
    port map (
            O => \N__25374\,
            I => \N__25368\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__25371\,
            I => \quad_counter0.a_delay_counter_4\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__25368\,
            I => \quad_counter0.a_delay_counter_4\
        );

    \I__2300\ : InMux
    port map (
            O => \N__25363\,
            I => \N__25359\
        );

    \I__2299\ : InMux
    port map (
            O => \N__25362\,
            I => \N__25356\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__25359\,
            I => \quad_counter0.a_delay_counter_11\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__25356\,
            I => \quad_counter0.a_delay_counter_11\
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__25351\,
            I => \N__25347\
        );

    \I__2295\ : InMux
    port map (
            O => \N__25350\,
            I => \N__25344\
        );

    \I__2294\ : InMux
    port map (
            O => \N__25347\,
            I => \N__25341\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__25344\,
            I => \quad_counter0.a_delay_counter_14\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__25341\,
            I => \quad_counter0.a_delay_counter_14\
        );

    \I__2291\ : InMux
    port map (
            O => \N__25336\,
            I => \N__25332\
        );

    \I__2290\ : InMux
    port map (
            O => \N__25335\,
            I => \N__25329\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__25332\,
            I => \quad_counter0.a_delay_counter_13\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__25329\,
            I => \quad_counter0.a_delay_counter_13\
        );

    \I__2287\ : InMux
    port map (
            O => \N__25324\,
            I => \N__25321\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__25321\,
            I => \quad_counter0.n19\
        );

    \I__2285\ : SRMux
    port map (
            O => \N__25318\,
            I => \N__25315\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__25315\,
            I => \N__25312\
        );

    \I__2283\ : Span4Mux_h
    port map (
            O => \N__25312\,
            I => \N__25309\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__25309\,
            I => \c0.n18649\
        );

    \I__2281\ : SRMux
    port map (
            O => \N__25306\,
            I => \N__25303\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__25303\,
            I => \c0.n18639\
        );

    \I__2279\ : SRMux
    port map (
            O => \N__25300\,
            I => \N__25297\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__25297\,
            I => \N__25294\
        );

    \I__2277\ : Span4Mux_v
    port map (
            O => \N__25294\,
            I => \N__25291\
        );

    \I__2276\ : Odrv4
    port map (
            O => \N__25291\,
            I => \c0.n18663\
        );

    \I__2275\ : SRMux
    port map (
            O => \N__25288\,
            I => \N__25285\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__25285\,
            I => \N__25281\
        );

    \I__2273\ : SRMux
    port map (
            O => \N__25284\,
            I => \N__25278\
        );

    \I__2272\ : Span4Mux_h
    port map (
            O => \N__25281\,
            I => \N__25272\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__25278\,
            I => \N__25272\
        );

    \I__2270\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25269\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__25272\,
            I => \a_delay_counter_15__N_2916\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__25269\,
            I => \a_delay_counter_15__N_2916\
        );

    \I__2267\ : InMux
    port map (
            O => \N__25264\,
            I => \N__25261\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__25261\,
            I => \quad_counter0.n13266\
        );

    \I__2265\ : InMux
    port map (
            O => \N__25258\,
            I => \N__25253\
        );

    \I__2264\ : InMux
    port map (
            O => \N__25257\,
            I => \N__25250\
        );

    \I__2263\ : InMux
    port map (
            O => \N__25256\,
            I => \N__25247\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__25253\,
            I => \quad_counter0.b_delay_counter_14\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__25250\,
            I => \quad_counter0.b_delay_counter_14\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__25247\,
            I => \quad_counter0.b_delay_counter_14\
        );

    \I__2259\ : InMux
    port map (
            O => \N__25240\,
            I => \N__25237\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__25237\,
            I => \quad_counter0.n13248\
        );

    \I__2257\ : InMux
    port map (
            O => \N__25234\,
            I => \N__25229\
        );

    \I__2256\ : InMux
    port map (
            O => \N__25233\,
            I => \N__25226\
        );

    \I__2255\ : InMux
    port map (
            O => \N__25232\,
            I => \N__25223\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__25229\,
            I => \N__25220\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__25226\,
            I => \quad_counter0.b_delay_counter_8\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__25223\,
            I => \quad_counter0.b_delay_counter_8\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__25220\,
            I => \quad_counter0.b_delay_counter_8\
        );

    \I__2250\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25210\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__25210\,
            I => \N__25207\
        );

    \I__2248\ : Odrv4
    port map (
            O => \N__25207\,
            I => \quad_counter0.n13203\
        );

    \I__2247\ : InMux
    port map (
            O => \N__25204\,
            I => \N__25199\
        );

    \I__2246\ : InMux
    port map (
            O => \N__25203\,
            I => \N__25196\
        );

    \I__2245\ : CascadeMux
    port map (
            O => \N__25202\,
            I => \N__25193\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__25199\,
            I => \N__25188\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__25196\,
            I => \N__25188\
        );

    \I__2242\ : InMux
    port map (
            O => \N__25193\,
            I => \N__25185\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__25188\,
            I => \quad_counter0.b_delay_counter_6\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__25185\,
            I => \quad_counter0.b_delay_counter_6\
        );

    \I__2239\ : InMux
    port map (
            O => \N__25180\,
            I => \N__25176\
        );

    \I__2238\ : InMux
    port map (
            O => \N__25179\,
            I => \N__25173\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__25176\,
            I => \N__25167\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__25173\,
            I => \N__25167\
        );

    \I__2235\ : InMux
    port map (
            O => \N__25172\,
            I => \N__25164\
        );

    \I__2234\ : Odrv4
    port map (
            O => \N__25167\,
            I => \quad_counter0.b_delay_counter_0\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__25164\,
            I => \quad_counter0.b_delay_counter_0\
        );

    \I__2232\ : InMux
    port map (
            O => \N__25159\,
            I => \N__25156\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__25156\,
            I => \quad_counter0.n13251\
        );

    \I__2230\ : InMux
    port map (
            O => \N__25153\,
            I => \N__25148\
        );

    \I__2229\ : InMux
    port map (
            O => \N__25152\,
            I => \N__25145\
        );

    \I__2228\ : InMux
    port map (
            O => \N__25151\,
            I => \N__25142\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__25148\,
            I => \quad_counter0.b_delay_counter_9\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__25145\,
            I => \quad_counter0.b_delay_counter_9\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__25142\,
            I => \quad_counter0.b_delay_counter_9\
        );

    \I__2224\ : InMux
    port map (
            O => \N__25135\,
            I => \N__25132\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__25132\,
            I => \N__25129\
        );

    \I__2222\ : Odrv4
    port map (
            O => \N__25129\,
            I => \quad_counter0.n13194\
        );

    \I__2221\ : InMux
    port map (
            O => \N__25126\,
            I => \N__25122\
        );

    \I__2220\ : InMux
    port map (
            O => \N__25125\,
            I => \N__25119\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__25122\,
            I => \N__25113\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__25119\,
            I => \N__25113\
        );

    \I__2217\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25110\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__25113\,
            I => \quad_counter0.b_delay_counter_3\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__25110\,
            I => \quad_counter0.b_delay_counter_3\
        );

    \I__2214\ : InMux
    port map (
            O => \N__25105\,
            I => \N__25102\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__25102\,
            I => \N__25099\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__25099\,
            I => \quad_counter0.n13200\
        );

    \I__2211\ : InMux
    port map (
            O => \N__25096\,
            I => \N__25092\
        );

    \I__2210\ : InMux
    port map (
            O => \N__25095\,
            I => \N__25089\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__25092\,
            I => \N__25083\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__25089\,
            I => \N__25083\
        );

    \I__2207\ : InMux
    port map (
            O => \N__25088\,
            I => \N__25080\
        );

    \I__2206\ : Odrv12
    port map (
            O => \N__25083\,
            I => \quad_counter0.b_delay_counter_5\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__25080\,
            I => \quad_counter0.b_delay_counter_5\
        );

    \I__2204\ : InMux
    port map (
            O => \N__25075\,
            I => \quad_counter0.n17216\
        );

    \I__2203\ : InMux
    port map (
            O => \N__25072\,
            I => \N__25068\
        );

    \I__2202\ : InMux
    port map (
            O => \N__25071\,
            I => \N__25065\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__25068\,
            I => \N__25059\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__25065\,
            I => \N__25059\
        );

    \I__2199\ : InMux
    port map (
            O => \N__25064\,
            I => \N__25056\
        );

    \I__2198\ : Span4Mux_v
    port map (
            O => \N__25059\,
            I => \N__25051\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__25056\,
            I => \N__25051\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__25051\,
            I => \quad_counter0.b_delay_counter_11\
        );

    \I__2195\ : InMux
    port map (
            O => \N__25048\,
            I => \N__25045\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__25045\,
            I => \N__25042\
        );

    \I__2193\ : Odrv12
    port map (
            O => \N__25042\,
            I => \quad_counter0.n13257\
        );

    \I__2192\ : InMux
    port map (
            O => \N__25039\,
            I => \quad_counter0.n17217\
        );

    \I__2191\ : InMux
    port map (
            O => \N__25036\,
            I => \quad_counter0.n17218\
        );

    \I__2190\ : InMux
    port map (
            O => \N__25033\,
            I => \N__25028\
        );

    \I__2189\ : InMux
    port map (
            O => \N__25032\,
            I => \N__25025\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__25031\,
            I => \N__25022\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__25028\,
            I => \N__25017\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__25025\,
            I => \N__25017\
        );

    \I__2185\ : InMux
    port map (
            O => \N__25022\,
            I => \N__25014\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__25017\,
            I => \quad_counter0.b_delay_counter_13\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__25014\,
            I => \quad_counter0.b_delay_counter_13\
        );

    \I__2182\ : InMux
    port map (
            O => \N__25009\,
            I => \N__25006\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__25006\,
            I => \N__25003\
        );

    \I__2180\ : Odrv4
    port map (
            O => \N__25003\,
            I => \quad_counter0.n13263\
        );

    \I__2179\ : InMux
    port map (
            O => \N__25000\,
            I => \quad_counter0.n17219\
        );

    \I__2178\ : InMux
    port map (
            O => \N__24997\,
            I => \quad_counter0.n17220\
        );

    \I__2177\ : InMux
    port map (
            O => \N__24994\,
            I => \quad_counter0.n17221\
        );

    \I__2176\ : InMux
    port map (
            O => \N__24991\,
            I => \N__24988\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__24988\,
            I => \quad_counter0.n13260\
        );

    \I__2174\ : InMux
    port map (
            O => \N__24985\,
            I => \N__24980\
        );

    \I__2173\ : InMux
    port map (
            O => \N__24984\,
            I => \N__24977\
        );

    \I__2172\ : InMux
    port map (
            O => \N__24983\,
            I => \N__24974\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__24980\,
            I => \quad_counter0.b_delay_counter_12\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__24977\,
            I => \quad_counter0.b_delay_counter_12\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__24974\,
            I => \quad_counter0.b_delay_counter_12\
        );

    \I__2168\ : InMux
    port map (
            O => \N__24967\,
            I => \N__24964\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__24964\,
            I => \N__24961\
        );

    \I__2166\ : Odrv4
    port map (
            O => \N__24961\,
            I => \quad_counter0.n13444\
        );

    \I__2165\ : InMux
    port map (
            O => \N__24958\,
            I => \N__24955\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__24955\,
            I => \quad_counter0.n13182\
        );

    \I__2163\ : InMux
    port map (
            O => \N__24952\,
            I => \quad_counter0.n17207\
        );

    \I__2162\ : InMux
    port map (
            O => \N__24949\,
            I => \quad_counter0.n17208\
        );

    \I__2161\ : InMux
    port map (
            O => \N__24946\,
            I => \quad_counter0.n17209\
        );

    \I__2160\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24939\
        );

    \I__2159\ : InMux
    port map (
            O => \N__24942\,
            I => \N__24936\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__24939\,
            I => \N__24933\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__24936\,
            I => \N__24929\
        );

    \I__2156\ : Span4Mux_v
    port map (
            O => \N__24933\,
            I => \N__24926\
        );

    \I__2155\ : InMux
    port map (
            O => \N__24932\,
            I => \N__24923\
        );

    \I__2154\ : Span4Mux_v
    port map (
            O => \N__24929\,
            I => \N__24916\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__24926\,
            I => \N__24916\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__24923\,
            I => \N__24916\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__24916\,
            I => \quad_counter0.b_delay_counter_4\
        );

    \I__2150\ : InMux
    port map (
            O => \N__24913\,
            I => \N__24910\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__24910\,
            I => \N__24907\
        );

    \I__2148\ : Span4Mux_h
    port map (
            O => \N__24907\,
            I => \N__24904\
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__24904\,
            I => \quad_counter0.n13197\
        );

    \I__2146\ : InMux
    port map (
            O => \N__24901\,
            I => \quad_counter0.n17210\
        );

    \I__2145\ : InMux
    port map (
            O => \N__24898\,
            I => \quad_counter0.n17211\
        );

    \I__2144\ : InMux
    port map (
            O => \N__24895\,
            I => \quad_counter0.n17212\
        );

    \I__2143\ : CascadeMux
    port map (
            O => \N__24892\,
            I => \N__24887\
        );

    \I__2142\ : InMux
    port map (
            O => \N__24891\,
            I => \N__24884\
        );

    \I__2141\ : InMux
    port map (
            O => \N__24890\,
            I => \N__24881\
        );

    \I__2140\ : InMux
    port map (
            O => \N__24887\,
            I => \N__24878\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__24884\,
            I => \quad_counter0.b_delay_counter_7\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__24881\,
            I => \quad_counter0.b_delay_counter_7\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__24878\,
            I => \quad_counter0.b_delay_counter_7\
        );

    \I__2136\ : InMux
    port map (
            O => \N__24871\,
            I => \N__24868\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__24868\,
            I => \quad_counter0.n13214\
        );

    \I__2134\ : InMux
    port map (
            O => \N__24865\,
            I => \quad_counter0.n17213\
        );

    \I__2133\ : InMux
    port map (
            O => \N__24862\,
            I => \bfn_9_15_0_\
        );

    \I__2132\ : InMux
    port map (
            O => \N__24859\,
            I => \quad_counter0.n17215\
        );

    \I__2131\ : InMux
    port map (
            O => \N__24856\,
            I => \N__24850\
        );

    \I__2130\ : InMux
    port map (
            O => \N__24855\,
            I => \N__24850\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__24850\,
            I => data_out_frame_5_1
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__24847\,
            I => \N__24844\
        );

    \I__2127\ : InMux
    port map (
            O => \N__24844\,
            I => \N__24838\
        );

    \I__2126\ : InMux
    port map (
            O => \N__24843\,
            I => \N__24838\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__24838\,
            I => data_out_frame_7_6
        );

    \I__2124\ : InMux
    port map (
            O => \N__24835\,
            I => \bfn_9_14_0_\
        );

    \I__2123\ : InMux
    port map (
            O => \N__24832\,
            I => \N__24827\
        );

    \I__2122\ : InMux
    port map (
            O => \N__24831\,
            I => \N__24824\
        );

    \I__2121\ : InMux
    port map (
            O => \N__24830\,
            I => \N__24821\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__24827\,
            I => \quad_counter0.b_delay_counter_1\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__24824\,
            I => \quad_counter0.b_delay_counter_1\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__24821\,
            I => \quad_counter0.b_delay_counter_1\
        );

    \I__2117\ : InMux
    port map (
            O => \N__24814\,
            I => \N__24808\
        );

    \I__2116\ : InMux
    port map (
            O => \N__24813\,
            I => \N__24808\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__24808\,
            I => data_out_frame_6_6
        );

    \I__2114\ : InMux
    port map (
            O => \N__24805\,
            I => \quad_counter0.n17236\
        );

    \I__2113\ : InMux
    port map (
            O => \N__24802\,
            I => \quad_counter0.n17227\
        );

    \I__2112\ : InMux
    port map (
            O => \N__24799\,
            I => \quad_counter0.n17228\
        );

    \I__2111\ : InMux
    port map (
            O => \N__24796\,
            I => \bfn_9_8_0_\
        );

    \I__2110\ : InMux
    port map (
            O => \N__24793\,
            I => \quad_counter0.n17230\
        );

    \I__2109\ : InMux
    port map (
            O => \N__24790\,
            I => \quad_counter0.n17231\
        );

    \I__2108\ : InMux
    port map (
            O => \N__24787\,
            I => \quad_counter0.n17232\
        );

    \I__2107\ : InMux
    port map (
            O => \N__24784\,
            I => \quad_counter0.n17233\
        );

    \I__2106\ : InMux
    port map (
            O => \N__24781\,
            I => \quad_counter0.n17234\
        );

    \I__2105\ : InMux
    port map (
            O => \N__24778\,
            I => \quad_counter0.n17235\
        );

    \I__2104\ : SRMux
    port map (
            O => \N__24775\,
            I => \N__24772\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__24772\,
            I => \c0.n18661\
        );

    \I__2102\ : InMux
    port map (
            O => \N__24769\,
            I => \N__24766\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__24766\,
            I => n39
        );

    \I__2100\ : InMux
    port map (
            O => \N__24763\,
            I => \bfn_9_7_0_\
        );

    \I__2099\ : InMux
    port map (
            O => \N__24760\,
            I => \quad_counter0.n17222\
        );

    \I__2098\ : InMux
    port map (
            O => \N__24757\,
            I => \quad_counter0.n17223\
        );

    \I__2097\ : InMux
    port map (
            O => \N__24754\,
            I => \quad_counter0.n17224\
        );

    \I__2096\ : InMux
    port map (
            O => \N__24751\,
            I => \quad_counter0.n17225\
        );

    \I__2095\ : InMux
    port map (
            O => \N__24748\,
            I => \quad_counter0.n17226\
        );

    \I__2094\ : IoInMux
    port map (
            O => \N__24745\,
            I => \N__24742\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__24742\,
            I => \N__24739\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__24739\,
            I => tx_enable
        );

    \I__2091\ : IoInMux
    port map (
            O => \N__24736\,
            I => \N__24733\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__24733\,
            I => \N__24729\
        );

    \I__2089\ : InMux
    port map (
            O => \N__24732\,
            I => \N__24726\
        );

    \I__2088\ : IoSpan4Mux
    port map (
            O => \N__24729\,
            I => \N__24723\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__24726\,
            I => \N__24720\
        );

    \I__2086\ : Span4Mux_s3_v
    port map (
            O => \N__24723\,
            I => \N__24717\
        );

    \I__2085\ : Span4Mux_h
    port map (
            O => \N__24720\,
            I => \N__24714\
        );

    \I__2084\ : Sp12to4
    port map (
            O => \N__24717\,
            I => \N__24711\
        );

    \I__2083\ : Span4Mux_v
    port map (
            O => \N__24714\,
            I => \N__24708\
        );

    \I__2082\ : Span12Mux_s11_v
    port map (
            O => \N__24711\,
            I => \N__24703\
        );

    \I__2081\ : Sp12to4
    port map (
            O => \N__24708\,
            I => \N__24703\
        );

    \I__2080\ : Span12Mux_v
    port map (
            O => \N__24703\,
            I => \N__24700\
        );

    \I__2079\ : Odrv12
    port map (
            O => \N__24700\,
            I => \LED_c\
        );

    \I__2078\ : SRMux
    port map (
            O => \N__24697\,
            I => \N__24694\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__24694\,
            I => \N__24691\
        );

    \I__2076\ : Span4Mux_h
    port map (
            O => \N__24691\,
            I => \N__24688\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__24688\,
            I => \c0.n18673\
        );

    \I__2074\ : IoInMux
    port map (
            O => \N__24685\,
            I => \N__24682\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__24682\,
            I => \N__24679\
        );

    \I__2072\ : IoSpan4Mux
    port map (
            O => \N__24679\,
            I => \N__24676\
        );

    \I__2071\ : IoSpan4Mux
    port map (
            O => \N__24676\,
            I => \N__24673\
        );

    \I__2070\ : IoSpan4Mux
    port map (
            O => \N__24673\,
            I => \N__24670\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__24670\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n17321\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n17329\,
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n17337\,
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n17345\,
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_10_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n17289\,
            carryinitout => \bfn_10_10_0_\
        );

    \IN_MUX_bfv_10_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n17297\,
            carryinitout => \bfn_10_11_0_\
        );

    \IN_MUX_bfv_10_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n17305\,
            carryinitout => \bfn_10_12_0_\
        );

    \IN_MUX_bfv_10_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n17313\,
            carryinitout => \bfn_10_13_0_\
        );

    \IN_MUX_bfv_12_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_5_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n17244\,
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_12_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_8_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n17259\,
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n17214\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n17229\,
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_18_0_\
        );

    \IN_MUX_bfv_10_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx.n17281\,
            carryinitout => \bfn_10_19_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_14_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_5_0_\
        );

    \IN_MUX_bfv_14_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17180_THRU_CRY_2_THRU_CO\,
            carryinitout => \bfn_14_6_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17181_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17182_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17183_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17184_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17185_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17186_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17187_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17188_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17189_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17190_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17191_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17192_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17193_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17194_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17195_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17196_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_14_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17197_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_23_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17198_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_24_0_\
        );

    \IN_MUX_bfv_14_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17199_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_25_0_\
        );

    \IN_MUX_bfv_14_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17200_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_26_0_\
        );

    \IN_MUX_bfv_14_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17201_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_27_0_\
        );

    \IN_MUX_bfv_14_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17202_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_28_0_\
        );

    \IN_MUX_bfv_14_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17203_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_29_0_\
        );

    \IN_MUX_bfv_14_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17204_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_30_0_\
        );

    \IN_MUX_bfv_14_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17205_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_31_0_\
        );

    \IN_MUX_bfv_14_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n17206_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_32_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__24685\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_I_0_1_lut_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34182\,
            lcout => tx_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_R_49_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24732\,
            lcout => \c0.rx.r_Rx_Data_R\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i0_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35721\,
            in1 => \N__31127\,
            in2 => \_gnd_net_\,
            in3 => \N__25720\,
            lcout => encoder0_position_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71023\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i4_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__26595\,
            in1 => \N__26478\,
            in2 => \_gnd_net_\,
            in3 => \N__24913\,
            lcout => \quad_counter0.b_delay_counter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71001\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.quadB_delayed_62_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26594\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \quadB_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70991\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i9_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29397\,
            in2 => \_gnd_net_\,
            in3 => \N__40555\,
            lcout => \c0.FRAME_MATCHER_state_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70993\,
            ce => 'H',
            sr => \N__24697\
        );

    \c0.i1_2_lut_adj_924_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29396\,
            in2 => \_gnd_net_\,
            in3 => \N__41472\,
            lcout => \c0.n18673\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_249_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27632\,
            in2 => \_gnd_net_\,
            in3 => \N__41449\,
            lcout => \c0.n18661\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i15_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27633\,
            in2 => \_gnd_net_\,
            in3 => \N__40554\,
            lcout => \c0.FRAME_MATCHER_state_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71007\,
            ce => 'H',
            sr => \N__24775\
        );

    \quad_counter0.a_delay_counter__i0_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__25277\,
            in1 => \N__24769\,
            in2 => \N__25477\,
            in3 => \N__25616\,
            lcout => a_delay_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71100\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_85_2_lut_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25473\,
            in2 => \_gnd_net_\,
            in3 => \N__24763\,
            lcout => n39,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \quad_counter0.n17222\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.a_delay_counter__i1_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25530\,
            in2 => \_gnd_net_\,
            in3 => \N__24760\,
            lcout => \quad_counter0.a_delay_counter_1\,
            ltout => OPEN,
            carryin => \quad_counter0.n17222\,
            carryout => \quad_counter0.n17223\,
            clk => \N__71086\,
            ce => \N__25617\,
            sr => \N__25284\
        );

    \quad_counter0.a_delay_counter__i2_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25453\,
            in2 => \_gnd_net_\,
            in3 => \N__24757\,
            lcout => \quad_counter0.a_delay_counter_2\,
            ltout => OPEN,
            carryin => \quad_counter0.n17223\,
            carryout => \quad_counter0.n17224\,
            clk => \N__71086\,
            ce => \N__25617\,
            sr => \N__25284\
        );

    \quad_counter0.a_delay_counter__i3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25393\,
            in2 => \_gnd_net_\,
            in3 => \N__24754\,
            lcout => \quad_counter0.a_delay_counter_3\,
            ltout => OPEN,
            carryin => \quad_counter0.n17224\,
            carryout => \quad_counter0.n17225\,
            clk => \N__71086\,
            ce => \N__25617\,
            sr => \N__25284\
        );

    \quad_counter0.a_delay_counter__i4_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25375\,
            in2 => \_gnd_net_\,
            in3 => \N__24751\,
            lcout => \quad_counter0.a_delay_counter_4\,
            ltout => OPEN,
            carryin => \quad_counter0.n17225\,
            carryout => \quad_counter0.n17226\,
            clk => \N__71086\,
            ce => \N__25617\,
            sr => \N__25284\
        );

    \quad_counter0.a_delay_counter__i5_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25432\,
            in2 => \_gnd_net_\,
            in3 => \N__24748\,
            lcout => \quad_counter0.a_delay_counter_5\,
            ltout => OPEN,
            carryin => \quad_counter0.n17226\,
            carryout => \quad_counter0.n17227\,
            clk => \N__71086\,
            ce => \N__25617\,
            sr => \N__25284\
        );

    \quad_counter0.a_delay_counter__i6_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25516\,
            in2 => \_gnd_net_\,
            in3 => \N__24802\,
            lcout => \quad_counter0.a_delay_counter_6\,
            ltout => OPEN,
            carryin => \quad_counter0.n17227\,
            carryout => \quad_counter0.n17228\,
            clk => \N__71086\,
            ce => \N__25617\,
            sr => \N__25284\
        );

    \quad_counter0.a_delay_counter__i7_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25492\,
            in2 => \_gnd_net_\,
            in3 => \N__24799\,
            lcout => \quad_counter0.a_delay_counter_7\,
            ltout => OPEN,
            carryin => \quad_counter0.n17228\,
            carryout => \quad_counter0.n17229\,
            clk => \N__71086\,
            ce => \N__25617\,
            sr => \N__25284\
        );

    \quad_counter0.a_delay_counter__i8_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25543\,
            in2 => \_gnd_net_\,
            in3 => \N__24796\,
            lcout => \quad_counter0.a_delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \quad_counter0.n17230\,
            clk => \N__71072\,
            ce => \N__25624\,
            sr => \N__25288\
        );

    \quad_counter0.a_delay_counter__i9_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25504\,
            in2 => \_gnd_net_\,
            in3 => \N__24793\,
            lcout => \quad_counter0.a_delay_counter_9\,
            ltout => OPEN,
            carryin => \quad_counter0.n17230\,
            carryout => \quad_counter0.n17231\,
            clk => \N__71072\,
            ce => \N__25624\,
            sr => \N__25288\
        );

    \quad_counter0.a_delay_counter__i10_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25420\,
            in2 => \_gnd_net_\,
            in3 => \N__24790\,
            lcout => \quad_counter0.a_delay_counter_10\,
            ltout => OPEN,
            carryin => \quad_counter0.n17231\,
            carryout => \quad_counter0.n17232\,
            clk => \N__71072\,
            ce => \N__25624\,
            sr => \N__25288\
        );

    \quad_counter0.a_delay_counter__i11_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25363\,
            in2 => \_gnd_net_\,
            in3 => \N__24787\,
            lcout => \quad_counter0.a_delay_counter_11\,
            ltout => OPEN,
            carryin => \quad_counter0.n17232\,
            carryout => \quad_counter0.n17233\,
            clk => \N__71072\,
            ce => \N__25624\,
            sr => \N__25288\
        );

    \quad_counter0.a_delay_counter__i12_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25407\,
            in2 => \_gnd_net_\,
            in3 => \N__24784\,
            lcout => \quad_counter0.a_delay_counter_12\,
            ltout => OPEN,
            carryin => \quad_counter0.n17233\,
            carryout => \quad_counter0.n17234\,
            clk => \N__71072\,
            ce => \N__25624\,
            sr => \N__25288\
        );

    \quad_counter0.a_delay_counter__i13_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25336\,
            in2 => \_gnd_net_\,
            in3 => \N__24781\,
            lcout => \quad_counter0.a_delay_counter_13\,
            ltout => OPEN,
            carryin => \quad_counter0.n17234\,
            carryout => \quad_counter0.n17235\,
            clk => \N__71072\,
            ce => \N__25624\,
            sr => \N__25288\
        );

    \quad_counter0.a_delay_counter__i14_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25350\,
            in2 => \_gnd_net_\,
            in3 => \N__24778\,
            lcout => \quad_counter0.a_delay_counter_14\,
            ltout => OPEN,
            carryin => \quad_counter0.n17235\,
            carryout => \quad_counter0.n17236\,
            clk => \N__71072\,
            ce => \N__25624\,
            sr => \N__25288\
        );

    \quad_counter0.a_delay_counter__i15_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25555\,
            in2 => \_gnd_net_\,
            in3 => \N__24805\,
            lcout => \quad_counter0.a_delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71072\,
            ce => \N__25624\,
            sr => \N__25288\
        );

    \quad_counter0.B_delayed_68_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26928\,
            lcout => \quad_counter0.B_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.B_65_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010101000"
        )
    port map (
            in0 => \N__26927\,
            in1 => \N__26257\,
            in2 => \N__26494\,
            in3 => \N__26614\,
            lcout => \B_filtered\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i1060_1_lut_2_lut_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__26881\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26903\,
            lcout => \quad_counter0.n2228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.A_filtered_I_0_2_lut_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__26882\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26904\,
            lcout => \quad_counter0.count_direction\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i2_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35720\,
            in1 => \N__25698\,
            in2 => \_gnd_net_\,
            in3 => \N__25681\,
            lcout => encoder0_position_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__2__5364_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25699\,
            in1 => \N__28473\,
            in2 => \_gnd_net_\,
            in3 => \N__46918\,
            lcout => data_out_frame_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i21_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35731\,
            in1 => \N__33458\,
            in2 => \_gnd_net_\,
            in3 => \N__25801\,
            lcout => encoder0_position_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i18_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35712\,
            in1 => \N__35756\,
            in2 => \_gnd_net_\,
            in3 => \N__25828\,
            lcout => encoder0_position_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i19_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__33002\,
            in1 => \N__35716\,
            in2 => \_gnd_net_\,
            in3 => \N__25819\,
            lcout => encoder0_position_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i20_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35713\,
            in1 => \N__27107\,
            in2 => \_gnd_net_\,
            in3 => \N__25810\,
            lcout => encoder0_position_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i11_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__26613\,
            in1 => \N__26493\,
            in2 => \_gnd_net_\,
            in3 => \N__25048\,
            lcout => \quad_counter0.b_delay_counter_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i22_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35714\,
            in1 => \N__25790\,
            in2 => \_gnd_net_\,
            in3 => \N__25771\,
            lcout => encoder0_position_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i23_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25762\,
            in1 => \N__33965\,
            in2 => \_gnd_net_\,
            in3 => \N__35717\,
            lcout => encoder0_position_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i24_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35715\,
            in1 => \N__32885\,
            in2 => \_gnd_net_\,
            in3 => \N__26011\,
            lcout => encoder0_position_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i25_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26002\,
            in1 => \N__27149\,
            in2 => \_gnd_net_\,
            in3 => \N__35718\,
            lcout => encoder0_position_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__6__5384_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46824\,
            in2 => \N__27055\,
            in3 => \N__24814\,
            lcout => data_out_frame_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71024\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__1__5397_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__41059\,
            in1 => \N__24856\,
            in2 => \N__46904\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71024\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24843\,
            in1 => \N__24813\,
            in2 => \_gnd_net_\,
            in3 => \N__40915\,
            lcout => \c0.n5_adj_3471\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__3__5363_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33204\,
            in1 => \N__25672\,
            in2 => \_gnd_net_\,
            in3 => \N__46826\,
            lcout => data_out_frame_9_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71024\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17971_3_lut_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__40914\,
            in1 => \N__24855\,
            in2 => \_gnd_net_\,
            in3 => \N__36965\,
            lcout => \c0.n21559\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__6__5376_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46825\,
            in2 => \N__24847\,
            in3 => \N__25791\,
            lcout => data_out_frame_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71024\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27085\,
            in1 => \N__26962\,
            in2 => \_gnd_net_\,
            in3 => \N__40935\,
            lcout => \c0.n5_adj_3033\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i13_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100001000100"
        )
    port map (
            in0 => \N__26615\,
            in1 => \N__25009\,
            in2 => \_gnd_net_\,
            in3 => \N__26483\,
            lcout => \quad_counter0.b_delay_counter_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71014\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i1_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100001000100"
        )
    port map (
            in0 => \N__26482\,
            in1 => \N__24958\,
            in2 => \_gnd_net_\,
            in3 => \N__26616\,
            lcout => \quad_counter0.b_delay_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71014\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i11_4_lut_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26032\,
            in1 => \N__25064\,
            in2 => \N__24892\,
            in3 => \N__24932\,
            lcout => \quad_counter0.n27_adj_2992\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i10_4_lut_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24830\,
            in1 => \N__26312\,
            in2 => \N__25031\,
            in3 => \N__25234\,
            lcout => \quad_counter0.n26_adj_2991\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i7_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000001010"
        )
    port map (
            in0 => \N__24871\,
            in1 => \_gnd_net_\,
            in2 => \N__26620\,
            in3 => \N__26484\,
            lcout => \quad_counter0.b_delay_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71014\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_2_lut_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25180\,
            in1 => \N__25179\,
            in2 => \N__26227\,
            in3 => \N__24835\,
            lcout => \quad_counter0.n13444\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \quad_counter0.n17207\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_3_lut_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__24832\,
            in1 => \N__24831\,
            in2 => \N__26231\,
            in3 => \N__24952\,
            lcout => \quad_counter0.n13182\,
            ltout => OPEN,
            carryin => \quad_counter0.n17207\,
            carryout => \quad_counter0.n17208\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_4_lut_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__26374\,
            in1 => \N__26373\,
            in2 => \N__26228\,
            in3 => \N__24949\,
            lcout => \quad_counter0.n13187\,
            ltout => OPEN,
            carryin => \quad_counter0.n17208\,
            carryout => \quad_counter0.n17209\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_5_lut_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25126\,
            in1 => \N__25125\,
            in2 => \N__26232\,
            in3 => \N__24946\,
            lcout => \quad_counter0.n13194\,
            ltout => OPEN,
            carryin => \quad_counter0.n17209\,
            carryout => \quad_counter0.n17210\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_6_lut_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__24942\,
            in1 => \N__24943\,
            in2 => \N__26229\,
            in3 => \N__24901\,
            lcout => \quad_counter0.n13197\,
            ltout => OPEN,
            carryin => \quad_counter0.n17210\,
            carryout => \quad_counter0.n17211\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_7_lut_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25096\,
            in1 => \N__25095\,
            in2 => \N__26233\,
            in3 => \N__24898\,
            lcout => \quad_counter0.n13200\,
            ltout => OPEN,
            carryin => \quad_counter0.n17211\,
            carryout => \quad_counter0.n17212\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_8_lut_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25204\,
            in1 => \N__25203\,
            in2 => \N__26230\,
            in3 => \N__24895\,
            lcout => \quad_counter0.n13203\,
            ltout => OPEN,
            carryin => \quad_counter0.n17212\,
            carryout => \quad_counter0.n17213\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_9_lut_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__24891\,
            in1 => \N__24890\,
            in2 => \N__26234\,
            in3 => \N__24865\,
            lcout => \quad_counter0.n13214\,
            ltout => OPEN,
            carryin => \quad_counter0.n17213\,
            carryout => \quad_counter0.n17214\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_10_lut_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25233\,
            in1 => \N__25232\,
            in2 => \N__26235\,
            in3 => \N__24862\,
            lcout => \quad_counter0.n13248\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \quad_counter0.n17215\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_11_lut_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25153\,
            in1 => \N__25152\,
            in2 => \N__26239\,
            in3 => \N__24859\,
            lcout => \quad_counter0.n13251\,
            ltout => OPEN,
            carryin => \quad_counter0.n17215\,
            carryout => \quad_counter0.n17216\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_12_lut_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__26031\,
            in1 => \N__26030\,
            in2 => \N__26236\,
            in3 => \N__25075\,
            lcout => \quad_counter0.n13254\,
            ltout => OPEN,
            carryin => \quad_counter0.n17216\,
            carryout => \quad_counter0.n17217\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_13_lut_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25072\,
            in1 => \N__25071\,
            in2 => \N__26240\,
            in3 => \N__25039\,
            lcout => \quad_counter0.n13257\,
            ltout => OPEN,
            carryin => \quad_counter0.n17217\,
            carryout => \quad_counter0.n17218\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_14_lut_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__24985\,
            in1 => \N__24984\,
            in2 => \N__26237\,
            in3 => \N__25036\,
            lcout => \quad_counter0.n13260\,
            ltout => OPEN,
            carryin => \quad_counter0.n17218\,
            carryout => \quad_counter0.n17219\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_15_lut_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25033\,
            in1 => \N__25032\,
            in2 => \N__26241\,
            in3 => \N__25000\,
            lcout => \quad_counter0.n13263\,
            ltout => OPEN,
            carryin => \quad_counter0.n17219\,
            carryout => \quad_counter0.n17220\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_16_lut_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25258\,
            in1 => \N__25257\,
            in2 => \N__26238\,
            in3 => \N__24997\,
            lcout => \quad_counter0.n13266\,
            ltout => OPEN,
            carryin => \quad_counter0.n17220\,
            carryout => \quad_counter0.n17221\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_17_lut_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__26313\,
            in1 => \N__26314\,
            in2 => \N__26242\,
            in3 => \N__24994\,
            lcout => \quad_counter0.n13269\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i12_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__26604\,
            in1 => \N__26486\,
            in2 => \_gnd_net_\,
            in3 => \N__24991\,
            lcout => \quad_counter0.b_delay_counter_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70995\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i12_4_lut_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__25256\,
            in1 => \N__24983\,
            in2 => \N__26366\,
            in3 => \N__25088\,
            lcout => \quad_counter0.n28_adj_2990\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i0_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__26603\,
            in1 => \N__26485\,
            in2 => \_gnd_net_\,
            in3 => \N__24967\,
            lcout => \quad_counter0.b_delay_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70995\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i14_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__26488\,
            in1 => \N__26605\,
            in2 => \_gnd_net_\,
            in3 => \N__25264\,
            lcout => \quad_counter0.b_delay_counter_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70995\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i8_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__26607\,
            in1 => \N__26487\,
            in2 => \_gnd_net_\,
            in3 => \N__25240\,
            lcout => \quad_counter0.b_delay_counter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70995\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i6_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__26489\,
            in1 => \N__26606\,
            in2 => \_gnd_net_\,
            in3 => \N__25213\,
            lcout => \quad_counter0.b_delay_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70995\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i9_4_lut_adj_206_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__25151\,
            in1 => \N__25118\,
            in2 => \N__25202\,
            in3 => \N__25172\,
            lcout => \quad_counter0.n25_adj_2993\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i9_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__26490\,
            in1 => \N__26608\,
            in2 => \_gnd_net_\,
            in3 => \N__25159\,
            lcout => \quad_counter0.b_delay_counter_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70995\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i3_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__26541\,
            in1 => \N__26491\,
            in2 => \_gnd_net_\,
            in3 => \N__25135\,
            lcout => \quad_counter0.b_delay_counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70992\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i5_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__26542\,
            in1 => \N__26492\,
            in2 => \_gnd_net_\,
            in3 => \N__25105\,
            lcout => \quad_counter0.b_delay_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70992\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i25_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29624\,
            in2 => \_gnd_net_\,
            in3 => \N__40542\,
            lcout => \c0.FRAME_MATCHER_state_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70996\,
            ce => 'H',
            sr => \N__25318\
        );

    \c0.i1_2_lut_adj_435_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29816\,
            in2 => \_gnd_net_\,
            in3 => \N__41471\,
            lcout => \c0.n18639\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_368_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29618\,
            in2 => \_gnd_net_\,
            in3 => \N__41470\,
            lcout => \c0.n18649\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i27_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40544\,
            in2 => \_gnd_net_\,
            in3 => \N__29817\,
            lcout => \c0.FRAME_MATCHER_state_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71008\,
            ce => 'H',
            sr => \N__25306\
        );

    \c0.i1_2_lut_adj_247_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29423\,
            in2 => \_gnd_net_\,
            in3 => \N__41393\,
            lcout => \c0.n18663\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i14_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29424\,
            in2 => \_gnd_net_\,
            in3 => \N__40540\,
            lcout => \c0.FRAME_MATCHER_state_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71025\,
            ce => 'H',
            sr => \N__25300\
        );

    \c0.i1_2_lut_adj_258_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27611\,
            in2 => \_gnd_net_\,
            in3 => \N__41469\,
            lcout => \c0.n18671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i24_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40541\,
            in2 => \_gnd_net_\,
            in3 => \N__29771\,
            lcout => \c0.FRAME_MATCHER_state_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71046\,
            ce => 'H',
            sr => \N__27952\
        );

    \quad_counter1.quadA_delayed_61_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28206\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \quadA_delayed_adj_3584\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71131\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.quadA_I_0_73_2_lut_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__25598\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25565\,
            lcout => \a_delay_counter_15__N_2916\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.A_63_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111001000000"
        )
    port map (
            in0 => \N__25441\,
            in1 => \N__25567\,
            in2 => \N__25600\,
            in3 => \N__26880\,
            lcout => \A_filtered\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71101\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101100110"
        )
    port map (
            in0 => \N__25566\,
            in1 => \N__25594\,
            in2 => \_gnd_net_\,
            in3 => \N__25440\,
            lcout => n12447,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.quadA_delayed_61_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25599\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \quadA_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71101\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i7_4_lut_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25554\,
            in1 => \N__25542\,
            in2 => \N__25531\,
            in3 => \N__25515\,
            lcout => OPEN,
            ltout => \quad_counter0.n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i9_4_lut_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25503\,
            in1 => \N__25491\,
            in2 => \N__25480\,
            in3 => \N__25381\,
            lcout => OPEN,
            ltout => \quad_counter0.n20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i2_4_lut_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__25324\,
            in1 => \N__25472\,
            in2 => \N__25456\,
            in3 => \N__25452\,
            lcout => n11349,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i3_4_lut_adj_205_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25431\,
            in1 => \N__25419\,
            in2 => \N__25408\,
            in3 => \N__25392\,
            lcout => \quad_counter0.n20954\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i1_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35640\,
            in1 => \N__27326\,
            in2 => \_gnd_net_\,
            in3 => \N__25708\,
            lcout => encoder0_position_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71073\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i8_4_lut_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25374\,
            in1 => \N__25362\,
            in2 => \N__25351\,
            in3 => \N__25335\,
            lcout => \quad_counter0.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i3_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35641\,
            in1 => \N__25661\,
            in2 => \_gnd_net_\,
            in3 => \N__25642\,
            lcout => encoder0_position_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71073\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_1_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25895\,
            in2 => \N__25955\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \quad_counter0.n17282\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_2_lut_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25726\,
            in2 => \N__31140\,
            in3 => \N__25711\,
            lcout => n2279,
            ltout => OPEN,
            carryin => \quad_counter0.n17282\,
            carryout => \quad_counter0.n17283\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_3_lut_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25896\,
            in2 => \N__27327\,
            in3 => \N__25702\,
            lcout => n2278,
            ltout => OPEN,
            carryin => \quad_counter0.n17283\,
            carryout => \quad_counter0.n17284\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_4_lut_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25697\,
            in2 => \N__25954\,
            in3 => \N__25675\,
            lcout => n2277,
            ltout => OPEN,
            carryin => \quad_counter0.n17284\,
            carryout => \quad_counter0.n17285\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_5_lut_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25900\,
            in2 => \N__25671\,
            in3 => \N__25636\,
            lcout => n2276,
            ltout => OPEN,
            carryin => \quad_counter0.n17285\,
            carryout => \quad_counter0.n17286\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_6_lut_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25905\,
            in2 => \N__27211\,
            in3 => \N__25633\,
            lcout => n2275,
            ltout => OPEN,
            carryin => \quad_counter0.n17286\,
            carryout => \quad_counter0.n17287\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_7_lut_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25901\,
            in2 => \N__26074\,
            in3 => \N__25630\,
            lcout => n2274,
            ltout => OPEN,
            carryin => \quad_counter0.n17287\,
            carryout => \quad_counter0.n17288\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_8_lut_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25906\,
            in2 => \N__27442\,
            in3 => \N__25627\,
            lcout => n2273,
            ltout => OPEN,
            carryin => \quad_counter0.n17288\,
            carryout => \quad_counter0.n17289\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_9_lut_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25907\,
            in2 => \N__27403\,
            in3 => \N__25753\,
            lcout => n2272,
            ltout => OPEN,
            carryin => \bfn_10_10_0_\,
            carryout => \quad_counter0.n17290\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_10_lut_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25911\,
            in2 => \N__30721\,
            in3 => \N__25750\,
            lcout => n2271,
            ltout => OPEN,
            carryin => \quad_counter0.n17290\,
            carryout => \quad_counter0.n17291\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_11_lut_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25908\,
            in2 => \N__30790\,
            in3 => \N__25747\,
            lcout => n2270,
            ltout => OPEN,
            carryin => \quad_counter0.n17291\,
            carryout => \quad_counter0.n17292\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_12_lut_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25912\,
            in2 => \N__27130\,
            in3 => \N__25744\,
            lcout => n2269,
            ltout => OPEN,
            carryin => \quad_counter0.n17292\,
            carryout => \quad_counter0.n17293\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_13_lut_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25909\,
            in2 => \N__33258\,
            in3 => \N__25741\,
            lcout => n2268,
            ltout => OPEN,
            carryin => \quad_counter0.n17293\,
            carryout => \quad_counter0.n17294\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_14_lut_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25913\,
            in2 => \N__28842\,
            in3 => \N__25738\,
            lcout => n2267,
            ltout => OPEN,
            carryin => \quad_counter0.n17294\,
            carryout => \quad_counter0.n17295\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_15_lut_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25910\,
            in2 => \N__28674\,
            in3 => \N__25735\,
            lcout => n2266,
            ltout => OPEN,
            carryin => \quad_counter0.n17295\,
            carryout => \quad_counter0.n17296\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_16_lut_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25914\,
            in2 => \N__27249\,
            in3 => \N__25732\,
            lcout => n2265,
            ltout => OPEN,
            carryin => \quad_counter0.n17296\,
            carryout => \quad_counter0.n17297\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_17_lut_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25956\,
            in2 => \N__27003\,
            in3 => \N__25729\,
            lcout => n2264,
            ltout => OPEN,
            carryin => \bfn_10_11_0_\,
            carryout => \quad_counter0.n17298\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_18_lut_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25959\,
            in2 => \N__27273\,
            in3 => \N__25834\,
            lcout => n2263,
            ltout => OPEN,
            carryin => \quad_counter0.n17298\,
            carryout => \quad_counter0.n17299\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_19_lut_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28721\,
            in2 => \N__25977\,
            in3 => \N__25831\,
            lcout => n2262,
            ltout => OPEN,
            carryin => \quad_counter0.n17299\,
            carryout => \quad_counter0.n17300\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_20_lut_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25963\,
            in2 => \N__35760\,
            in3 => \N__25822\,
            lcout => n2261,
            ltout => OPEN,
            carryin => \quad_counter0.n17300\,
            carryout => \quad_counter0.n17301\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_21_lut_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25957\,
            in2 => \N__33003\,
            in3 => \N__25813\,
            lcout => n2260,
            ltout => OPEN,
            carryin => \quad_counter0.n17301\,
            carryout => \quad_counter0.n17302\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_22_lut_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25964\,
            in2 => \N__27108\,
            in3 => \N__25804\,
            lcout => n2259,
            ltout => OPEN,
            carryin => \quad_counter0.n17302\,
            carryout => \quad_counter0.n17303\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_23_lut_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25958\,
            in2 => \N__33462\,
            in3 => \N__25795\,
            lcout => n2258,
            ltout => OPEN,
            carryin => \quad_counter0.n17303\,
            carryout => \quad_counter0.n17304\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_24_lut_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25965\,
            in2 => \N__25792\,
            in3 => \N__25765\,
            lcout => n2257,
            ltout => OPEN,
            carryin => \quad_counter0.n17304\,
            carryout => \quad_counter0.n17305\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_25_lut_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25966\,
            in2 => \N__33969\,
            in3 => \N__25756\,
            lcout => n2256,
            ltout => OPEN,
            carryin => \bfn_10_12_0_\,
            carryout => \quad_counter0.n17306\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_26_lut_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25970\,
            in2 => \N__32889\,
            in3 => \N__26005\,
            lcout => n2255,
            ltout => OPEN,
            carryin => \quad_counter0.n17306\,
            carryout => \quad_counter0.n17307\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_27_lut_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25967\,
            in2 => \N__27153\,
            in3 => \N__25996\,
            lcout => n2254,
            ltout => OPEN,
            carryin => \quad_counter0.n17307\,
            carryout => \quad_counter0.n17308\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_28_lut_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25971\,
            in2 => \N__35895\,
            in3 => \N__25993\,
            lcout => n2253,
            ltout => OPEN,
            carryin => \quad_counter0.n17308\,
            carryout => \quad_counter0.n17309\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_29_lut_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25968\,
            in2 => \N__35547\,
            in3 => \N__25990\,
            lcout => n2252,
            ltout => OPEN,
            carryin => \quad_counter0.n17309\,
            carryout => \quad_counter0.n17310\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_30_lut_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25972\,
            in2 => \N__27297\,
            in3 => \N__25987\,
            lcout => n2251,
            ltout => OPEN,
            carryin => \quad_counter0.n17310\,
            carryout => \quad_counter0.n17311\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_31_lut_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25969\,
            in2 => \N__33354\,
            in3 => \N__25984\,
            lcout => n2250,
            ltout => OPEN,
            carryin => \quad_counter0.n17311\,
            carryout => \quad_counter0.n17312\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_32_lut_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25973\,
            in2 => \N__27051\,
            in3 => \N__25981\,
            lcout => n2249,
            ltout => OPEN,
            carryin => \quad_counter0.n17312\,
            carryout => \quad_counter0.n17313\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_601_33_lut_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__43454\,
            in1 => \N__25978\,
            in2 => \_gnd_net_\,
            in3 => \N__25837\,
            lcout => n2248,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__0__5350_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30121\,
            in1 => \N__33606\,
            in2 => \_gnd_net_\,
            in3 => \N__46903\,
            lcout => data_out_frame_11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i4_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35709\,
            in1 => \N__27203\,
            in2 => \_gnd_net_\,
            in3 => \N__26119\,
            lcout => encoder0_position_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__3__5203_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__36033\,
            in1 => \N__46889\,
            in2 => \_gnd_net_\,
            in3 => \N__50362\,
            lcout => data_out_frame_29_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i7_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27398\,
            in1 => \N__35711\,
            in2 => \_gnd_net_\,
            in3 => \N__26107\,
            lcout => encoder0_position_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i5_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__35710\,
            in1 => \_gnd_net_\,
            in2 => \N__26073\,
            in3 => \N__26098\,
            lcout => encoder0_position_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i31_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35719\,
            in1 => \N__43455\,
            in2 => \_gnd_net_\,
            in3 => \N__26089\,
            lcout => encoder0_position_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17718_4_lut_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__26083\,
            in1 => \N__36953\,
            in2 => \N__33430\,
            in3 => \N__36700\,
            lcout => \c0.n21305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__5__5361_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26069\,
            in1 => \N__33102\,
            in2 => \_gnd_net_\,
            in3 => \N__46901\,
            lcout => data_out_frame_9_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71010\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n21629_bdd_4_lut_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__36699\,
            in1 => \N__26046\,
            in2 => \N__27226\,
            in3 => \N__26125\,
            lcout => \c0.n21632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__6__5360_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26047\,
            in1 => \N__27435\,
            in2 => \_gnd_net_\,
            in3 => \N__46902\,
            lcout => data_out_frame_9_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71010\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i10_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__26473\,
            in1 => \N__26610\,
            in2 => \_gnd_net_\,
            in3 => \N__26038\,
            lcout => \quad_counter0.b_delay_counter_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71003\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i15_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__26474\,
            in1 => \N__26611\,
            in2 => \_gnd_net_\,
            in3 => \N__26320\,
            lcout => \quad_counter0.b_delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71003\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__6__5352_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30646\,
            in1 => \N__26134\,
            in2 => \_gnd_net_\,
            in3 => \N__46723\,
            lcout => data_out_frame_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71003\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i15_4_lut_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26290\,
            in1 => \N__26281\,
            in2 => \N__26272\,
            in3 => \N__26263\,
            lcout => n11347,
            ltout => \n11347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i18016_4_lut_3_lut_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__26612\,
            in1 => \_gnd_net_\,
            in2 => \N__26245\,
            in3 => \N__26472\,
            lcout => \quad_counter0.n21603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_18044_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__26133\,
            in1 => \N__40857\,
            in2 => \N__28651\,
            in3 => \N__36701\,
            lcout => \c0.n21629\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i2_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__29282\,
            in1 => \N__29145\,
            in2 => \_gnd_net_\,
            in3 => \N__27556\,
            lcout => \c0.r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70998\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__4__5354_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36082\,
            in1 => \N__27472\,
            in2 => \_gnd_net_\,
            in3 => \N__46939\,
            lcout => data_out_frame_10_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70998\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__7__5367_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46938\,
            in1 => \N__27004\,
            in2 => \_gnd_net_\,
            in3 => \N__27168\,
            lcout => data_out_frame_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70998\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i0_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__29328\,
            in1 => \N__34065\,
            in2 => \N__29163\,
            in3 => \N__27523\,
            lcout => \c0.r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70998\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i2_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__26609\,
            in1 => \N__26471\,
            in2 => \_gnd_net_\,
            in3 => \N__26383\,
            lcout => \quad_counter0.b_delay_counter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70998\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i17744_3_lut_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28939\,
            in1 => \N__34161\,
            in2 => \_gnd_net_\,
            in3 => \N__34064\,
            lcout => OPEN,
            ltout => \c0.n21331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13772_4_lut_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__29280\,
            in1 => \N__27412\,
            in2 => \N__26347\,
            in3 => \N__29005\,
            lcout => OPEN,
            ltout => \c0.n17354_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_45_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__29032\,
            in1 => \N__26341\,
            in2 => \N__26344\,
            in3 => \N__29281\,
            lcout => tx_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70994\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17934_2_lut_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__29159\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27543\,
            lcout => \c0.n21521\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_4_lut_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__26712\,
            in1 => \N__26667\,
            in2 => \N__26731\,
            in3 => \N__26697\,
            lcout => OPEN,
            ltout => \c0.tx.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i12488_4_lut_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__26682\,
            in1 => \N__26652\,
            in2 => \N__26335\,
            in3 => \N__26637\,
            lcout => \c0.n15938\,
            ltout => \c0.n15938_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_4_lut_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34062\,
            in2 => \N__26332\,
            in3 => \N__29158\,
            lcout => \c0.tx.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i0_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26329\,
            in2 => \_gnd_net_\,
            in3 => \N__26323\,
            lcout => \c0.tx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_10_18_0_\,
            carryout => \c0.tx.n17274\,
            clk => \N__70999\,
            ce => \N__29199\,
            sr => \N__27651\
        );

    \c0.tx.r_Clock_Count__i1_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26730\,
            in2 => \_gnd_net_\,
            in3 => \N__26716\,
            lcout => \c0.tx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \c0.tx.n17274\,
            carryout => \c0.tx.n17275\,
            clk => \N__70999\,
            ce => \N__29199\,
            sr => \N__27651\
        );

    \c0.tx.r_Clock_Count__i2_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26713\,
            in2 => \_gnd_net_\,
            in3 => \N__26701\,
            lcout => \c0.tx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \c0.tx.n17275\,
            carryout => \c0.tx.n17276\,
            clk => \N__70999\,
            ce => \N__29199\,
            sr => \N__27651\
        );

    \c0.tx.r_Clock_Count__i3_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26698\,
            in2 => \_gnd_net_\,
            in3 => \N__26686\,
            lcout => \c0.tx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \c0.tx.n17276\,
            carryout => \c0.tx.n17277\,
            clk => \N__70999\,
            ce => \N__29199\,
            sr => \N__27651\
        );

    \c0.tx.r_Clock_Count__i4_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26683\,
            in2 => \_gnd_net_\,
            in3 => \N__26671\,
            lcout => \c0.tx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \c0.tx.n17277\,
            carryout => \c0.tx.n17278\,
            clk => \N__70999\,
            ce => \N__29199\,
            sr => \N__27651\
        );

    \c0.tx.r_Clock_Count__i5_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26668\,
            in2 => \_gnd_net_\,
            in3 => \N__26656\,
            lcout => \c0.tx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \c0.tx.n17278\,
            carryout => \c0.tx.n17279\,
            clk => \N__70999\,
            ce => \N__29199\,
            sr => \N__27651\
        );

    \c0.tx.r_Clock_Count__i6_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26653\,
            in2 => \_gnd_net_\,
            in3 => \N__26641\,
            lcout => \c0.tx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \c0.tx.n17279\,
            carryout => \c0.tx.n17280\,
            clk => \N__70999\,
            ce => \N__29199\,
            sr => \N__27651\
        );

    \c0.tx.r_Clock_Count__i7_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26638\,
            in2 => \_gnd_net_\,
            in3 => \N__26626\,
            lcout => \c0.tx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \c0.tx.n17280\,
            carryout => \c0.tx.n17281\,
            clk => \N__70999\,
            ce => \N__29199\,
            sr => \N__27651\
        );

    \c0.tx.r_Clock_Count__i8_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27681\,
            in2 => \_gnd_net_\,
            in3 => \N__26623\,
            lcout => \c0.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71004\,
            ce => \N__29203\,
            sr => \N__27655\
        );

    \c0.FRAME_MATCHER_state_i21_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31506\,
            in2 => \_gnd_net_\,
            in3 => \N__40480\,
            lcout => \c0.FRAME_MATCHER_state_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71017\,
            ce => 'H',
            sr => \N__31480\
        );

    \c0.FRAME_MATCHER_state_i6_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29548\,
            in2 => \_gnd_net_\,
            in3 => \N__40524\,
            lcout => \c0.FRAME_MATCHER_state_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71027\,
            ce => 'H',
            sr => \N__27568\
        );

    \c0.FRAME_MATCHER_state_i10_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27612\,
            in2 => \_gnd_net_\,
            in3 => \N__40525\,
            lcout => \c0.FRAME_MATCHER_state_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71036\,
            ce => 'H',
            sr => \N__26755\
        );

    \c0.FRAME_MATCHER_state_i13_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27770\,
            in2 => \_gnd_net_\,
            in3 => \N__40527\,
            lcout => \c0.FRAME_MATCHER_state_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71048\,
            ce => 'H',
            sr => \N__27751\
        );

    \c0.FRAME_MATCHER_state_i28_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29591\,
            in2 => \_gnd_net_\,
            in3 => \N__40529\,
            lcout => \c0.FRAME_MATCHER_state_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71060\,
            ce => 'H',
            sr => \N__26746\
        );

    \c0.i1_2_lut_adj_485_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29590\,
            in2 => \_gnd_net_\,
            in3 => \N__41476\,
            lcout => \c0.n18617\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.quadB_I_0_79_2_lut_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__26815\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26780\,
            lcout => \b_delay_counter_15__N_2933\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.quadB_delayed_62_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26816\,
            lcout => \quadB_delayed_adj_3585\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i9_4_lut_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__28026\,
            in1 => \N__27867\,
            in2 => \N__28075\,
            in3 => \N__27926\,
            lcout => OPEN,
            ltout => \quad_counter1.n25_adj_3577_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i15_4_lut_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26824\,
            in1 => \N__26767\,
            in2 => \N__26734\,
            in3 => \N__26761\,
            lcout => n11343,
            ltout => \n11343_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110010000"
        )
    port map (
            in0 => \N__26781\,
            in1 => \N__26817\,
            in2 => \N__26830\,
            in3 => \N__28231\,
            lcout => n12417,
            ltout => \n12417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.b_delay_counter__i0_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__27927\,
            in1 => \N__28245\,
            in2 => \N__26827\,
            in3 => \N__27913\,
            lcout => b_delay_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71132\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i12_4_lut_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__28089\,
            in1 => \N__28056\,
            in2 => \N__27886\,
            in3 => \N__28302\,
            lcout => \quad_counter1.n28_adj_3574\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.B_65_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011001000"
        )
    port map (
            in0 => \N__26818\,
            in1 => \N__29903\,
            in2 => \N__26791\,
            in3 => \N__26782\,
            lcout => \B_filtered_adj_3582\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71132\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i10_4_lut_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28284\,
            in1 => \N__28317\,
            in2 => \N__27904\,
            in3 => \N__28041\,
            lcout => \quad_counter1.n26_adj_3575\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i11_4_lut_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27996\,
            in1 => \N__28011\,
            in2 => \N__27982\,
            in3 => \N__27852\,
            lcout => \quad_counter1.n27_adj_3576\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.A_63_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111001000000"
        )
    port map (
            in0 => \N__26938\,
            in1 => \N__28213\,
            in2 => \N__28174\,
            in3 => \N__29857\,
            lcout => \A_filtered_adj_3581\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71102\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_951_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101100110"
        )
    port map (
            in0 => \N__28212\,
            in1 => \N__28170\,
            in2 => \_gnd_net_\,
            in3 => \N__26937\,
            lcout => n12477,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i3_4_lut_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28428\,
            in1 => \N__28530\,
            in2 => \N__28597\,
            in3 => \N__26890\,
            lcout => OPEN,
            ltout => \quad_counter1.n16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i11_4_lut_adj_946_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28443\,
            in1 => \N__28398\,
            in2 => \N__26944\,
            in3 => \N__26848\,
            lcout => OPEN,
            ltout => \quad_counter1.n24_adj_3578_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i12_4_lut_adj_947_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28116\,
            in1 => \N__28563\,
            in2 => \N__26941\,
            in3 => \N__28147\,
            lcout => n11351,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i30_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36247\,
            in1 => \N__30638\,
            in2 => \_gnd_net_\,
            in3 => \N__30616\,
            lcout => encoder1_position_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i3_4_lut_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26854\,
            in1 => \N__26883\,
            in2 => \N__26929\,
            in3 => \N__26908\,
            lcout => count_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i2_2_lut_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28548\,
            in2 => \_gnd_net_\,
            in3 => \N__28383\,
            lcout => \quad_counter1.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.A_delayed_67_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26884\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \quad_counter0.A_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i9_4_lut_adj_945_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28578\,
            in1 => \N__28413\,
            in2 => \N__28369\,
            in3 => \N__28332\,
            lcout => \quad_counter1.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i10_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35632\,
            in1 => \N__27128\,
            in2 => \_gnd_net_\,
            in3 => \N__26842\,
            lcout => encoder0_position_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71061\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i11_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__33257\,
            in1 => \N__35636\,
            in2 => \_gnd_net_\,
            in3 => \N__26836\,
            lcout => encoder0_position_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71061\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i12_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35633\,
            in1 => \N__28838\,
            in2 => \_gnd_net_\,
            in3 => \N__27028\,
            lcout => encoder0_position_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71061\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i13_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28673\,
            in1 => \N__35637\,
            in2 => \_gnd_net_\,
            in3 => \N__27022\,
            lcout => encoder0_position_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71061\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i14_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35634\,
            in1 => \N__27245\,
            in2 => \_gnd_net_\,
            in3 => \N__27016\,
            lcout => encoder0_position_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71061\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i15_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26996\,
            in1 => \N__35638\,
            in2 => \_gnd_net_\,
            in3 => \N__27010\,
            lcout => encoder0_position_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71061\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i16_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35635\,
            in1 => \N__27269\,
            in2 => \_gnd_net_\,
            in3 => \N__26974\,
            lcout => encoder0_position_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71061\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i17_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28725\,
            in1 => \N__35639\,
            in2 => \_gnd_net_\,
            in3 => \N__26968\,
            lcout => encoder0_position_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71061\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i18_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__33290\,
            in1 => \N__36248\,
            in2 => \_gnd_net_\,
            in3 => \N__30427\,
            lcout => encoder1_position_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__3__5387_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35548\,
            in1 => \N__35499\,
            in2 => \_gnd_net_\,
            in3 => \N__46934\,
            lcout => data_out_frame_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__4__5386_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46931\,
            in1 => \N__27298\,
            in2 => \_gnd_net_\,
            in3 => \N__26958\,
            lcout => data_out_frame_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__1__5389_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27345\,
            in1 => \N__27154\,
            in2 => \_gnd_net_\,
            in3 => \N__46933\,
            lcout => data_out_frame_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__2__5372_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46932\,
            in1 => \N__27129\,
            in2 => \_gnd_net_\,
            in3 => \N__28459\,
            lcout => data_out_frame_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__4__5378_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27109\,
            in1 => \N__27081\,
            in2 => \_gnd_net_\,
            in3 => \N__46935\,
            lcout => data_out_frame_7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i26_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35728\,
            in1 => \N__35891\,
            in2 => \_gnd_net_\,
            in3 => \N__27067\,
            lcout => encoder0_position_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i4_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30908\,
            in1 => \N__36258\,
            in2 => \_gnd_net_\,
            in3 => \N__30055\,
            lcout => encoder1_position_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i19_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36256\,
            in1 => \N__30407\,
            in2 => \_gnd_net_\,
            in3 => \N__30388\,
            lcout => encoder1_position_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i30_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35729\,
            in1 => \N__27047\,
            in2 => \_gnd_net_\,
            in3 => \N__27061\,
            lcout => encoder0_position_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17712_4_lut_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__33307\,
            in1 => \N__32749\,
            in2 => \N__36986\,
            in3 => \N__40919\,
            lcout => \c0.n21299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i7_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36257\,
            in1 => \N__29978\,
            in2 => \_gnd_net_\,
            in3 => \N__29959\,
            lcout => encoder1_position_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i8_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36356\,
            in1 => \N__36259\,
            in2 => \_gnd_net_\,
            in3 => \N__29944\,
            lcout => encoder1_position_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28704\,
            in1 => \N__27346\,
            in2 => \_gnd_net_\,
            in3 => \N__40905\,
            lcout => \c0.n5_adj_3102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__1__5365_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27331\,
            in1 => \N__31242\,
            in2 => \_gnd_net_\,
            in3 => \N__46736\,
            lcout => data_out_frame_9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71028\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i28_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27293\,
            in1 => \N__35688\,
            in2 => \_gnd_net_\,
            in3 => \N__27304\,
            lcout => encoder0_position_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71028\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__0__5382_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27274\,
            in1 => \N__33321\,
            in2 => \_gnd_net_\,
            in3 => \N__46735\,
            lcout => \c0.data_out_frame_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71028\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__6__5368_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46733\,
            in1 => \N__27250\,
            in2 => \_gnd_net_\,
            in3 => \N__27225\,
            lcout => data_out_frame_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71028\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__4__5362_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46734\,
            in1 => \N__27207\,
            in2 => \_gnd_net_\,
            in3 => \N__30828\,
            lcout => data_out_frame_9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71028\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17982_4_lut_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__36765\,
            in1 => \N__36952\,
            in2 => \N__27367\,
            in3 => \N__27184\,
            lcout => \c0.n21570\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17714_4_lut_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__29071\,
            in1 => \N__28693\,
            in2 => \N__37465\,
            in3 => \N__27178\,
            lcout => \c0.n21301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n21623_bdd_4_lut_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101111001000"
        )
    port map (
            in0 => \N__27375\,
            in1 => \N__33217\,
            in2 => \N__36766\,
            in3 => \N__27169\,
            lcout => OPEN,
            ltout => \c0.n21626_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17984_4_lut_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__36764\,
            in1 => \N__27358\,
            in2 => \N__27406\,
            in3 => \N__36951\,
            lcout => \c0.n21572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__7__5359_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27376\,
            in1 => \N__27402\,
            in2 => \_gnd_net_\,
            in3 => \N__46930\,
            lcout => data_out_frame_9_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__3__5347_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46929\,
            in1 => \N__30411\,
            in2 => \_gnd_net_\,
            in3 => \N__28869\,
            lcout => data_out_frame_11_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40855\,
            in1 => \N__28815\,
            in2 => \_gnd_net_\,
            in3 => \N__28741\,
            lcout => \c0.n11_adj_3472\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28960\,
            in1 => \N__28881\,
            in2 => \_gnd_net_\,
            in3 => \N__40853\,
            lcout => \c0.n11_adj_3479\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30889\,
            in1 => \N__37027\,
            in2 => \_gnd_net_\,
            in3 => \N__40854\,
            lcout => OPEN,
            ltout => \c0.n11_adj_3444_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17702_4_lut_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__36930\,
            in1 => \N__36702\,
            in2 => \N__27352\,
            in3 => \N__27460\,
            lcout => OPEN,
            ltout => \c0.n21289_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17989_4_lut_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__36703\,
            in1 => \N__30802\,
            in2 => \N__27349\,
            in3 => \N__36931\,
            lcout => \c0.n21577\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_adj_220_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29144\,
            in2 => \_gnd_net_\,
            in3 => \N__30955\,
            lcout => n6866,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_651_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__27687\,
            in1 => \N__34063\,
            in2 => \_gnd_net_\,
            in3 => \N__27514\,
            lcout => \c0.n55\,
            ltout => \c0.n55_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27490\,
            in3 => \N__29143\,
            lcout => OPEN,
            ltout => \c0.n14301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i1_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__29284\,
            in1 => \N__27484\,
            in2 => \N__27487\,
            in3 => \N__34085\,
            lcout => \r_SM_Main_1_adj_3592\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71005\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12492_2_lut_3_lut_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__27515\,
            in1 => \N__29142\,
            in2 => \_gnd_net_\,
            in3 => \N__27688\,
            lcout => \c0.n15942\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Active_47_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010011110000"
        )
    port map (
            in0 => \N__29283\,
            in1 => \N__27478\,
            in2 => \N__31295\,
            in3 => \N__29233\,
            lcout => tx_active,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71005\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17701_3_lut_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28768\,
            in1 => \N__27471\,
            in2 => \_gnd_net_\,
            in3 => \N__40856\,
            lcout => \c0.n21288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i6_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35687\,
            in1 => \N__27431\,
            in2 => \_gnd_net_\,
            in3 => \N__27454\,
            lcout => encoder0_position_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71005\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17930_3_lut_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__34060\,
            in1 => \N__29162\,
            in2 => \_gnd_net_\,
            in3 => \N__29056\,
            lcout => \c0.n21517\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_3_lut_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__29269\,
            in1 => \N__34059\,
            in2 => \_gnd_net_\,
            in3 => \N__27516\,
            lcout => \c0.tx.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17919_2_lut_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34226\,
            in2 => \_gnd_net_\,
            in3 => \N__29057\,
            lcout => OPEN,
            ltout => \c0.n21506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i2_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100011001100"
        )
    port map (
            in0 => \N__29272\,
            in1 => \N__27542\,
            in2 => \N__27559\,
            in3 => \N__28988\,
            lcout => \c0.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70997\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17898_4_lut_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__34228\,
            in1 => \N__27555\,
            in2 => \N__27544\,
            in3 => \N__29055\,
            lcout => OPEN,
            ltout => \c0.n21414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_4_lut_4_lut_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__29270\,
            in1 => \N__30943\,
            in2 => \N__27526\,
            in3 => \N__34061\,
            lcout => \c0.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i1_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110000001100"
        )
    port map (
            in0 => \N__34229\,
            in1 => \N__29058\,
            in2 => \N__28993\,
            in3 => \N__29271\,
            lcout => \c0.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__70997\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n21611_bdd_4_lut_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011000010"
        )
    port map (
            in0 => \N__31186\,
            in1 => \N__33991\,
            in2 => \N__34233\,
            in3 => \N__28945\,
            lcout => \c0.n21614\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_transmit_5164_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__39492\,
            in1 => \N__39071\,
            in2 => \N__38985\,
            in3 => \N__31519\,
            lcout => \c0.r_SM_Main_2_N_2547_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71006\,
            ce => 'H',
            sr => \N__31447\
        );

    \c0.i12472_2_lut_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__27517\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27678\,
            lcout => \c0.n15920\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_2_lut_4_lut_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__29161\,
            in1 => \N__34096\,
            in2 => \N__30952\,
            in3 => \N__29303\,
            lcout => n9377,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_3_lut_adj_219_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__27679\,
            in1 => \N__29160\,
            in2 => \_gnd_net_\,
            in3 => \N__27496\,
            lcout => OPEN,
            ltout => \c0.tx.n21179_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i18012_4_lut_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__27697\,
            in1 => \N__34097\,
            in2 => \N__27691\,
            in3 => \N__27680\,
            lcout => \c0.tx.n12759\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i26_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27798\,
            in2 => \_gnd_net_\,
            in3 => \N__40533\,
            lcout => \c0.FRAME_MATCHER_state_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71011\,
            ce => 'H',
            sr => \N__27784\
        );

    \c0.FRAME_MATCHER_state_i23_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40543\,
            in2 => \_gnd_net_\,
            in3 => \N__27737\,
            lcout => \c0.FRAME_MATCHER_state_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71019\,
            ce => 'H',
            sr => \N__27838\
        );

    \c0.FRAME_MATCHER_state_i31_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29356\,
            in2 => \_gnd_net_\,
            in3 => \N__40443\,
            lcout => \c0.FRAME_MATCHER_state_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71029\,
            ce => 'H',
            sr => \N__29083\
        );

    \c0.i4_4_lut_adj_688_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27771\,
            in1 => \N__27634\,
            in2 => \N__27613\,
            in3 => \N__27590\,
            lcout => \c0.n10_adj_3488\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i11_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27592\,
            in2 => \_gnd_net_\,
            in3 => \N__40522\,
            lcout => \c0.FRAME_MATCHER_state_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71038\,
            ce => 'H',
            sr => \N__27580\
        );

    \c0.i1_2_lut_adj_267_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27591\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41456\,
            lcout => \c0.n18669\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_268_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27718\,
            in2 => \_gnd_net_\,
            in3 => \N__41457\,
            lcout => \c0.n18651\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_269_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41458\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29553\,
            lcout => \c0.n18679\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_363_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27739\,
            in2 => \_gnd_net_\,
            in3 => \N__41459\,
            lcout => \c0.n18637\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_686_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27804\,
            in1 => \N__31502\,
            in2 => \N__29500\,
            in3 => \N__27824\,
            lcout => \c0.n10_adj_3438\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i22_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27826\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40523\,
            lcout => \c0.FRAME_MATCHER_state_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71050\,
            ce => 'H',
            sr => \N__27814\
        );

    \c0.i1_2_lut_adj_346_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27825\,
            in2 => \_gnd_net_\,
            in3 => \N__41462\,
            lcout => \c0.n18635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_370_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27805\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41463\,
            lcout => \c0.n18623\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_260_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27772\,
            in2 => \_gnd_net_\,
            in3 => \N__41460\,
            lcout => \c0.n18665\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_263_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41461\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29797\,
            lcout => \c0.n18641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_677_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34932\,
            in1 => \N__27738\,
            in2 => \N__31666\,
            in3 => \N__27710\,
            lcout => \c0.n16_adj_3484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i20_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__40526\,
            in1 => \_gnd_net_\,
            in2 => \N__27717\,
            in3 => \_gnd_net_\,
            lcout => \c0.FRAME_MATCHER_state_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71062\,
            ce => 'H',
            sr => \N__27964\
        );

    \c0.i1_2_lut_adj_366_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29775\,
            in2 => \_gnd_net_\,
            in3 => \N__41464\,
            lcout => \c0.n18625\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_851_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29735\,
            in2 => \_gnd_net_\,
            in3 => \N__41465\,
            lcout => \c0.n18677\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i19_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29796\,
            lcout => \c0.FRAME_MATCHER_state_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71074\,
            ce => 'H',
            sr => \N__27940\
        );

    \c0.FRAME_MATCHER_state_i3_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29452\,
            in2 => \_gnd_net_\,
            in3 => \N__40553\,
            lcout => \c0.FRAME_MATCHER_state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71087\,
            ce => 'H',
            sr => \N__29437\
        );

    \quad_counter1.add_86_2_lut_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27928\,
            in2 => \_gnd_net_\,
            in3 => \N__27907\,
            lcout => n187,
            ltout => OPEN,
            carryin => \bfn_12_5_0_\,
            carryout => \quad_counter1.n17237\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.b_delay_counter__i1_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27903\,
            in2 => \_gnd_net_\,
            in3 => \N__27889\,
            lcout => \quad_counter1.b_delay_counter_1\,
            ltout => OPEN,
            carryin => \quad_counter1.n17237\,
            carryout => \quad_counter1.n17238\,
            clk => \N__71149\,
            ce => \N__28273\,
            sr => \N__28244\
        );

    \quad_counter1.b_delay_counter__i2_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27885\,
            in2 => \_gnd_net_\,
            in3 => \N__27871\,
            lcout => \quad_counter1.b_delay_counter_2\,
            ltout => OPEN,
            carryin => \quad_counter1.n17238\,
            carryout => \quad_counter1.n17239\,
            clk => \N__71149\,
            ce => \N__28273\,
            sr => \N__28244\
        );

    \quad_counter1.b_delay_counter__i3_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27868\,
            in2 => \_gnd_net_\,
            in3 => \N__27856\,
            lcout => \quad_counter1.b_delay_counter_3\,
            ltout => OPEN,
            carryin => \quad_counter1.n17239\,
            carryout => \quad_counter1.n17240\,
            clk => \N__71149\,
            ce => \N__28273\,
            sr => \N__28244\
        );

    \quad_counter1.b_delay_counter__i4_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27853\,
            in2 => \_gnd_net_\,
            in3 => \N__27841\,
            lcout => \quad_counter1.b_delay_counter_4\,
            ltout => OPEN,
            carryin => \quad_counter1.n17240\,
            carryout => \quad_counter1.n17241\,
            clk => \N__71149\,
            ce => \N__28273\,
            sr => \N__28244\
        );

    \quad_counter1.b_delay_counter__i5_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28090\,
            in2 => \_gnd_net_\,
            in3 => \N__28078\,
            lcout => \quad_counter1.b_delay_counter_5\,
            ltout => OPEN,
            carryin => \quad_counter1.n17241\,
            carryout => \quad_counter1.n17242\,
            clk => \N__71149\,
            ce => \N__28273\,
            sr => \N__28244\
        );

    \quad_counter1.b_delay_counter__i6_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28074\,
            in2 => \_gnd_net_\,
            in3 => \N__28060\,
            lcout => \quad_counter1.b_delay_counter_6\,
            ltout => OPEN,
            carryin => \quad_counter1.n17242\,
            carryout => \quad_counter1.n17243\,
            clk => \N__71149\,
            ce => \N__28273\,
            sr => \N__28244\
        );

    \quad_counter1.b_delay_counter__i7_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28057\,
            in2 => \_gnd_net_\,
            in3 => \N__28045\,
            lcout => \quad_counter1.b_delay_counter_7\,
            ltout => OPEN,
            carryin => \quad_counter1.n17243\,
            carryout => \quad_counter1.n17244\,
            clk => \N__71149\,
            ce => \N__28273\,
            sr => \N__28244\
        );

    \quad_counter1.b_delay_counter__i8_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28042\,
            in2 => \_gnd_net_\,
            in3 => \N__28030\,
            lcout => \quad_counter1.b_delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \quad_counter1.n17245\,
            clk => \N__71134\,
            ce => \N__28266\,
            sr => \N__28246\
        );

    \quad_counter1.b_delay_counter__i9_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28027\,
            in2 => \_gnd_net_\,
            in3 => \N__28015\,
            lcout => \quad_counter1.b_delay_counter_9\,
            ltout => OPEN,
            carryin => \quad_counter1.n17245\,
            carryout => \quad_counter1.n17246\,
            clk => \N__71134\,
            ce => \N__28266\,
            sr => \N__28246\
        );

    \quad_counter1.b_delay_counter__i10_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28012\,
            in2 => \_gnd_net_\,
            in3 => \N__28000\,
            lcout => \quad_counter1.b_delay_counter_10\,
            ltout => OPEN,
            carryin => \quad_counter1.n17246\,
            carryout => \quad_counter1.n17247\,
            clk => \N__71134\,
            ce => \N__28266\,
            sr => \N__28246\
        );

    \quad_counter1.b_delay_counter__i11_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27997\,
            in2 => \_gnd_net_\,
            in3 => \N__27985\,
            lcout => \quad_counter1.b_delay_counter_11\,
            ltout => OPEN,
            carryin => \quad_counter1.n17247\,
            carryout => \quad_counter1.n17248\,
            clk => \N__71134\,
            ce => \N__28266\,
            sr => \N__28246\
        );

    \quad_counter1.b_delay_counter__i12_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27981\,
            in2 => \_gnd_net_\,
            in3 => \N__27967\,
            lcout => \quad_counter1.b_delay_counter_12\,
            ltout => OPEN,
            carryin => \quad_counter1.n17248\,
            carryout => \quad_counter1.n17249\,
            clk => \N__71134\,
            ce => \N__28266\,
            sr => \N__28246\
        );

    \quad_counter1.b_delay_counter__i13_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28318\,
            in2 => \_gnd_net_\,
            in3 => \N__28306\,
            lcout => \quad_counter1.b_delay_counter_13\,
            ltout => OPEN,
            carryin => \quad_counter1.n17249\,
            carryout => \quad_counter1.n17250\,
            clk => \N__71134\,
            ce => \N__28266\,
            sr => \N__28246\
        );

    \quad_counter1.b_delay_counter__i14_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28303\,
            in2 => \_gnd_net_\,
            in3 => \N__28291\,
            lcout => \quad_counter1.b_delay_counter_14\,
            ltout => OPEN,
            carryin => \quad_counter1.n17250\,
            carryout => \quad_counter1.n17251\,
            clk => \N__71134\,
            ce => \N__28266\,
            sr => \N__28246\
        );

    \quad_counter1.b_delay_counter__i15_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28285\,
            in2 => \_gnd_net_\,
            in3 => \N__28288\,
            lcout => \quad_counter1.b_delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71134\,
            ce => \N__28266\,
            sr => \N__28246\
        );

    \quad_counter1.quadA_I_0_73_2_lut_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28205\,
            in2 => \_gnd_net_\,
            in3 => \N__28169\,
            lcout => \a_delay_counter_15__N_2916_adj_3589\,
            ltout => \a_delay_counter_15__N_2916_adj_3589_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.a_delay_counter__i0_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__28126\,
            in1 => \N__28140\,
            in2 => \N__28150\,
            in3 => \N__28508\,
            lcout => a_delay_counter_0_adj_3583,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i7_3_lut_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__28351\,
            in1 => \N__28139\,
            in2 => \_gnd_net_\,
            in3 => \N__28101\,
            lcout => \quad_counter1.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_85_2_lut_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28141\,
            in2 => \_gnd_net_\,
            in3 => \N__28120\,
            lcout => n39_adj_3587,
            ltout => OPEN,
            carryin => \bfn_12_8_0_\,
            carryout => \quad_counter1.n17252\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.a_delay_counter__i1_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28117\,
            in2 => \_gnd_net_\,
            in3 => \N__28105\,
            lcout => \quad_counter1.a_delay_counter_1\,
            ltout => OPEN,
            carryin => \quad_counter1.n17252\,
            carryout => \quad_counter1.n17253\,
            clk => \N__71104\,
            ce => \N__28515\,
            sr => \N__28491\
        );

    \quad_counter1.a_delay_counter__i2_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28102\,
            in2 => \_gnd_net_\,
            in3 => \N__28447\,
            lcout => \quad_counter1.a_delay_counter_2\,
            ltout => OPEN,
            carryin => \quad_counter1.n17253\,
            carryout => \quad_counter1.n17254\,
            clk => \N__71104\,
            ce => \N__28515\,
            sr => \N__28491\
        );

    \quad_counter1.a_delay_counter__i3_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28444\,
            in2 => \_gnd_net_\,
            in3 => \N__28432\,
            lcout => \quad_counter1.a_delay_counter_3\,
            ltout => OPEN,
            carryin => \quad_counter1.n17254\,
            carryout => \quad_counter1.n17255\,
            clk => \N__71104\,
            ce => \N__28515\,
            sr => \N__28491\
        );

    \quad_counter1.a_delay_counter__i4_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28429\,
            in2 => \_gnd_net_\,
            in3 => \N__28417\,
            lcout => \quad_counter1.a_delay_counter_4\,
            ltout => OPEN,
            carryin => \quad_counter1.n17255\,
            carryout => \quad_counter1.n17256\,
            clk => \N__71104\,
            ce => \N__28515\,
            sr => \N__28491\
        );

    \quad_counter1.a_delay_counter__i5_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28414\,
            in2 => \_gnd_net_\,
            in3 => \N__28402\,
            lcout => \quad_counter1.a_delay_counter_5\,
            ltout => OPEN,
            carryin => \quad_counter1.n17256\,
            carryout => \quad_counter1.n17257\,
            clk => \N__71104\,
            ce => \N__28515\,
            sr => \N__28491\
        );

    \quad_counter1.a_delay_counter__i6_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28399\,
            in2 => \_gnd_net_\,
            in3 => \N__28387\,
            lcout => \quad_counter1.a_delay_counter_6\,
            ltout => OPEN,
            carryin => \quad_counter1.n17257\,
            carryout => \quad_counter1.n17258\,
            clk => \N__71104\,
            ce => \N__28515\,
            sr => \N__28491\
        );

    \quad_counter1.a_delay_counter__i7_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28384\,
            in2 => \_gnd_net_\,
            in3 => \N__28372\,
            lcout => \quad_counter1.a_delay_counter_7\,
            ltout => OPEN,
            carryin => \quad_counter1.n17258\,
            carryout => \quad_counter1.n17259\,
            clk => \N__71104\,
            ce => \N__28515\,
            sr => \N__28491\
        );

    \quad_counter1.a_delay_counter__i8_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28368\,
            in2 => \_gnd_net_\,
            in3 => \N__28354\,
            lcout => \quad_counter1.a_delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \quad_counter1.n17260\,
            clk => \N__71088\,
            ce => \N__28519\,
            sr => \N__28492\
        );

    \quad_counter1.a_delay_counter__i9_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28350\,
            in2 => \_gnd_net_\,
            in3 => \N__28336\,
            lcout => \quad_counter1.a_delay_counter_9\,
            ltout => OPEN,
            carryin => \quad_counter1.n17260\,
            carryout => \quad_counter1.n17261\,
            clk => \N__71088\,
            ce => \N__28519\,
            sr => \N__28492\
        );

    \quad_counter1.a_delay_counter__i10_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28333\,
            in2 => \_gnd_net_\,
            in3 => \N__28321\,
            lcout => \quad_counter1.a_delay_counter_10\,
            ltout => OPEN,
            carryin => \quad_counter1.n17261\,
            carryout => \quad_counter1.n17262\,
            clk => \N__71088\,
            ce => \N__28519\,
            sr => \N__28492\
        );

    \quad_counter1.a_delay_counter__i11_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28596\,
            in2 => \_gnd_net_\,
            in3 => \N__28582\,
            lcout => \quad_counter1.a_delay_counter_11\,
            ltout => OPEN,
            carryin => \quad_counter1.n17262\,
            carryout => \quad_counter1.n17263\,
            clk => \N__71088\,
            ce => \N__28519\,
            sr => \N__28492\
        );

    \quad_counter1.a_delay_counter__i12_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28579\,
            in2 => \_gnd_net_\,
            in3 => \N__28567\,
            lcout => \quad_counter1.a_delay_counter_12\,
            ltout => OPEN,
            carryin => \quad_counter1.n17263\,
            carryout => \quad_counter1.n17264\,
            clk => \N__71088\,
            ce => \N__28519\,
            sr => \N__28492\
        );

    \quad_counter1.a_delay_counter__i13_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28564\,
            in2 => \_gnd_net_\,
            in3 => \N__28552\,
            lcout => \quad_counter1.a_delay_counter_13\,
            ltout => OPEN,
            carryin => \quad_counter1.n17264\,
            carryout => \quad_counter1.n17265\,
            clk => \N__71088\,
            ce => \N__28519\,
            sr => \N__28492\
        );

    \quad_counter1.a_delay_counter__i14_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28549\,
            in2 => \_gnd_net_\,
            in3 => \N__28537\,
            lcout => \quad_counter1.a_delay_counter_14\,
            ltout => OPEN,
            carryin => \quad_counter1.n17265\,
            carryout => \quad_counter1.n17266\,
            clk => \N__71088\,
            ce => \N__28519\,
            sr => \N__28492\
        );

    \quad_counter1.a_delay_counter__i15_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28531\,
            in2 => \_gnd_net_\,
            in3 => \N__28534\,
            lcout => \quad_counter1.a_delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71088\,
            ce => \N__28519\,
            sr => \N__28492\
        );

    \quad_counter1.count_i0_i9_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36177\,
            in1 => \N__31163\,
            in2 => \_gnd_net_\,
            in3 => \N__29929\,
            lcout => encoder1_position_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i10_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30287\,
            in1 => \N__36178\,
            in2 => \_gnd_net_\,
            in3 => \N__30268\,
            lcout => encoder1_position_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i11_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36174\,
            in1 => \N__30251\,
            in2 => \_gnd_net_\,
            in3 => \N__30232\,
            lcout => encoder1_position_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n21647_bdd_4_lut_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__28474\,
            in1 => \N__36756\,
            in2 => \N__32824\,
            in3 => \N__28458\,
            lcout => \c0.n21650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i13_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36175\,
            in1 => \N__30218\,
            in2 => \_gnd_net_\,
            in3 => \N__30196\,
            lcout => encoder1_position_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i14_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30185\,
            in1 => \N__36179\,
            in2 => \_gnd_net_\,
            in3 => \N__30163\,
            lcout => encoder1_position_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i15_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36176\,
            in1 => \N__30149\,
            in2 => \_gnd_net_\,
            in3 => \N__30130\,
            lcout => encoder1_position_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i16_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30116\,
            in1 => \N__36180\,
            in2 => \_gnd_net_\,
            in3 => \N__30094\,
            lcout => encoder1_position_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17976_4_lut_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__36954\,
            in1 => \N__28618\,
            in2 => \N__36760\,
            in3 => \N__31006\,
            lcout => OPEN,
            ltout => \c0.n21564_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_3_lut_4_lut_adj_607_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__37336\,
            in1 => \N__37450\,
            in2 => \N__28612\,
            in3 => \N__35779\,
            lcout => n10_adj_3593,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i20_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30368\,
            in1 => \N__36246\,
            in2 => \_gnd_net_\,
            in3 => \N__30349\,
            lcout => encoder1_position_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71063\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i9_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30782\,
            in1 => \N__35730\,
            in2 => \_gnd_net_\,
            in3 => \N__28609\,
            lcout => encoder0_position_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71063\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i22_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36245\,
            in1 => \N__30335\,
            in2 => \_gnd_net_\,
            in3 => \N__30316\,
            lcout => encoder1_position_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71063\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i17_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31052\,
            in1 => \N__36224\,
            in2 => \_gnd_net_\,
            in3 => \N__30085\,
            lcout => encoder1_position_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i29_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__33350\,
            in1 => \N__35724\,
            in2 => \_gnd_net_\,
            in3 => \N__28687\,
            lcout => encoder0_position_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i24_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__36221\,
            in1 => \_gnd_net_\,
            in2 => \N__30762\,
            in3 => \N__30304\,
            lcout => encoder1_position_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__5__5337_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30220\,
            in1 => \N__30439\,
            in2 => \_gnd_net_\,
            in3 => \N__46732\,
            lcout => data_out_frame_12_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i26_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36222\,
            in1 => \N__32799\,
            in2 => \_gnd_net_\,
            in3 => \N__30694\,
            lcout => encoder1_position_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i27_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30661\,
            in1 => \N__36223\,
            in2 => \_gnd_net_\,
            in3 => \N__30680\,
            lcout => encoder1_position_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__5__5369_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46730\,
            in1 => \N__28678\,
            in2 => \_gnd_net_\,
            in3 => \N__33126\,
            lcout => data_out_frame_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__6__5344_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30336\,
            in1 => \N__28644\,
            in2 => \_gnd_net_\,
            in3 => \N__46731\,
            lcout => data_out_frame_11_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i8_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28630\,
            in1 => \N__35723\,
            in2 => \_gnd_net_\,
            in3 => \N__30714\,
            lcout => encoder0_position_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71039\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i2_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36260\,
            in1 => \N__31079\,
            in2 => \_gnd_net_\,
            in3 => \N__30073\,
            lcout => encoder1_position_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71039\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__4__5346_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30373\,
            in1 => \N__28767\,
            in2 => \_gnd_net_\,
            in3 => \N__46726\,
            lcout => data_out_frame_11_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71039\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__36475\,
            in1 => \N__36939\,
            in2 => \N__28753\,
            in3 => \N__36698\,
            lcout => \c0.n21653\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__6__5336_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30187\,
            in1 => \N__28740\,
            in2 => \_gnd_net_\,
            in3 => \N__46727\,
            lcout => data_out_frame_12_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71039\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i6_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36261\,
            in1 => \N__30029\,
            in2 => \_gnd_net_\,
            in3 => \N__30007\,
            lcout => encoder1_position_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71039\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__1__5381_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28726\,
            in1 => \N__28705\,
            in2 => \_gnd_net_\,
            in3 => \N__46728\,
            lcout => data_out_frame_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71039\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_475_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40975\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36940\,
            lcout => \c0.n6_adj_3324\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__2__5340_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30292\,
            in1 => \N__46923\,
            in2 => \_gnd_net_\,
            in3 => \N__31018\,
            lcout => data_out_frame_12_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__3__5331_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__46920\,
            in1 => \_gnd_net_\,
            in2 => \N__28894\,
            in3 => \N__33036\,
            lcout => data_out_frame_13_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__3__5355_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30685\,
            in1 => \N__46922\,
            in2 => \_gnd_net_\,
            in3 => \N__28855\,
            lcout => data_out_frame_10_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40881\,
            in1 => \N__28890\,
            in2 => \_gnd_net_\,
            in3 => \N__28909\,
            lcout => \c0.n11_adj_3404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__7__5335_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46919\,
            in1 => \N__30154\,
            in2 => \_gnd_net_\,
            in3 => \N__28882\,
            lcout => data_out_frame_12_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_18054_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__40880\,
            in1 => \N__36746\,
            in2 => \N__28870\,
            in3 => \N__28854\,
            lcout => \c0.n21641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__4__5370_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46921\,
            in1 => \N__28846\,
            in2 => \_gnd_net_\,
            in3 => \N__30814\,
            lcout => data_out_frame_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__6__5328_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30033\,
            in1 => \N__28816\,
            in2 => \_gnd_net_\,
            in3 => \N__46737\,
            lcout => data_out_frame_13_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71020\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_3_lut_4_lut_adj_609_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__28804\,
            in1 => \N__33556\,
            in2 => \N__37451\,
            in3 => \N__37341\,
            lcout => \c0.n7_adj_3333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n21653_bdd_4_lut_4_lut_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010011000"
        )
    port map (
            in0 => \N__40824\,
            in1 => \N__28798\,
            in2 => \N__30736\,
            in3 => \N__36908\,
            lcout => n21656,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17720_4_lut_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__37423\,
            in1 => \N__37523\,
            in2 => \N__35839\,
            in3 => \N__28789\,
            lcout => OPEN,
            ltout => \c0.n21307_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_3_lut_4_lut_adj_619_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__37342\,
            in1 => \N__28777\,
            in2 => \N__28771\,
            in3 => \N__37428\,
            lcout => n9_adj_3588,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17990_4_lut_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__37422\,
            in1 => \N__37522\,
            in2 => \N__33073\,
            in3 => \N__28975\,
            lcout => OPEN,
            ltout => \n21578_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i23_4_lut_adj_953_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__37340\,
            in1 => \N__37424\,
            in2 => \N__28969\,
            in3 => \N__28966\,
            lcout => n9_adj_3591,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__7__5327_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46622\,
            in1 => \N__29991\,
            in2 => \_gnd_net_\,
            in3 => \N__28959\,
            lcout => data_out_frame_13_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71012\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17927_2_lut_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31199\,
            in2 => \_gnd_net_\,
            in3 => \N__34084\,
            lcout => \c0.n21467\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i17743_3_lut_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34227\,
            in1 => \N__33931\,
            in2 => \_gnd_net_\,
            in3 => \N__28920\,
            lcout => \c0.tx.n21330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i6_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__33785\,
            in1 => \N__28921\,
            in2 => \N__33886\,
            in3 => \N__28927\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71012\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_643_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__36876\,
            in1 => \N__37316\,
            in2 => \_gnd_net_\,
            in3 => \N__36621\,
            lcout => \c0.n9753\,
            ltout => \c0.n9753_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_647_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28912\,
            in3 => \N__40823\,
            lcout => \c0.n9755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__3__5339_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30259\,
            in1 => \N__28908\,
            in2 => \_gnd_net_\,
            in3 => \N__46623\,
            lcout => data_out_frame_12_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71012\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17972_3_lut_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__37301\,
            in1 => \N__40739\,
            in2 => \_gnd_net_\,
            in3 => \N__36588\,
            lcout => \c0.n21456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_3_lut_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29059\,
            in1 => \N__29020\,
            in2 => \_gnd_net_\,
            in3 => \N__29038\,
            lcout => \c0.n32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i17742_3_lut_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34220\,
            in1 => \N__30853\,
            in2 => \_gnd_net_\,
            in3 => \N__29214\,
            lcout => \c0.n21329\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i0_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__29304\,
            in1 => \N__28992\,
            in2 => \_gnd_net_\,
            in3 => \N__34222\,
            lcout => \c0.r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_2__I_0_i2_3_lut_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34221\,
            in1 => \N__31362\,
            in2 => \_gnd_net_\,
            in3 => \N__31323\,
            lcout => OPEN,
            ltout => \c0.n2_adj_3556_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_3_lut_adj_904_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34098\,
            in2 => \N__29023\,
            in3 => \N__34160\,
            lcout => \c0.n7_adj_3557\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_935_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111100000"
        )
    port map (
            in0 => \N__34168\,
            in1 => \N__29186\,
            in2 => \N__29170\,
            in3 => \N__29014\,
            lcout => OPEN,
            ltout => \c0.n19001_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i31_3_lut_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29298\,
            in2 => \N__29008\,
            in3 => \N__29089\,
            lcout => \c0.n30_adj_3559\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_690_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39590\,
            in2 => \_gnd_net_\,
            in3 => \N__38968\,
            lcout => \c0.n6_adj_3338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_4_lut_4_lut_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__34095\,
            in1 => \N__29302\,
            in2 => \N__29329\,
            in3 => \N__29169\,
            lcout => \c0.n12498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_3_lut_4_lut_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001111"
        )
    port map (
            in0 => \N__29168\,
            in1 => \N__29324\,
            in2 => \N__29305\,
            in3 => \N__34094\,
            lcout => n4_adj_3580,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i4_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__33765\,
            in1 => \N__29215\,
            in2 => \N__33877\,
            in3 => \N__29224\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71013\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_1_lut_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34092\,
            lcout => \c0.n12512\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_3_lut_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34093\,
            in1 => \N__29164\,
            in2 => \_gnd_net_\,
            in3 => \N__34169\,
            lcout => \c0.n19023\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_691_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__37149\,
            in1 => \N__29527\,
            in2 => \_gnd_net_\,
            in3 => \N__37128\,
            lcout => \c0.n19052\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_2_lut_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56126\,
            in2 => \_gnd_net_\,
            in3 => \N__39232\,
            lcout => \c0.rx.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_390_Select_2_i2_4_lut_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__38972\,
            in1 => \N__42505\,
            in2 => \N__39076\,
            in3 => \N__35419\,
            lcout => n8112,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12190_4_lut_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001000"
        )
    port map (
            in0 => \N__29650\,
            in1 => \N__40284\,
            in2 => \N__38167\,
            in3 => \N__38194\,
            lcout => \c0.n4812\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_229_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29355\,
            in2 => \_gnd_net_\,
            in3 => \N__41404\,
            lcout => \c0.n18609\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17645_2_lut_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39486\,
            in2 => \_gnd_net_\,
            in3 => \N__29523\,
            lcout => \c0.n21231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_adj_915_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__31575\,
            in1 => \N__38245\,
            in2 => \N__31429\,
            in3 => \N__38325\,
            lcout => \c0.n21053\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_425_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38361\,
            in2 => \_gnd_net_\,
            in3 => \N__35208\,
            lcout => \c0.FRAME_MATCHER_state_31_N_1864_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_22_i6_2_lut_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60695\,
            in2 => \_gnd_net_\,
            in3 => \N__34390\,
            lcout => \c0.n6_adj_3178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_689_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__29425\,
            in1 => \N__29404\,
            in2 => \_gnd_net_\,
            in3 => \N__29377\,
            lcout => \c0.n15850\,
            ltout => \c0.n15850_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29469\,
            in1 => \N__29560\,
            in2 => \N__29371\,
            in3 => \N__29335\,
            lcout => \c0.n11427\,
            ltout => \c0.n11427_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_279_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29368\,
            in3 => \N__39568\,
            lcout => n11289,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_682_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40324\,
            in1 => \N__29365\,
            in2 => \N__29749\,
            in3 => \N__29354\,
            lcout => \c0.n19045\,
            ltout => \c0.n19045_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_586_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41505\,
            in1 => \N__29736\,
            in2 => \N__29338\,
            in3 => \N__29549\,
            lcout => \c0.n4_adj_3046\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_577_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29569\,
            in1 => \N__29626\,
            in2 => \N__29635\,
            in3 => \N__29599\,
            lcout => \c0.n70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_687_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__29625\,
            in1 => \N__29598\,
            in2 => \_gnd_net_\,
            in3 => \N__29568\,
            lcout => \c0.n19050\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_594_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29737\,
            in1 => \N__29470\,
            in2 => \N__29554\,
            in3 => \N__41506\,
            lcout => \c0.n63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_50_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29509\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \r_Rx_Data\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_511_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__42518\,
            in1 => \N__37960\,
            in2 => \N__29695\,
            in3 => \N__31543\,
            lcout => \c0.n18601\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_251_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29495\,
            in2 => \_gnd_net_\,
            in3 => \N__41435\,
            lcout => \c0.n18659\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i16_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29496\,
            in2 => \_gnd_net_\,
            in3 => \N__40545\,
            lcout => \c0.FRAME_MATCHER_state_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71077\,
            ce => 'H',
            sr => \N__29476\
        );

    \c0.i3_4_lut_adj_674_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31627\,
            in1 => \N__35472\,
            in2 => \N__31690\,
            in3 => \N__29450\,
            lcout => \c0.n19146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_858_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29451\,
            in2 => \_gnd_net_\,
            in3 => \N__41467\,
            lcout => \c0.n18633\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_680_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29824\,
            in1 => \N__29792\,
            in2 => \N__29694\,
            in3 => \N__29776\,
            lcout => \c0.n17_adj_3486\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_923_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41468\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31688\,
            lcout => \c0.n18681\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i7_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29729\,
            in2 => \_gnd_net_\,
            in3 => \N__40548\,
            lcout => \c0.FRAME_MATCHER_state_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71103\,
            ce => 'H',
            sr => \N__29707\
        );

    \c0.FRAME_MATCHER_state_i30_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40549\,
            in2 => \_gnd_net_\,
            in3 => \N__29687\,
            lcout => \c0.FRAME_MATCHER_state_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71117\,
            ce => 'H',
            sr => \N__29665\
        );

    \c0.FRAME_MATCHER_state_i4_LC_12_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40550\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31626\,
            lcout => \c0.FRAME_MATCHER_state_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71133\,
            ce => 'H',
            sr => \N__31606\
        );

    \c0.FRAME_MATCHER_i_i3_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111010101"
        )
    port map (
            in0 => \N__38670\,
            in1 => \N__60710\,
            in2 => \N__40084\,
            in3 => \N__31723\,
            lcout => \c0.FRAME_MATCHER_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71150\,
            ce => 'H',
            sr => \N__46937\
        );

    \c0.select_357_Select_2_i6_2_lut_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__60709\,
            in1 => \_gnd_net_\,
            in2 => \N__59944\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.n6_adj_3143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i2_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__38984\,
            in1 => \N__31594\,
            in2 => \N__29653\,
            in3 => \N__35437\,
            lcout => \c0.FRAME_MATCHER_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71150\,
            ce => 'H',
            sr => \N__46937\
        );

    \c0.i1_2_lut_3_lut_adj_675_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__59921\,
            in1 => \N__60048\,
            in2 => \_gnd_net_\,
            in3 => \N__40071\,
            lcout => \c0.n4_adj_3227\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_63_i9_2_lut_3_lut_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111111"
        )
    port map (
            in0 => \N__60049\,
            in1 => \_gnd_net_\,
            in2 => \N__60263\,
            in3 => \N__59923\,
            lcout => \c0.n9_adj_3351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_64_i9_2_lut_3_lut_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__59922\,
            in1 => \N__60242\,
            in2 => \_gnd_net_\,
            in3 => \N__60047\,
            lcout => \c0.n9_adj_3251\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i3_4_lut_adj_948_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29913\,
            in1 => \N__29884\,
            in2 => \N__29869\,
            in3 => \N__29920\,
            lcout => count_enable_adj_3586,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.A_delayed_67_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29866\,
            lcout => \quad_counter1.A_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71136\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.A_filtered_I_0_2_lut_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29883\,
            in2 => \_gnd_net_\,
            in3 => \N__29868\,
            lcout => \quad_counter1.count_direction\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.B_delayed_68_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29914\,
            lcout => \quad_counter1.B_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i1063_1_lut_2_lut_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29882\,
            in2 => \_gnd_net_\,
            in3 => \N__29867\,
            lcout => \quad_counter1.n2301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_1_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30498\,
            in2 => \N__30564\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \quad_counter1.n17314\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_2_lut_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29833\,
            in2 => \N__37212\,
            in3 => \N__29827\,
            lcout => n2345,
            ltout => OPEN,
            carryin => \quad_counter1.n17314\,
            carryout => \quad_counter1.n17315\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_3_lut_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30499\,
            in2 => \N__33702\,
            in3 => \N__30076\,
            lcout => n2344,
            ltout => OPEN,
            carryin => \quad_counter1.n17315\,
            carryout => \quad_counter1.n17316\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_4_lut_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30505\,
            in2 => \N__31090\,
            in3 => \N__30061\,
            lcout => n2343,
            ltout => OPEN,
            carryin => \quad_counter1.n17316\,
            carryout => \quad_counter1.n17317\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_5_lut_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30500\,
            in2 => \N__33037\,
            in3 => \N__30058\,
            lcout => n2342,
            ltout => OPEN,
            carryin => \quad_counter1.n17317\,
            carryout => \quad_counter1.n17318\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_6_lut_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30506\,
            in2 => \N__30919\,
            in3 => \N__30043\,
            lcout => n2341,
            ltout => OPEN,
            carryin => \quad_counter1.n17318\,
            carryout => \quad_counter1.n17319\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_7_lut_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30501\,
            in2 => \N__32853\,
            in3 => \N__30040\,
            lcout => n2340,
            ltout => OPEN,
            carryin => \quad_counter1.n17319\,
            carryout => \quad_counter1.n17320\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_8_lut_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30507\,
            in2 => \N__30037\,
            in3 => \N__29995\,
            lcout => n2339,
            ltout => OPEN,
            carryin => \quad_counter1.n17320\,
            carryout => \quad_counter1.n17321\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_9_lut_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30565\,
            in2 => \N__29992\,
            in3 => \N__29947\,
            lcout => n2338,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \quad_counter1.n17322\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_10_lut_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30569\,
            in2 => \N__36369\,
            in3 => \N__29932\,
            lcout => n2337,
            ltout => OPEN,
            carryin => \quad_counter1.n17322\,
            carryout => \quad_counter1.n17323\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_11_lut_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30566\,
            in2 => \N__31167\,
            in3 => \N__29923\,
            lcout => n2336,
            ltout => OPEN,
            carryin => \quad_counter1.n17323\,
            carryout => \quad_counter1.n17324\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_12_lut_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30570\,
            in2 => \N__30291\,
            in3 => \N__30262\,
            lcout => n2335,
            ltout => OPEN,
            carryin => \quad_counter1.n17324\,
            carryout => \quad_counter1.n17325\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_13_lut_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30567\,
            in2 => \N__30255\,
            in3 => \N__30226\,
            lcout => n2334,
            ltout => OPEN,
            carryin => \quad_counter1.n17325\,
            carryout => \quad_counter1.n17326\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_14_lut_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30571\,
            in2 => \N__37060\,
            in3 => \N__30223\,
            lcout => n2333,
            ltout => OPEN,
            carryin => \quad_counter1.n17326\,
            carryout => \quad_counter1.n17327\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_15_lut_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30568\,
            in2 => \N__30219\,
            in3 => \N__30190\,
            lcout => n2332,
            ltout => OPEN,
            carryin => \quad_counter1.n17327\,
            carryout => \quad_counter1.n17328\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_16_lut_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30572\,
            in2 => \N__30186\,
            in3 => \N__30157\,
            lcout => n2331,
            ltout => OPEN,
            carryin => \quad_counter1.n17328\,
            carryout => \quad_counter1.n17329\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_17_lut_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30573\,
            in2 => \N__30153\,
            in3 => \N__30124\,
            lcout => n2330,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \quad_counter1.n17330\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_18_lut_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30577\,
            in2 => \N__30117\,
            in3 => \N__30088\,
            lcout => n2329,
            ltout => OPEN,
            carryin => \quad_counter1.n17330\,
            carryout => \quad_counter1.n17331\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_19_lut_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30574\,
            in2 => \N__31056\,
            in3 => \N__30079\,
            lcout => n2328,
            ltout => OPEN,
            carryin => \quad_counter1.n17331\,
            carryout => \quad_counter1.n17332\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_20_lut_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30578\,
            in2 => \N__33294\,
            in3 => \N__30418\,
            lcout => n2327,
            ltout => OPEN,
            carryin => \quad_counter1.n17332\,
            carryout => \quad_counter1.n17333\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_21_lut_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30575\,
            in2 => \N__30415\,
            in3 => \N__30376\,
            lcout => n2326,
            ltout => OPEN,
            carryin => \quad_counter1.n17333\,
            carryout => \quad_counter1.n17334\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_22_lut_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30579\,
            in2 => \N__30372\,
            in3 => \N__30343\,
            lcout => n2325,
            ltout => OPEN,
            carryin => \quad_counter1.n17334\,
            carryout => \quad_counter1.n17335\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_23_lut_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30576\,
            in2 => \N__32965\,
            in3 => \N__30340\,
            lcout => n2324,
            ltout => OPEN,
            carryin => \quad_counter1.n17335\,
            carryout => \quad_counter1.n17336\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_24_lut_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30580\,
            in2 => \N__30337\,
            in3 => \N__30310\,
            lcout => n2323,
            ltout => OPEN,
            carryin => \quad_counter1.n17336\,
            carryout => \quad_counter1.n17337\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_25_lut_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30581\,
            in2 => \N__36322\,
            in3 => \N__30307\,
            lcout => n2322,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \quad_counter1.n17338\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_26_lut_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30752\,
            in2 => \N__30598\,
            in3 => \N__30298\,
            lcout => n2321,
            ltout => OPEN,
            carryin => \quad_counter1.n17338\,
            carryout => \quad_counter1.n17339\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_27_lut_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30585\,
            in2 => \N__31111\,
            in3 => \N__30295\,
            lcout => n2320,
            ltout => OPEN,
            carryin => \quad_counter1.n17339\,
            carryout => \quad_counter1.n17340\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_28_lut_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32798\,
            in2 => \N__30599\,
            in3 => \N__30688\,
            lcout => n2319,
            ltout => OPEN,
            carryin => \quad_counter1.n17340\,
            carryout => \quad_counter1.n17341\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_29_lut_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30589\,
            in2 => \N__30684\,
            in3 => \N__30655\,
            lcout => n2318,
            ltout => OPEN,
            carryin => \quad_counter1.n17341\,
            carryout => \quad_counter1.n17342\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_30_lut_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36078\,
            in2 => \N__30600\,
            in3 => \N__30652\,
            lcout => n2317,
            ltout => OPEN,
            carryin => \quad_counter1.n17342\,
            carryout => \quad_counter1.n17343\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_31_lut_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30593\,
            in2 => \N__33391\,
            in3 => \N__30649\,
            lcout => n2316,
            ltout => OPEN,
            carryin => \quad_counter1.n17343\,
            carryout => \quad_counter1.n17344\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_32_lut_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30642\,
            in2 => \N__30601\,
            in3 => \N__30604\,
            lcout => n2315,
            ltout => OPEN,
            carryin => \quad_counter1.n17344\,
            carryout => \quad_counter1.n17345\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_635_33_lut_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__30869\,
            in1 => \N__30597\,
            in2 => \_gnd_net_\,
            in3 => \N__30457\,
            lcout => n2314,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i31_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36229\,
            in1 => \N__30454\,
            in2 => \_gnd_net_\,
            in3 => \N__30870\,
            lcout => encoder1_position_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i0_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30448\,
            in1 => \N__36230\,
            in2 => \_gnd_net_\,
            in3 => \N__37211\,
            lcout => encoder1_position_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30970\,
            in1 => \N__30438\,
            in2 => \_gnd_net_\,
            in3 => \N__40884\,
            lcout => \c0.n11_adj_3462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__4__5330_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46724\,
            in1 => \N__30918\,
            in2 => \_gnd_net_\,
            in3 => \N__30885\,
            lcout => data_out_frame_13_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__7__5351_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30871\,
            in1 => \N__33231\,
            in2 => \_gnd_net_\,
            in3 => \N__46725\,
            lcout => data_out_frame_10_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i25_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36228\,
            in1 => \N__31109\,
            in2 => \_gnd_net_\,
            in3 => \N__30859\,
            lcout => encoder1_position_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i5_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__33799\,
            in1 => \N__33873\,
            in2 => \N__30852\,
            in3 => \N__37243\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71040\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17700_3_lut_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30832\,
            in1 => \N__30813\,
            in2 => \_gnd_net_\,
            in3 => \N__40885\,
            lcout => \c0.n21287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__1__5373_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46646\,
            in1 => \N__30786\,
            in2 => \_gnd_net_\,
            in3 => \N__31218\,
            lcout => data_out_frame_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71040\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__0__5358_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30763\,
            in1 => \N__33628\,
            in2 => \_gnd_net_\,
            in3 => \N__46648\,
            lcout => data_out_frame_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71040\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_0__4__5434_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__39493\,
            in1 => \N__30735\,
            in2 => \N__38996\,
            in3 => \N__37091\,
            lcout => \c0.data_out_frame_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71040\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__0__5374_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30713\,
            in1 => \N__33591\,
            in2 => \_gnd_net_\,
            in3 => \N__46650\,
            lcout => data_out_frame_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71040\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__0__5366_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46647\,
            in1 => \N__31144\,
            in2 => \_gnd_net_\,
            in3 => \N__33573\,
            lcout => data_out_frame_9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71040\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__1__5357_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31110\,
            in1 => \N__30994\,
            in2 => \_gnd_net_\,
            in3 => \N__46649\,
            lcout => data_out_frame_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71040\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__2__5332_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46651\,
            in2 => \N__31033\,
            in3 => \N__31086\,
            lcout => data_out_frame_13_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__1__5349_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__30981\,
            in1 => \N__31060\,
            in2 => \N__46765\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame_11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__40883\,
            in1 => \_gnd_net_\,
            in2 => \N__31032\,
            in3 => \N__31017\,
            lcout => \c0.n11_adj_3108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_18029_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__30993\,
            in1 => \N__40882\,
            in2 => \N__30982\,
            in3 => \N__36633\,
            lcout => \c0.n21605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i276_3_lut_4_lut_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111011"
        )
    port map (
            in0 => \N__30953\,
            in1 => \N__33507\,
            in2 => \N__31302\,
            in3 => \N__31272\,
            lcout => \c0.n700\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__5__5329_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__32857\,
            in1 => \N__30969\,
            in2 => \N__46766\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame_13_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18009_3_lut_4_lut_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30954\,
            in1 => \N__33508\,
            in2 => \N__31303\,
            in3 => \N__31273\,
            lcout => \c0.tx_transmit_N_2443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_264_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37412\,
            in1 => \N__36864\,
            in2 => \N__37335\,
            in3 => \N__34264\,
            lcout => \c0.n15842\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17978_4_lut_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__36624\,
            in1 => \N__31264\,
            in2 => \N__36926\,
            in3 => \N__33163\,
            lcout => \c0.n21566\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i0_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__33800\,
            in1 => \N__31201\,
            in2 => \N__33885\,
            in3 => \N__31252\,
            lcout => \c0.r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71021\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n21605_bdd_4_lut_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__31246\,
            in1 => \N__31228\,
            in2 => \N__31222\,
            in3 => \N__36622\,
            lcout => OPEN,
            ltout => \c0.n21608_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17974_4_lut_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__36623\,
            in1 => \N__36885\,
            in2 => \N__31204\,
            in3 => \N__31342\,
            lcout => \c0.n21562\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17959_2_lut_2_lut_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31200\,
            in2 => \_gnd_net_\,
            in3 => \N__34083\,
            lcout => \c0.n21466\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__1__5341_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31174\,
            in1 => \N__31351\,
            in2 => \_gnd_net_\,
            in3 => \N__46645\,
            lcout => data_out_frame_12_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71009\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__5__5393_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46644\,
            in1 => \N__36448\,
            in2 => \_gnd_net_\,
            in3 => \N__33735\,
            lcout => data_out_frame_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71009\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_3_lut_4_lut_adj_610_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__37312\,
            in1 => \N__31375\,
            in2 => \N__37443\,
            in3 => \N__35953\,
            lcout => OPEN,
            ltout => \n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i3_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__33861\,
            in1 => \N__31366\,
            in2 => \N__31369\,
            in3 => \N__33798\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71009\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33670\,
            in1 => \N__31350\,
            in2 => \_gnd_net_\,
            in3 => \N__40738\,
            lcout => \c0.n11_adj_3104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i2_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__31324\,
            in1 => \N__33797\,
            in2 => \N__33878\,
            in3 => \N__31336\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71009\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1399__i0_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31536\,
            in2 => \N__40825\,
            in3 => \_gnd_net_\,
            lcout => \c0.byte_transmit_counter_0\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \c0.n17346\,
            clk => \N__71022\,
            ce => \N__31408\,
            sr => \N__31393\
        );

    \c0.byte_transmit_counter_1399__i1_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36589\,
            in2 => \_gnd_net_\,
            in3 => \N__31312\,
            lcout => \c0.byte_transmit_counter_1\,
            ltout => OPEN,
            carryin => \c0.n17346\,
            carryout => \c0.n17347\,
            clk => \N__71022\,
            ce => \N__31408\,
            sr => \N__31393\
        );

    \c0.byte_transmit_counter_1399__i2_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36925\,
            in2 => \_gnd_net_\,
            in3 => \N__31309\,
            lcout => \c0.byte_transmit_counter_2\,
            ltout => OPEN,
            carryin => \c0.n17347\,
            carryout => \c0.n17348\,
            clk => \N__71022\,
            ce => \N__31408\,
            sr => \N__31393\
        );

    \c0.byte_transmit_counter_1399__i3_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37311\,
            in2 => \_gnd_net_\,
            in3 => \N__31306\,
            lcout => byte_transmit_counter_3,
            ltout => OPEN,
            carryin => \c0.n17348\,
            carryout => \c0.n17349\,
            clk => \N__71022\,
            ce => \N__31408\,
            sr => \N__31393\
        );

    \c0.byte_transmit_counter_1399__i4_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37408\,
            in2 => \_gnd_net_\,
            in3 => \N__31459\,
            lcout => byte_transmit_counter_4,
            ltout => OPEN,
            carryin => \c0.n17349\,
            carryout => \c0.n17350\,
            clk => \N__71022\,
            ce => \N__31408\,
            sr => \N__31393\
        );

    \c0.byte_transmit_counter_1399__i5_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33848\,
            in2 => \_gnd_net_\,
            in3 => \N__31456\,
            lcout => byte_transmit_counter_5,
            ltout => OPEN,
            carryin => \c0.n17350\,
            carryout => \c0.n17351\,
            clk => \N__71022\,
            ce => \N__31408\,
            sr => \N__31393\
        );

    \c0.byte_transmit_counter_1399__i6_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33540\,
            in2 => \_gnd_net_\,
            in3 => \N__31453\,
            lcout => \c0.byte_transmit_counter_6\,
            ltout => OPEN,
            carryin => \c0.n17351\,
            carryout => \c0.n17352\,
            clk => \N__71022\,
            ce => \N__31408\,
            sr => \N__31393\
        );

    \c0.byte_transmit_counter_1399__i7_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33522\,
            in2 => \_gnd_net_\,
            in3 => \N__31450\,
            lcout => \c0.byte_transmit_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71022\,
            ce => \N__31408\,
            sr => \N__31393\
        );

    \c0.i18005_4_lut_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__42512\,
            in1 => \N__31440\,
            in2 => \N__31428\,
            in3 => \N__31468\,
            lcout => \c0.n12326\,
            ltout => \c0.n12326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18001_2_lut_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__39595\,
            in1 => \_gnd_net_\,
            in2 => \N__31396\,
            in3 => \_gnd_net_\,
            lcout => \c0.n12758\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_741_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40092\,
            in1 => \N__40267\,
            in2 => \N__59965\,
            in3 => \N__38193\,
            lcout => OPEN,
            ltout => \c0.n4_adj_3263_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12196_4_lut_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001010000"
        )
    port map (
            in0 => \N__38153\,
            in1 => \N__60272\,
            in2 => \N__31381\,
            in3 => \N__60115\,
            lcout => \c0.n936\,
            ltout => \c0.n936_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_671_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__42516\,
            in1 => \_gnd_net_\,
            in2 => \N__31378\,
            in3 => \N__42330\,
            lcout => \c0.n10_adj_3081\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17902_4_lut_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010110000"
        )
    port map (
            in0 => \N__31537\,
            in1 => \N__39596\,
            in2 => \N__42520\,
            in3 => \N__38848\,
            lcout => \c0.n21420\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_18_i6_2_lut_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__60692\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38046\,
            lcout => \c0.n6_adj_3186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_313_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31507\,
            in2 => \_gnd_net_\,
            in3 => \N__41403\,
            lcout => \c0.n18627\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_13_i6_2_lut_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__60691\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34848\,
            lcout => \c0.n6_adj_3162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_949_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100010"
        )
    port map (
            in0 => \N__42506\,
            in1 => \N__39075\,
            in2 => \N__38977\,
            in3 => \N__35418\,
            lcout => n20764,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_20_i6_2_lut_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60694\,
            in2 => \_gnd_net_\,
            in3 => \N__34483\,
            lcout => \c0.n6_adj_3182\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_19_i6_2_lut_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34594\,
            in2 => \_gnd_net_\,
            in3 => \N__60693\,
            lcout => \c0.n6_adj_3184\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_21_i6_2_lut_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__60690\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35079\,
            lcout => \c0.n6_adj_3180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16066_2_lut_4_lut_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110010"
        )
    port map (
            in0 => \N__38925\,
            in1 => \N__38841\,
            in2 => \N__39597\,
            in3 => \N__39064\,
            lcout => \c0.n19650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__38380\,
            in1 => \N__35095\,
            in2 => \N__34729\,
            in3 => \N__38326\,
            lcout => \c0.n5_adj_2999\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_17_i6_2_lut_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60689\,
            in2 => \_gnd_net_\,
            in3 => \N__35055\,
            lcout => \c0.n6_adj_3188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16054_2_lut_3_lut_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__42508\,
            in1 => \N__31571\,
            in2 => \_gnd_net_\,
            in3 => \N__42323\,
            lcout => \c0.n19638\,
            ltout => \c0.n19638_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17686_3_lut_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__38362\,
            in1 => \_gnd_net_\,
            in2 => \N__31588\,
            in3 => \N__34757\,
            lcout => \c0.n21273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_583_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__38247\,
            in1 => \N__38927\,
            in2 => \N__42519\,
            in3 => \N__39594\,
            lcout => \c0.n11432\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_877_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__42479\,
            in1 => \N__38926\,
            in2 => \N__39598\,
            in3 => \N__38246\,
            lcout => \c0.n63_adj_3146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_390_Select_2_i6_3_lut_4_lut_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__42324\,
            in1 => \N__34727\,
            in2 => \N__42507\,
            in3 => \N__35209\,
            lcout => OPEN,
            ltout => \c0.n6_adj_3521_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i2_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__34758\,
            in1 => \N__31585\,
            in2 => \N__31579\,
            in3 => \N__31696\,
            lcout => \FRAME_MATCHER_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71065\,
            ce => 'H',
            sr => \N__46738\
        );

    \c0.i1_3_lut_4_lut_adj_913_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__42329\,
            in1 => \N__38284\,
            in2 => \N__31576\,
            in3 => \N__38321\,
            lcout => \c0.n11_adj_3370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_254_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31662\,
            in2 => \_gnd_net_\,
            in3 => \N__41434\,
            lcout => \c0.n18657\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_797_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__35155\,
            in1 => \N__34951\,
            in2 => \N__35134\,
            in3 => \N__35207\,
            lcout => OPEN,
            ltout => \c0.n6_adj_3515_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_753_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__38476\,
            in1 => \N__31708\,
            in2 => \N__31699\,
            in3 => \N__38524\,
            lcout => \c0.n5_adj_3516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i29_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40490\,
            in2 => \_gnd_net_\,
            in3 => \N__34931\,
            lcout => \c0.FRAME_MATCHER_state_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71089\,
            ce => 'H',
            sr => \N__35218\
        );

    \c0.FRAME_MATCHER_state_i5_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31689\,
            in2 => \_gnd_net_\,
            in3 => \N__40515\,
            lcout => \c0.FRAME_MATCHER_state_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71105\,
            ce => 'H',
            sr => \N__31672\
        );

    \c0.FRAME_MATCHER_state_i17_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40546\,
            in2 => \_gnd_net_\,
            in3 => \N__31658\,
            lcout => \c0.FRAME_MATCHER_state_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71119\,
            ce => 'H',
            sr => \N__31636\
        );

    \c0.FRAME_MATCHER_state_i8_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35471\,
            in2 => \_gnd_net_\,
            in3 => \N__40547\,
            lcout => \c0.FRAME_MATCHER_state_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71135\,
            ce => 'H',
            sr => \N__35449\
        );

    \c0.i1_2_lut_adj_860_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31625\,
            in2 => \_gnd_net_\,
            in3 => \N__41466\,
            lcout => \c0.n18629\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_2_lut_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42170\,
            in1 => \N__60208\,
            in2 => \N__41829\,
            in3 => \_gnd_net_\,
            lcout => n16,
            ltout => OPEN,
            carryin => \bfn_14_5_0_\,
            carryout => \c0.n17176\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i1_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42196\,
            in1 => \N__60041\,
            in2 => \_gnd_net_\,
            in3 => \N__31597\,
            lcout => \c0.FRAME_MATCHER_i_1\,
            ltout => OPEN,
            carryin => \c0.n17176\,
            carryout => \c0.n17177\,
            clk => \N__71177\,
            ce => 'H',
            sr => \N__60511\
        );

    \c0.add_80_4_lut_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42171\,
            in1 => \N__59927\,
            in2 => \_gnd_net_\,
            in3 => \N__31726\,
            lcout => \c0.n2_adj_3144\,
            ltout => OPEN,
            carryin => \c0.n17177\,
            carryout => \c0.n17178\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_5_lut_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42195\,
            in1 => \N__40062\,
            in2 => \_gnd_net_\,
            in3 => \N__31717\,
            lcout => \c0.n2_adj_3145\,
            ltout => OPEN,
            carryin => \c0.n17178\,
            carryout => \c0.n17179\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_6_lut_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42169\,
            in1 => \N__40266\,
            in2 => \_gnd_net_\,
            in3 => \N__31714\,
            lcout => \c0.n2_adj_3147\,
            ltout => OPEN,
            carryin => \c0.n17179\,
            carryout => \c0.n17180\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_6_THRU_CRY_0_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32614\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17180\,
            carryout => \c0.n17180_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_6_THRU_CRY_1_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32704\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17180_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17180_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_6_THRU_CRY_2_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32618\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17180_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17180_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i5_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42197\,
            in1 => \N__49618\,
            in2 => \_gnd_net_\,
            in3 => \N__31711\,
            lcout => \c0.FRAME_MATCHER_i_5\,
            ltout => OPEN,
            carryin => \bfn_14_6_0_\,
            carryout => \c0.n17181\,
            clk => \N__71165\,
            ce => 'H',
            sr => \N__49597\
        );

    \c0.add_80_7_THRU_CRY_0_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32601\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17181\,
            carryout => \c0.n17181_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_7_THRU_CRY_1_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32701\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17181_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17181_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_7_THRU_CRY_2_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32605\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17181_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17181_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_7_THRU_CRY_3_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32702\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17181_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17181_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_7_THRU_CRY_4_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32609\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17181_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17181_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_7_THRU_CRY_5_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32703\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17181_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17181_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_7_THRU_CRY_6_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32613\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17181_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17181_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i6_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42200\,
            in1 => \N__40164\,
            in2 => \_gnd_net_\,
            in3 => \N__31729\,
            lcout => \c0.FRAME_MATCHER_i_6\,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \c0.n17182\,
            clk => \N__71152\,
            ce => 'H',
            sr => \N__35803\
        );

    \c0.add_80_8_THRU_CRY_0_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32588\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17182\,
            carryout => \c0.n17182_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_8_THRU_CRY_1_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32698\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17182_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17182_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_8_THRU_CRY_2_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32592\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17182_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17182_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_8_THRU_CRY_3_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32699\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17182_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17182_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_8_THRU_CRY_4_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32596\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17182_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17182_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_8_THRU_CRY_5_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32700\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17182_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17182_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_8_THRU_CRY_6_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32600\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17182_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17182_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i7_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42199\,
            in1 => \N__34424\,
            in2 => \_gnd_net_\,
            in3 => \N__31732\,
            lcout => \c0.FRAME_MATCHER_i_7\,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \c0.n17183\,
            clk => \N__71138\,
            ce => 'H',
            sr => \N__33481\
        );

    \c0.add_80_9_THRU_CRY_0_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32566\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17183\,
            carryout => \c0.n17183_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_9_THRU_CRY_1_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32695\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17183_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17183_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_9_THRU_CRY_2_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32570\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17183_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17183_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_9_THRU_CRY_3_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32696\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17183_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17183_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_9_THRU_CRY_4_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32574\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17183_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17183_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_9_THRU_CRY_5_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32697\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17183_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17183_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_9_THRU_CRY_6_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32578\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17183_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17183_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i8_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42198\,
            in1 => \N__34610\,
            in2 => \_gnd_net_\,
            in3 => \N__31735\,
            lcout => \c0.FRAME_MATCHER_i_8\,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \c0.n17184\,
            clk => \N__71122\,
            ce => 'H',
            sr => \N__32773\
        );

    \c0.add_80_10_THRU_CRY_0_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32408\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17184\,
            carryout => \c0.n17184_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_10_THRU_CRY_1_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32585\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17184_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17184_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_10_THRU_CRY_2_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32412\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17184_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17184_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_10_THRU_CRY_3_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32586\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17184_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17184_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_10_THRU_CRY_4_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32416\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17184_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17184_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_10_THRU_CRY_5_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32587\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17184_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17184_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_10_THRU_CRY_6_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32420\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17184_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17184_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i9_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42224\,
            in1 => \N__34802\,
            in2 => \_gnd_net_\,
            in3 => \N__31738\,
            lcout => \c0.FRAME_MATCHER_i_9\,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => \c0.n17185\,
            clk => \N__71106\,
            ce => 'H',
            sr => \N__31885\
        );

    \c0.add_80_11_THRU_CRY_0_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32395\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17185\,
            carryout => \c0.n17185_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_11_THRU_CRY_1_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32582\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17185_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17185_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_11_THRU_CRY_2_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32399\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17185_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17185_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_11_THRU_CRY_3_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32583\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17185_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17185_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_11_THRU_CRY_4_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32403\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17185_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17185_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_11_THRU_CRY_5_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32584\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17185_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17185_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_11_THRU_CRY_6_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32407\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17185_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17185_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i10_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42227\,
            in1 => \N__34892\,
            in2 => \_gnd_net_\,
            in3 => \N__31744\,
            lcout => \c0.FRAME_MATCHER_i_10\,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => \c0.n17186\,
            clk => \N__71090\,
            ce => 'H',
            sr => \N__33400\
        );

    \c0.add_80_12_THRU_CRY_0_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32382\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17186\,
            carryout => \c0.n17186_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_12_THRU_CRY_1_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32579\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17186_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17186_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_12_THRU_CRY_2_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32386\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17186_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17186_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_12_THRU_CRY_3_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32580\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17186_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17186_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_12_THRU_CRY_4_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32390\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17186_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17186_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_12_THRU_CRY_5_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32581\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17186_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17186_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_12_THRU_CRY_6_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32394\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17186_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17186_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i11_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42226\,
            in1 => \N__34323\,
            in2 => \_gnd_net_\,
            in3 => \N__31741\,
            lcout => \c0.FRAME_MATCHER_i_11\,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \c0.n17187\,
            clk => \N__71078\,
            ce => 'H',
            sr => \N__34405\
        );

    \c0.add_80_13_THRU_CRY_0_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32348\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17187\,
            carryout => \c0.n17187_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_13_THRU_CRY_1_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32563\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17187_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17187_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_13_THRU_CRY_2_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32352\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17187_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17187_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_13_THRU_CRY_3_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32564\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17187_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17187_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_13_THRU_CRY_4_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32356\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17187_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17187_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_13_THRU_CRY_5_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32565\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17187_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17187_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_13_THRU_CRY_6_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32360\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17187_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17187_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i12_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42225\,
            in1 => \N__34497\,
            in2 => \_gnd_net_\,
            in3 => \N__31747\,
            lcout => \c0.FRAME_MATCHER_i_12\,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \c0.n17188\,
            clk => \N__71066\,
            ce => 'H',
            sr => \N__34573\
        );

    \c0.add_80_14_THRU_CRY_0_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32193\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17188\,
            carryout => \c0.n17188_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_14_THRU_CRY_1_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32379\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17188_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17188_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_14_THRU_CRY_2_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32197\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17188_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17188_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_14_THRU_CRY_3_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32380\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17188_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17188_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_14_THRU_CRY_4_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32201\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17188_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17188_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_14_THRU_CRY_5_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32381\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17188_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17188_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_14_THRU_CRY_6_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32205\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17188_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17188_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i13_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42249\,
            in1 => \N__34835\,
            in2 => \_gnd_net_\,
            in3 => \N__31762\,
            lcout => \c0.FRAME_MATCHER_i_13\,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \c0.n17189\,
            clk => \N__71053\,
            ce => 'H',
            sr => \N__31759\
        );

    \c0.add_80_15_THRU_CRY_0_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32180\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17189\,
            carryout => \c0.n17189_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_15_THRU_CRY_1_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32376\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17189_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17189_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_15_THRU_CRY_2_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32184\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17189_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17189_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_15_THRU_CRY_3_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32377\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17189_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17189_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_15_THRU_CRY_4_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32188\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17189_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17189_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_15_THRU_CRY_5_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32378\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17189_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17189_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_15_THRU_CRY_6_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32192\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17189_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17189_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i14_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42252\,
            in1 => \N__34455\,
            in2 => \_gnd_net_\,
            in3 => \N__31765\,
            lcout => \c0.FRAME_MATCHER_i_14\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \c0.n17190\,
            clk => \N__71041\,
            ce => 'H',
            sr => \N__34522\
        );

    \c0.add_80_16_THRU_CRY_0_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32000\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17190\,
            carryout => \c0.n17190_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_16_THRU_CRY_1_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32071\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17190_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17190_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_16_THRU_CRY_2_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32004\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17190_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17190_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_16_THRU_CRY_3_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32072\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17190_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17190_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_16_THRU_CRY_4_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32008\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17190_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17190_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_16_THRU_CRY_5_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__32073\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17190_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17190_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_16_THRU_CRY_6_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32012\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17190_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17190_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i15_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42251\,
            in1 => \N__34868\,
            in2 => \_gnd_net_\,
            in3 => \N__31768\,
            lcout => \c0.FRAME_MATCHER_i_15\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \c0.n17191\,
            clk => \N__71032\,
            ce => 'H',
            sr => \N__33712\
        );

    \c0.add_80_17_THRU_CRY_0_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31993\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17191\,
            carryout => \c0.n17191_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_17_THRU_CRY_1_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31997\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17191_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17191_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_17_THRU_CRY_2_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31994\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17191_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17191_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_17_THRU_CRY_3_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31998\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17191_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17191_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_17_THRU_CRY_4_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31995\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17191_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17191_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_17_THRU_CRY_5_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31999\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17191_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17191_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_17_THRU_CRY_6_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31996\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17191_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17191_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i16_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42250\,
            in1 => \N__34355\,
            in2 => \_gnd_net_\,
            in3 => \N__31771\,
            lcout => \c0.FRAME_MATCHER_i_16\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \c0.n17192\,
            clk => \N__71015\,
            ce => 'H',
            sr => \N__33655\
        );

    \c0.add_80_18_THRU_CRY_0_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32013\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17192\,
            carryout => \c0.n17192_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_18_THRU_CRY_1_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32017\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17192_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17192_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_18_THRU_CRY_2_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32014\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17192_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17192_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_18_THRU_CRY_3_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32018\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17192_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17192_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_18_THRU_CRY_4_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32015\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17192_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17192_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_18_THRU_CRY_5_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32019\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17192_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17192_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_18_THRU_CRY_6_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32016\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17192_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17192_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i17_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42265\,
            in1 => \N__35042\,
            in2 => \_gnd_net_\,
            in3 => \N__31786\,
            lcout => \c0.FRAME_MATCHER_i_17\,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \c0.n17193\,
            clk => \N__71033\,
            ce => 'H',
            sr => \N__31783\
        );

    \c0.add_80_19_THRU_CRY_0_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32148\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17193\,
            carryout => \c0.n17193_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_19_THRU_CRY_1_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32152\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17193_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17193_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_19_THRU_CRY_2_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32149\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17193_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17193_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_19_THRU_CRY_3_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32153\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17193_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17193_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_19_THRU_CRY_4_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32150\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17193_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17193_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_19_THRU_CRY_5_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32154\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17193_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17193_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_19_THRU_CRY_6_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32151\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17193_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17193_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i18_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42266\,
            in1 => \N__38045\,
            in2 => \_gnd_net_\,
            in3 => \N__31798\,
            lcout => \c0.FRAME_MATCHER_i_18\,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \c0.n17194\,
            clk => \N__71042\,
            ce => 'H',
            sr => \N__31795\
        );

    \c0.add_80_20_THRU_CRY_0_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32155\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17194\,
            carryout => \c0.n17194_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_20_THRU_CRY_1_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32159\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17194_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17194_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_20_THRU_CRY_2_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32156\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17194_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17194_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_20_THRU_CRY_3_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32160\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17194_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17194_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_20_THRU_CRY_4_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32157\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17194_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17194_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_20_THRU_CRY_5_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32161\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17194_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17194_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_20_THRU_CRY_6_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32158\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17194_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17194_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i19_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42268\,
            in1 => \N__34589\,
            in2 => \_gnd_net_\,
            in3 => \N__31816\,
            lcout => \c0.FRAME_MATCHER_i_19\,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \c0.n17195\,
            clk => \N__71054\,
            ce => 'H',
            sr => \N__31813\
        );

    \c0.add_80_21_THRU_CRY_0_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32258\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17195\,
            carryout => \c0.n17195_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_21_THRU_CRY_1_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32262\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17195_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17195_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_21_THRU_CRY_2_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32259\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17195_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17195_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_21_THRU_CRY_3_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32263\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17195_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17195_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_21_THRU_CRY_4_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32260\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17195_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17195_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_21_THRU_CRY_5_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32264\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17195_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17195_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_21_THRU_CRY_6_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32261\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17195_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17195_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i20_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42267\,
            in1 => \N__34482\,
            in2 => \_gnd_net_\,
            in3 => \N__31801\,
            lcout => \c0.FRAME_MATCHER_i_20\,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \c0.n17196\,
            clk => \N__71067\,
            ce => 'H',
            sr => \N__31834\
        );

    \c0.add_80_22_THRU_CRY_0_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32458\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17196\,
            carryout => \c0.n17196_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_22_THRU_CRY_1_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32462\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17196_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17196_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_22_THRU_CRY_2_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32459\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17196_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17196_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_22_THRU_CRY_3_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32463\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17196_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17196_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_22_THRU_CRY_4_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32460\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17196_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17196_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_22_THRU_CRY_5_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32464\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17196_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17196_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_22_THRU_CRY_6_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32461\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17196_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17196_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i21_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42140\,
            in1 => \N__35078\,
            in2 => \_gnd_net_\,
            in3 => \N__31828\,
            lcout => \c0.FRAME_MATCHER_i_21\,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => \c0.n17197\,
            clk => \N__71079\,
            ce => 'H',
            sr => \N__31825\
        );

    \c0.add_80_23_THRU_CRY_0_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32465\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17197\,
            carryout => \c0.n17197_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_23_THRU_CRY_1_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32469\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17197_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17197_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_23_THRU_CRY_2_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32466\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17197_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17197_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_23_THRU_CRY_3_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32470\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17197_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17197_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_23_THRU_CRY_4_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32467\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17197_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17197_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_23_THRU_CRY_5_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32471\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17197_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17197_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_23_THRU_CRY_6_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32468\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17197_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17197_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i22_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42145\,
            in1 => \N__34382\,
            in2 => \_gnd_net_\,
            in3 => \N__31849\,
            lcout => \c0.FRAME_MATCHER_i_22\,
            ltout => OPEN,
            carryin => \bfn_14_23_0_\,
            carryout => \c0.n17198\,
            clk => \N__71091\,
            ce => 'H',
            sr => \N__31846\
        );

    \c0.add_80_24_THRU_CRY_0_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32472\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17198\,
            carryout => \c0.n17198_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_24_THRU_CRY_1_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32476\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17198_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17198_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_24_THRU_CRY_2_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32473\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17198_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17198_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_24_THRU_CRY_3_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32477\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17198_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17198_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_24_THRU_CRY_4_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32474\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17198_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17198_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_24_THRU_CRY_5_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32478\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17198_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17198_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_24_THRU_CRY_6_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32475\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17198_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17198_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i23_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42141\,
            in1 => \N__38018\,
            in2 => \_gnd_net_\,
            in3 => \N__31852\,
            lcout => \c0.FRAME_MATCHER_i_23\,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => \c0.n17199\,
            clk => \N__71107\,
            ce => 'H',
            sr => \N__35164\
        );

    \c0.add_80_25_THRU_CRY_0_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32479\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17199\,
            carryout => \c0.n17199_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_25_THRU_CRY_1_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32483\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17199_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17199_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_25_THRU_CRY_2_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32480\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17199_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17199_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_25_THRU_CRY_3_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32484\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17199_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17199_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_25_THRU_CRY_4_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32481\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17199_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17199_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_25_THRU_CRY_5_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32485\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17199_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17199_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_25_THRU_CRY_6_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32482\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17199_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17199_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i24_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42127\,
            in1 => \N__35013\,
            in2 => \_gnd_net_\,
            in3 => \N__31855\,
            lcout => \c0.FRAME_MATCHER_i_24\,
            ltout => OPEN,
            carryin => \bfn_14_25_0_\,
            carryout => \c0.n17200\,
            clk => \N__71121\,
            ce => 'H',
            sr => \N__34996\
        );

    \c0.add_80_26_THRU_CRY_0_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32619\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17200\,
            carryout => \c0.n17200_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_26_THRU_CRY_1_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32623\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17200_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17200_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_26_THRU_CRY_2_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32620\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17200_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17200_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_26_THRU_CRY_3_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32624\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17200_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17200_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_26_THRU_CRY_4_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32621\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17200_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17200_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_26_THRU_CRY_5_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32625\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17200_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17200_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_26_THRU_CRY_6_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32622\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17200_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17200_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i25_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42142\,
            in1 => \N__34551\,
            in2 => \_gnd_net_\,
            in3 => \N__31858\,
            lcout => \c0.FRAME_MATCHER_i_25\,
            ltout => OPEN,
            carryin => \bfn_14_26_0_\,
            carryout => \c0.n17201\,
            clk => \N__71137\,
            ce => 'H',
            sr => \N__34537\
        );

    \c0.add_80_27_THRU_CRY_0_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32626\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17201\,
            carryout => \c0.n17201_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_27_THRU_CRY_1_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32630\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17201_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17201_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_27_THRU_CRY_2_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32627\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17201_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17201_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_27_THRU_CRY_3_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32631\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17201_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17201_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_27_THRU_CRY_4_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32628\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17201_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17201_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_27_THRU_CRY_5_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32632\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17201_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17201_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_27_THRU_CRY_6_LC_14_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32629\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17201_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17201_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i26_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42143\,
            in1 => \N__35375\,
            in2 => \_gnd_net_\,
            in3 => \N__31861\,
            lcout => \c0.FRAME_MATCHER_i_26\,
            ltout => OPEN,
            carryin => \bfn_14_27_0_\,
            carryout => \c0.n17202\,
            clk => \N__71151\,
            ce => 'H',
            sr => \N__35353\
        );

    \c0.add_80_28_THRU_CRY_0_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32633\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17202\,
            carryout => \c0.n17202_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_28_THRU_CRY_1_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32637\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17202_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17202_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_28_THRU_CRY_2_LC_14_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32634\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17202_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17202_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_28_THRU_CRY_3_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32638\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17202_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17202_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_28_THRU_CRY_4_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32635\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17202_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17202_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_28_THRU_CRY_5_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32639\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17202_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17202_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_28_THRU_CRY_6_LC_14_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32636\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17202_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17202_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i27_LC_14_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42125\,
            in1 => \N__35327\,
            in2 => \_gnd_net_\,
            in3 => \N__31864\,
            lcout => \c0.FRAME_MATCHER_i_27\,
            ltout => OPEN,
            carryin => \bfn_14_28_0_\,
            carryout => \c0.n17203\,
            clk => \N__71164\,
            ce => 'H',
            sr => \N__35308\
        );

    \c0.add_80_29_THRU_CRY_0_LC_14_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32640\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17203\,
            carryout => \c0.n17203_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_29_THRU_CRY_1_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32644\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17203_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17203_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_29_THRU_CRY_2_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32641\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17203_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17203_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_29_THRU_CRY_3_LC_14_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32645\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17203_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17203_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_29_THRU_CRY_4_LC_14_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32642\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17203_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17203_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_29_THRU_CRY_5_LC_14_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32646\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17203_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17203_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_29_THRU_CRY_6_LC_14_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32643\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17203_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17203_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i28_LC_14_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42126\,
            in1 => \N__35291\,
            in2 => \_gnd_net_\,
            in3 => \N__31870\,
            lcout => \c0.FRAME_MATCHER_i_28\,
            ltout => OPEN,
            carryin => \bfn_14_29_0_\,
            carryout => \c0.n17204\,
            clk => \N__71176\,
            ce => 'H',
            sr => \N__35272\
        );

    \c0.add_80_30_THRU_CRY_0_LC_14_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32705\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17204\,
            carryout => \c0.n17204_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_30_THRU_CRY_1_LC_14_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32709\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17204_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17204_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_30_THRU_CRY_2_LC_14_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32706\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17204_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17204_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_30_THRU_CRY_3_LC_14_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32710\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17204_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17204_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_30_THRU_CRY_4_LC_14_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32707\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17204_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17204_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_30_THRU_CRY_5_LC_14_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32711\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17204_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17204_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_30_THRU_CRY_6_LC_14_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32708\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17204_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17204_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i29_LC_14_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42131\,
            in1 => \N__37985\,
            in2 => \_gnd_net_\,
            in3 => \N__31867\,
            lcout => \c0.FRAME_MATCHER_i_29\,
            ltout => OPEN,
            carryin => \bfn_14_30_0_\,
            carryout => \c0.n17205\,
            clk => \N__71188\,
            ce => 'H',
            sr => \N__35344\
        );

    \c0.add_80_31_THRU_CRY_0_LC_14_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32712\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17205\,
            carryout => \c0.n17205_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_31_THRU_CRY_1_LC_14_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32716\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17205_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17205_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_31_THRU_CRY_2_LC_14_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32713\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17205_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17205_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_31_THRU_CRY_3_LC_14_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32717\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17205_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17205_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_31_THRU_CRY_4_LC_14_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32714\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17205_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17205_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_31_THRU_CRY_5_LC_14_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32718\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17205_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17205_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_31_THRU_CRY_6_LC_14_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32715\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17205_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17205_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i30_LC_14_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42121\,
            in1 => \N__35246\,
            in2 => \_gnd_net_\,
            in3 => \N__31873\,
            lcout => \c0.FRAME_MATCHER_i_30\,
            ltout => OPEN,
            carryin => \bfn_14_31_0_\,
            carryout => \c0.n17206\,
            clk => \N__71199\,
            ce => 'H',
            sr => \N__35227\
        );

    \c0.add_80_32_THRU_CRY_0_LC_14_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32719\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17206\,
            carryout => \c0.n17206_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_32_THRU_CRY_1_LC_14_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32723\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17206_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n17206_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_32_THRU_CRY_2_LC_14_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32720\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17206_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n17206_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_32_THRU_CRY_3_LC_14_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32724\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17206_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n17206_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_32_THRU_CRY_4_LC_14_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32721\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17206_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n17206_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_32_THRU_CRY_5_LC_14_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32725\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17206_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n17206_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_80_32_THRU_CRY_6_LC_14_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32722\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n17206_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n17206_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i31_LC_14_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42144\,
            in1 => \N__38135\,
            in2 => \_gnd_net_\,
            in3 => \N__31915\,
            lcout => \c0.FRAME_MATCHER_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71212\,
            ce => 'H',
            sr => \N__35263\
        );

    \c0.FRAME_MATCHER_i_i0_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__60652\,
            in1 => \N__31912\,
            in2 => \N__60235\,
            in3 => \N__31897\,
            lcout => \FRAME_MATCHER_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71154\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_9_i6_2_lut_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34809\,
            in2 => \_gnd_net_\,
            in3 => \N__60651\,
            lcout => \c0.n6_adj_3155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__5__5345_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32964\,
            in1 => \N__33141\,
            in2 => \_gnd_net_\,
            in3 => \N__46692\,
            lcout => data_out_frame_11_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71154\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__0__5390_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46691\,
            in1 => \N__32896\,
            in2 => \_gnd_net_\,
            in3 => \N__32763\,
            lcout => data_out_frame_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71154\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i5_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36254\,
            in1 => \N__32843\,
            in2 => \_gnd_net_\,
            in3 => \N__32866\,
            lcout => encoder1_position_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71139\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__32781\,
            in1 => \N__40924\,
            in2 => \N__33646\,
            in3 => \N__36758\,
            lcout => \c0.n21647\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__2__5356_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32806\,
            in1 => \N__32782\,
            in2 => \_gnd_net_\,
            in3 => \N__46914\,
            lcout => data_out_frame_10_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71139\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_8_i6_2_lut_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60650\,
            in2 => \_gnd_net_\,
            in3 => \N__34614\,
            lcout => \c0.n6_adj_3154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__5__5209_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110010101010"
        )
    port map (
            in0 => \N__37488\,
            in1 => \N__62180\,
            in2 => \N__54479\,
            in3 => \N__46915\,
            lcout => data_out_frame_28_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71139\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13745_4_lut_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000001100"
        )
    port map (
            in0 => \N__32764\,
            in1 => \N__40925\,
            in2 => \N__36987\,
            in3 => \N__36755\,
            lcout => \c0.n6_adj_3321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i1_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__33689\,
            in1 => \N__36226\,
            in2 => \_gnd_net_\,
            in3 => \N__32737\,
            lcout => encoder1_position_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__4__5210_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__46860\,
            in1 => \N__62182\,
            in2 => \N__61132\,
            in3 => \N__33063\,
            lcout => data_out_frame_28_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_210_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__37231\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39352\,
            lcout => n11461,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i3_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36225\,
            in1 => \N__33023\,
            in2 => \_gnd_net_\,
            in3 => \N__33049\,
            lcout => encoder1_position_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__3__5379_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33004\,
            in1 => \N__35515\,
            in2 => \_gnd_net_\,
            in3 => \N__46799\,
            lcout => data_out_frame_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101000100"
        )
    port map (
            in0 => \N__36966\,
            in1 => \N__33439\,
            in2 => \N__33088\,
            in3 => \N__40904\,
            lcout => OPEN,
            ltout => \c0.n6_adj_3379_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17727_4_lut_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__36731\,
            in1 => \N__35485\,
            in2 => \N__32980\,
            in3 => \N__36967\,
            lcout => \c0.n21314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i21_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36249\,
            in1 => \N__32977\,
            in2 => \_gnd_net_\,
            in3 => \N__32957\,
            lcout => encoder1_position_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i45_2_lut_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52996\,
            in2 => \_gnd_net_\,
            in3 => \N__38786\,
            lcout => \c0.n160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17733_4_lut_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__32938\,
            in1 => \N__32923\,
            in2 => \N__36757\,
            in3 => \N__36968\,
            lcout => \c0.n21320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i23_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36250\,
            in1 => \N__36311\,
            in2 => \_gnd_net_\,
            in3 => \N__32911\,
            lcout => encoder1_position_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_52_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__37810\,
            in1 => \N__37870\,
            in2 => \N__53036\,
            in3 => \N__34273\,
            lcout => rx_data_ready,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__3__5371_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__46796\,
            in1 => \_gnd_net_\,
            in2 => \N__33178\,
            in3 => \N__33265\,
            lcout => data_out_frame_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_18039_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__36723\,
            in1 => \N__33235\,
            in2 => \N__36292\,
            in3 => \N__40908\,
            lcout => \c0.n21623\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n21641_bdd_4_lut_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__33205\,
            in1 => \N__33190\,
            in2 => \N__33177\,
            in3 => \N__36726\,
            lcout => \c0.n21644\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_rx_data_ready_prev_5165_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53011\,
            lcout => \c0.FRAME_MATCHER_rx_data_ready_prev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_18049_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__40907\,
            in1 => \N__33366\,
            in2 => \N__33148\,
            in3 => \N__36724\,
            lcout => OPEN,
            ltout => \c0.n21635_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n21635_bdd_4_lut_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__36725\,
            in1 => \N__33127\,
            in2 => \N__33112\,
            in3 => \N__33109\,
            lcout => \c0.n21638\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__3__5395_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46795\,
            in1 => \N__38740\,
            in2 => \_gnd_net_\,
            in3 => \N__33087\,
            lcout => data_out_frame_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__3__5211_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011001100"
        )
    port map (
            in0 => \N__61131\,
            in1 => \N__36019\,
            in2 => \N__56860\,
            in3 => \N__46798\,
            lcout => \c0.data_out_frame_28_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17910_2_lut_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35814\,
            in2 => \_gnd_net_\,
            in3 => \N__36736\,
            lcout => \c0.n21470\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i179_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__68612\,
            in1 => \N__67526\,
            in2 => \_gnd_net_\,
            in3 => \N__58871\,
            lcout => data_in_frame_22_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17955_3_lut_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__36048\,
            in1 => \N__36976\,
            in2 => \_gnd_net_\,
            in3 => \N__40900\,
            lcout => \c0.n21542\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i29_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36227\,
            in1 => \N__33383\,
            in2 => \_gnd_net_\,
            in3 => \N__33412\,
            lcout => encoder1_position_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_10_i6_2_lut_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34896\,
            in2 => \_gnd_net_\,
            in3 => \N__60688\,
            lcout => \c0.n6_adj_3156\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__5__5353_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33367\,
            in1 => \N__33384\,
            in2 => \_gnd_net_\,
            in3 => \N__46797\,
            lcout => data_out_frame_10_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__5__5385_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46779\,
            in1 => \N__33355\,
            in2 => \_gnd_net_\,
            in3 => \N__33906\,
            lcout => data_out_frame_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71068\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13744_3_lut_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36727\,
            in1 => \N__33325\,
            in2 => \_gnd_net_\,
            in3 => \N__36459\,
            lcout => \c0.n17150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__2__5348_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33295\,
            in1 => \N__33642\,
            in2 => \_gnd_net_\,
            in3 => \N__46780\,
            lcout => data_out_frame_11_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71068\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_18034_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__33627\,
            in1 => \N__40893\,
            in2 => \N__33613\,
            in3 => \N__36728\,
            lcout => OPEN,
            ltout => \c0.n21617_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n21617_bdd_4_lut_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__36729\,
            in1 => \N__33592\,
            in2 => \N__33577\,
            in3 => \N__33574\,
            lcout => OPEN,
            ltout => \c0.n21620_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17986_4_lut_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__36376\,
            in1 => \N__36950\,
            in2 => \N__33559\,
            in3 => \N__36730\,
            lcout => \c0.n21574\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_271_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__33879\,
            in1 => \N__33544\,
            in2 => \_gnd_net_\,
            in3 => \N__33526\,
            lcout => \c0.n7235\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i4_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110111011101"
        )
    port map (
            in0 => \N__38674\,
            in1 => \N__33496\,
            in2 => \N__40265\,
            in3 => \N__60687\,
            lcout => \c0.FRAME_MATCHER_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71055\,
            ce => 'H',
            sr => \N__46729\
        );

    \c0.select_357_Select_7_i6_2_lut_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60686\,
            in2 => \_gnd_net_\,
            in3 => \N__34441\,
            lcout => \c0.n6_adj_3151\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17721_4_lut_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__36696\,
            in1 => \N__36959\,
            in2 => \N__33721\,
            in3 => \N__33892\,
            lcout => \c0.n21308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__5__5377_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33916\,
            in1 => \N__33466\,
            in2 => \_gnd_net_\,
            in3 => \N__46888\,
            lcout => data_out_frame_7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71043\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40846\,
            in1 => \N__33946\,
            in2 => \_gnd_net_\,
            in3 => \N__43441\,
            lcout => \c0.n5_adj_3475\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i7_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__37531\,
            in1 => \N__33930\,
            in2 => \N__33805\,
            in3 => \N__33881\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71043\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40845\,
            in1 => \N__33915\,
            in2 => \_gnd_net_\,
            in3 => \N__33907\,
            lcout => \c0.n5_adj_3447\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i1_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33880\,
            in1 => \N__33801\,
            in2 => \N__34119\,
            in3 => \N__35926\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71043\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17958_4_lut_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011000100"
        )
    port map (
            in0 => \N__36958\,
            in1 => \N__40844\,
            in2 => \N__33742\,
            in3 => \N__36695\,
            lcout => \c0.n21546\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_15_i6_2_lut_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34869\,
            in2 => \_gnd_net_\,
            in3 => \N__60653\,
            lcout => \c0.n6_adj_3192\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__1__5333_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33703\,
            in1 => \N__33669\,
            in2 => \_gnd_net_\,
            in3 => \N__46642\,
            lcout => data_out_frame_13_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71026\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_16_i6_2_lut_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60654\,
            in2 => \_gnd_net_\,
            in3 => \N__34356\,
            lcout => \c0.n6_adj_3190\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i11148_4_lut_3_lut_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__37920\,
            in1 => \N__56193\,
            in2 => \_gnd_net_\,
            in3 => \N__39231\,
            lcout => OPEN,
            ltout => \c0.rx.n14601_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i0_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000001010100"
        )
    port map (
            in0 => \N__37800\,
            in1 => \N__37858\,
            in2 => \N__34276\,
            in3 => \N__37537\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71026\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_4_lut_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100000101"
        )
    port map (
            in0 => \N__37857\,
            in1 => \N__37799\,
            in2 => \N__37929\,
            in3 => \N__37749\,
            lcout => n12301,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12241_2_lut_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40826\,
            in2 => \_gnd_net_\,
            in3 => \N__36707\,
            lcout => \c0.n15685\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__37851\,
            in1 => \N__37805\,
            in2 => \N__34252\,
            in3 => \N__37912\,
            lcout => \c0.rx.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i7_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39194\,
            in2 => \_gnd_net_\,
            in3 => \N__34633\,
            lcout => \c0.rx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_4_lut_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__37852\,
            in1 => \N__37806\,
            in2 => \N__37753\,
            in3 => \N__37913\,
            lcout => n12492,
            ltout => \n12492_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i9378_3_lut_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39433\,
            in2 => \N__34237\,
            in3 => \N__37853\,
            lcout => n12835,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_o_bdd_4_lut_4_lut_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__34234\,
            in1 => \N__34175\,
            in2 => \N__34120\,
            in3 => \N__34099\,
            lcout => \c0.n21611\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__7__5375_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33979\,
            in1 => \N__33945\,
            in2 => \_gnd_net_\,
            in3 => \N__46887\,
            lcout => data_out_frame_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i0_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__39192\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34309\,
            lcout => \c0.rx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i2_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39193\,
            in2 => \_gnd_net_\,
            in3 => \N__34297\,
            lcout => \c0.rx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_2_lut_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__37652\,
            in1 => \N__37654\,
            in2 => \N__34683\,
            in3 => \N__34303\,
            lcout => n13179,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \c0.rx.n17267\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_3_lut_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__37621\,
            in1 => \N__37617\,
            in2 => \N__34687\,
            in3 => \N__34300\,
            lcout => \c0.rx.n9\,
            ltout => OPEN,
            carryin => \c0.rx.n17267\,
            carryout => \c0.rx.n17268\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_4_lut_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__37687\,
            in1 => \N__37683\,
            in2 => \N__34684\,
            in3 => \N__34291\,
            lcout => n12908,
            ltout => OPEN,
            carryin => \c0.rx.n17268\,
            carryout => \c0.rx.n17269\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_5_lut_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__39151\,
            in1 => \N__39150\,
            in2 => \N__34688\,
            in3 => \N__34288\,
            lcout => n12911,
            ltout => OPEN,
            carryin => \c0.rx.n17269\,
            carryout => \c0.rx.n17270\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_6_lut_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38107\,
            in1 => \N__38106\,
            in2 => \N__34685\,
            in3 => \N__34285\,
            lcout => n12914,
            ltout => OPEN,
            carryin => \c0.rx.n17270\,
            carryout => \c0.rx.n17271\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_7_lut_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38083\,
            in1 => \N__38082\,
            in2 => \N__34689\,
            in3 => \N__34282\,
            lcout => n12917,
            ltout => OPEN,
            carryin => \c0.rx.n17271\,
            carryout => \c0.rx.n17272\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_8_lut_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__37723\,
            in1 => \N__37722\,
            in2 => \N__34686\,
            in3 => \N__34279\,
            lcout => n12920,
            ltout => OPEN,
            carryin => \c0.rx.n17272\,
            carryout => \c0.rx.n17273\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_9_lut_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__39289\,
            in1 => \N__39290\,
            in2 => \N__34690\,
            in3 => \N__34636\,
            lcout => \c0.rx.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_431_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49672\,
            in1 => \N__34557\,
            in2 => \N__34627\,
            in3 => \N__34590\,
            lcout => \c0.n45_adj_3262\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_12_i6_2_lut_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__60618\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34507\,
            lcout => \c0.n6_adj_3161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_25_i6_2_lut_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34558\,
            in2 => \_gnd_net_\,
            in3 => \N__60620\,
            lcout => \c0.n6_adj_3172\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_14_i6_2_lut_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__60619\,
            in1 => \N__34464\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n6_adj_3194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_427_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34506\,
            in1 => \N__34481\,
            in2 => \N__34465\,
            in3 => \N__34440\,
            lcout => \c0.n43_adj_3257\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_11_i6_2_lut_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60617\,
            in2 => \_gnd_net_\,
            in3 => \N__34336\,
            lcout => \c0.n6_adj_3160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_502_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__40111\,
            in1 => \N__40286\,
            in2 => \N__49678\,
            in3 => \N__40201\,
            lcout => \c0.n12_adj_3361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_428_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34386\,
            in1 => \N__35380\,
            in2 => \N__34363\,
            in3 => \N__34335\,
            lcout => OPEN,
            ltout => \c0.n41_adj_3258_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_4_lut_adj_430_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35023\,
            in1 => \N__37966\,
            in2 => \N__34909\,
            in3 => \N__34906\,
            lcout => \c0.n50_adj_3261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_429_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34900\,
            in1 => \N__34873\,
            in2 => \N__35302\,
            in3 => \N__34849\,
            lcout => \c0.n40_adj_3259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_2_lut_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35332\,
            in2 => \_gnd_net_\,
            in3 => \N__34816\,
            lcout => OPEN,
            ltout => \c0.n39_adj_3260_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_4_lut_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34783\,
            in1 => \N__34777\,
            in2 => \N__34771\,
            in3 => \N__34768\,
            lcout => \c0.n11440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_930_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__42364\,
            in1 => \N__35173\,
            in2 => \N__34969\,
            in3 => \N__34699\,
            lcout => OPEN,
            ltout => \c0.n14_adj_3080_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i1_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__38354\,
            in1 => \N__34762\,
            in2 => \N__34744\,
            in3 => \N__34741\,
            lcout => \FRAME_MATCHER_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71093\,
            ce => 'H',
            sr => \N__46803\
        );

    \c0.i1_3_lut_4_lut_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__34728\,
            in1 => \N__34950\,
            in2 => \N__42496\,
            in3 => \N__42310\,
            lcout => \c0.n19119\,
            ltout => \c0.n19119_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_463_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__34965\,
            in1 => \_gnd_net_\,
            in2 => \N__34693\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.n5_adj_3306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i0_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__39567\,
            in1 => \N__34981\,
            in2 => \N__34972\,
            in3 => \N__38317\,
            lcout => \c0.FRAME_MATCHER_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71093\,
            ce => 'H',
            sr => \N__46803\
        );

    \c0.i1_2_lut_adj_460_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__35123\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35154\,
            lcout => \c0.n2_adj_3302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__5__5168_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__67983\,
            in1 => \N__53176\,
            in2 => \_gnd_net_\,
            in3 => \N__39743\,
            lcout => data_in_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_423_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38519\,
            in2 => \_gnd_net_\,
            in3 => \N__38413\,
            lcout => \c0.n9389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_581_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__39557\,
            in1 => \N__42427\,
            in2 => \N__38989\,
            in3 => \N__38258\,
            lcout => \c0.n11433\,
            ltout => \c0.n11433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_adj_757_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__42428\,
            in1 => \N__38211\,
            in2 => \N__34957\,
            in3 => \N__42293\,
            lcout => OPEN,
            ltout => \c0.n8_adj_3228_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_396_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000010000"
        )
    port map (
            in0 => \N__38976\,
            in1 => \N__42429\,
            in2 => \N__34954\,
            in3 => \N__35423\,
            lcout => \c0.n2103\,
            ltout => \c0.n2103_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_940_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38520\,
            in2 => \N__34936\,
            in3 => \N__38414\,
            lcout => \c0.n1_adj_3002\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__3__5194_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53195\,
            in1 => \N__39954\,
            in2 => \_gnd_net_\,
            in3 => \N__40012\,
            lcout => data_in_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_509_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41365\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34933\,
            lcout => \c0.n18653\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_657_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__38266\,
            in1 => \N__42459\,
            in2 => \_gnd_net_\,
            in3 => \N__39569\,
            lcout => n4_adj_3596,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__39891\,
            in1 => \N__38457\,
            in2 => \_gnd_net_\,
            in3 => \N__38469\,
            lcout => \c0.FRAME_MATCHER_state_31_N_1736_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_928_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__38458\,
            in1 => \N__42460\,
            in2 => \N__39895\,
            in3 => \N__38416\,
            lcout => \c0.FRAME_MATCHER_state_31_N_1736_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_23_i6_2_lut_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60633\,
            in2 => \_gnd_net_\,
            in3 => \N__38019\,
            lcout => \c0.n6_adj_3176\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_939_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__35150\,
            in1 => \N__38515\,
            in2 => \N__35133\,
            in3 => \N__38415\,
            lcout => \c0.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_424_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35012\,
            in1 => \N__35083\,
            in2 => \N__35059\,
            in3 => \N__35251\,
            lcout => \c0.n44_adj_3255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__5__5176_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53215\,
            in1 => \N__39744\,
            in2 => \_gnd_net_\,
            in3 => \N__41877\,
            lcout => data_in_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71153\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_24_i6_2_lut_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60583\,
            in2 => \_gnd_net_\,
            in3 => \N__35014\,
            lcout => \c0.n6_adj_3174\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_854_LC_15_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35473\,
            in2 => \_gnd_net_\,
            in3 => \N__41429\,
            lcout => \c0.n18675\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_4_lut_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__42328\,
            in1 => \N__42368\,
            in2 => \N__42497\,
            in3 => \N__35436\,
            lcout => n2108,
            ltout => \n2108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_26_i6_2_lut_LC_15_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35376\,
            in2 => \N__35356\,
            in3 => \_gnd_net_\,
            lcout => \c0.n6_adj_3170\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_29_i6_2_lut_LC_15_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60585\,
            in2 => \_gnd_net_\,
            in3 => \N__37992\,
            lcout => \c0.n6_adj_3165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_27_i6_2_lut_LC_15_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35328\,
            in2 => \_gnd_net_\,
            in3 => \N__60584\,
            lcout => \c0.n6_adj_3168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_28_i6_2_lut_LC_15_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35292\,
            in2 => \_gnd_net_\,
            in3 => \N__60632\,
            lcout => \c0.n6_adj_3166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_31_i6_2_lut_LC_15_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__60635\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38134\,
            lcout => \c0.n6_adj_3159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_30_i6_2_lut_LC_15_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35247\,
            in2 => \_gnd_net_\,
            in3 => \N__60634\,
            lcout => \c0.n6_adj_3164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_61_i9_2_lut_3_lut_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__60204\,
            in1 => \N__59977\,
            in2 => \_gnd_net_\,
            in3 => \N__60108\,
            lcout => \c0.n9_adj_3038\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_6_i6_2_lut_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60717\,
            in2 => \_gnd_net_\,
            in3 => \N__40186\,
            lcout => \c0.n6_adj_3150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_82_i11_2_lut_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49665\,
            in2 => \_gnd_net_\,
            in3 => \N__40185\,
            lcout => \c0.n11_adj_3093\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i12_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36255\,
            in1 => \N__37046\,
            in2 => \_gnd_net_\,
            in3 => \N__35791\,
            lcout => encoder1_position_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71156\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17732_4_lut_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__37466\,
            in1 => \N__38542\,
            in2 => \N__35999\,
            in3 => \N__35737\,
            lcout => \c0.n21319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__2__5380_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35767\,
            in1 => \N__35914\,
            in2 => \_gnd_net_\,
            in3 => \N__46859\,
            lcout => data_out_frame_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71140\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17730_4_lut_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__35902\,
            in1 => \N__36759\,
            in2 => \N__36988\,
            in3 => \N__35848\,
            lcout => \c0.n21317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i27_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35722\,
            in1 => \N__35529\,
            in2 => \_gnd_net_\,
            in3 => \N__35563\,
            lcout => encoder0_position_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71140\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35514\,
            in1 => \N__35503\,
            in2 => \_gnd_net_\,
            in3 => \N__40938\,
            lcout => \c0.n5_adj_3380\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17735_4_lut_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__37467\,
            in1 => \N__40654\,
            in2 => \N__36007\,
            in3 => \N__35479\,
            lcout => OPEN,
            ltout => \c0.n21322_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_3_lut_4_lut_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__37345\,
            in1 => \N__35941\,
            in2 => \N__35929\,
            in3 => \N__37468\,
            lcout => n10_adj_3594,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35913\,
            in1 => \N__35871\,
            in2 => \_gnd_net_\,
            in3 => \N__40937\,
            lcout => \c0.n5_adj_3106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_62_i9_2_lut_3_lut_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__60256\,
            in1 => \N__59978\,
            in2 => \_gnd_net_\,
            in3 => \N__60116\,
            lcout => \c0.n9_adj_3101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_0__2__5436_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__39490\,
            in1 => \N__35860\,
            in2 => \N__37092\,
            in3 => \N__39003\,
            lcout => \c0.data_out_frame_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__2__5388_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46856\,
            in1 => \N__35896\,
            in2 => \_gnd_net_\,
            in3 => \N__35872\,
            lcout => data_out_frame_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17928_2_lut_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36716\,
            in2 => \_gnd_net_\,
            in3 => \N__35859\,
            lcout => OPEN,
            ltout => \c0.n21473_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100000010000"
        )
    port map (
            in0 => \N__36969\,
            in1 => \N__40906\,
            in2 => \N__35851\,
            in3 => \N__36403\,
            lcout => \c0.n6_adj_3105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__6__5208_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__46855\,
            in1 => \N__50605\,
            in2 => \N__54481\,
            in3 => \N__35829\,
            lcout => data_out_frame_28_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_0__3__5435_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__39491\,
            in1 => \N__35815\,
            in2 => \N__37093\,
            in3 => \N__39004\,
            lcout => \c0.data_out_frame_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_3_lut_4_lut_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55511\,
            in1 => \N__51345\,
            in2 => \N__57379\,
            in3 => \N__51291\,
            lcout => \c0.n39_adj_3339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i101_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66194\,
            in1 => \N__67197\,
            in2 => \N__44624\,
            in3 => \N__72697\,
            lcout => \c0.data_in_frame_12_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__37183\,
            in1 => \N__36330\,
            in2 => \N__40936\,
            in3 => \_gnd_net_\,
            lcout => \c0.n11_adj_3325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__0__5342_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46848\,
            in2 => \N__36334\,
            in3 => \N__36370\,
            lcout => data_out_frame_12_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__7__5343_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__36318\,
            in1 => \N__36291\,
            in2 => \N__46916\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame_11_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i28_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36277\,
            in1 => \N__36262\,
            in2 => \_gnd_net_\,
            in3 => \N__36074\,
            lcout => encoder1_position_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__6__5392_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__36049\,
            in1 => \N__38632\,
            in2 => \N__46917\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36037\,
            in1 => \N__36018\,
            in2 => \_gnd_net_\,
            in3 => \N__40923\,
            lcout => OPEN,
            ltout => \c0.n26_adj_3382_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17729_4_lut_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__37464\,
            in1 => \N__36000\,
            in2 => \N__35965\,
            in3 => \N__35962\,
            lcout => \c0.n21316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__4__5394_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__46865\,
            in1 => \_gnd_net_\,
            in2 => \N__36487\,
            in3 => \N__38752\,
            lcout => data_out_frame_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17913_2_lut_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36483\,
            in2 => \_gnd_net_\,
            in3 => \N__40892\,
            lcout => \c0.n21465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__0__5398_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36460\,
            in1 => \N__39088\,
            in2 => \_gnd_net_\,
            in3 => \N__46866\,
            lcout => \c0.data_out_frame_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i5_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36441\,
            in1 => \N__55384\,
            in2 => \_gnd_net_\,
            in3 => \N__41096\,
            lcout => control_mode_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17980_4_lut_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__36430\,
            in1 => \N__36949\,
            in2 => \N__36418\,
            in3 => \N__36735\,
            lcout => \c0.n21568\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__2__5396_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46864\,
            in1 => \N__38620\,
            in2 => \_gnd_net_\,
            in3 => \N__36402\,
            lcout => data_out_frame_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i205_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66899\,
            in1 => \N__63395\,
            in2 => \N__59669\,
            in3 => \N__72711\,
            lcout => \c0.data_in_frame_25_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i146_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__71485\,
            in1 => \N__63937\,
            in2 => \_gnd_net_\,
            in3 => \N__45234\,
            lcout => data_in_frame_18_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i1_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39204\,
            in2 => \_gnd_net_\,
            in3 => \N__36388\,
            lcout => \c0.rx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i6_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__39205\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37165\,
            lcout => \c0.rx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__7__5391_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38722\,
            in1 => \N__37006\,
            in2 => \_gnd_net_\,
            in3 => \N__46764\,
            lcout => data_out_frame_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50863\,
            in1 => \N__54976\,
            in2 => \N__50944\,
            in3 => \N__50829\,
            lcout => \c0.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_243_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__37153\,
            in1 => \N__37135\,
            in2 => \N__37111\,
            in3 => \N__38812\,
            lcout => \c0.n12254\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__4__5338_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__37059\,
            in1 => \N__37023\,
            in2 => \N__46857\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame_12_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71056\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17988_3_lut_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__36960\,
            in1 => \N__37005\,
            in2 => \_gnd_net_\,
            in3 => \N__40886\,
            lcout => OPEN,
            ltout => \c0.n21576_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17715_4_lut_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__36994\,
            in1 => \N__36961\,
            in2 => \N__36769\,
            in3 => \N__36697\,
            lcout => OPEN,
            ltout => \c0.n21302_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17717_4_lut_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__46951\,
            in1 => \N__37524\,
            in2 => \N__36508\,
            in3 => \N__37462\,
            lcout => OPEN,
            ltout => \c0.n21304_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_3_lut_4_lut_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__37463\,
            in1 => \N__37344\,
            in2 => \N__36505\,
            in3 => \N__36502\,
            lcout => n9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17723_4_lut_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__37525\,
            in1 => \N__37460\,
            in2 => \N__37498\,
            in3 => \N__37474\,
            lcout => OPEN,
            ltout => \c0.n21310_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_3_lut_4_lut_adj_620_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__37461\,
            in1 => \N__37343\,
            in2 => \N__37255\,
            in3 => \N__37252\,
            lcout => n9_adj_3590,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i3_4_lut_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__37849\,
            in1 => \N__37796\,
            in2 => \N__37930\,
            in3 => \N__37744\,
            lcout => \c0.rx.n11302\,
            ltout => \c0.rx.n11302_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37219\,
            in3 => \N__39335\,
            lcout => n11466,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__0__5334_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37216\,
            in1 => \N__37182\,
            in2 => \_gnd_net_\,
            in3 => \N__46643\,
            lcout => data_out_frame_13_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71035\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i17914_2_lut_3_lut_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__56213\,
            in1 => \N__37927\,
            in2 => \_gnd_net_\,
            in3 => \N__39221\,
            lcout => OPEN,
            ltout => \c0.rx.n21451_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i1_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001110010"
        )
    port map (
            in0 => \N__37850\,
            in1 => \N__37570\,
            in2 => \N__37168\,
            in3 => \N__37797\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71035\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_516_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__40280\,
            in1 => \N__49677\,
            in2 => \N__40126\,
            in3 => \N__40200\,
            lcout => \c0.n12_adj_3006\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i147_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43116\,
            in1 => \N__63915\,
            in2 => \_gnd_net_\,
            in3 => \N__68622\,
            lcout => data_in_frame_18_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71035\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_adj_656_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63576\,
            in2 => \_gnd_net_\,
            in3 => \N__63651\,
            lcout => \c0.n27_adj_3455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_4_lut_adj_213_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__39136\,
            in1 => \N__37715\,
            in2 => \N__37564\,
            in3 => \N__39244\,
            lcout => \c0.rx.n15906\,
            ltout => \c0.rx.n15906_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_adj_208_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__39284\,
            in1 => \_gnd_net_\,
            in2 => \N__37573\,
            in3 => \N__37922\,
            lcout => \c0.rx.n20851\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_211_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37682\,
            in2 => \_gnd_net_\,
            in3 => \N__37610\,
            lcout => \c0.rx.n32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i2_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39285\,
            in2 => \_gnd_net_\,
            in3 => \N__37549\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71057\,
            ce => 'H',
            sr => \N__37555\
        );

    \c0.rx.i2_3_lut_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__37862\,
            in1 => \N__37921\,
            in2 => \_gnd_net_\,
            in3 => \N__37801\,
            lcout => \c0.rx.n20964\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i12463_2_lut_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39283\,
            in2 => \_gnd_net_\,
            in3 => \N__37548\,
            lcout => \r_SM_Main_2_N_2473_2\,
            ltout => \r_SM_Main_2_N_2473_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39432\,
            in2 => \N__37540\,
            in3 => \N__37923\,
            lcout => \c0.rx.n15926\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_215_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38104\,
            in2 => \_gnd_net_\,
            in3 => \N__38080\,
            lcout => \c0.rx.n11455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_214_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37680\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37648\,
            lcout => OPEN,
            ltout => \c0.rx.n35_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i5_4_lut_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100010"
        )
    port map (
            in0 => \N__37714\,
            in1 => \N__38059\,
            in2 => \N__37933\,
            in3 => \N__56154\,
            lcout => OPEN,
            ltout => \c0.rx.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i17900_4_lut_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110110011"
        )
    port map (
            in0 => \N__37585\,
            in1 => \N__37928\,
            in2 => \N__37873\,
            in3 => \N__39142\,
            lcout => OPEN,
            ltout => \c0.rx.n21406_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_adj_216_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__37863\,
            in1 => \N__37798\,
            in2 => \N__37756\,
            in3 => \N__37748\,
            lcout => n3792,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_3_lut_4_lut_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__37679\,
            in1 => \N__37713\,
            in2 => \N__37653\,
            in3 => \N__37608\,
            lcout => \c0.rx.n6_adj_2995\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__37681\,
            in1 => \N__37647\,
            in2 => \_gnd_net_\,
            in3 => \N__37609\,
            lcout => \c0.rx.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i4_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39190\,
            in2 => \_gnd_net_\,
            in3 => \N__37579\,
            lcout => \c0.rx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71082\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_925_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__44260\,
            in1 => \N__71623\,
            in2 => \_gnd_net_\,
            in3 => \N__59432\,
            lcout => n19129,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i5_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39191\,
            in2 => \_gnd_net_\,
            in3 => \N__38200\,
            lcout => \c0.rx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71082\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_432_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__40110\,
            in1 => \N__40285\,
            in2 => \_gnd_net_\,
            in3 => \N__38186\,
            lcout => OPEN,
            ltout => \c0.n11317_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12193_3_lut_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111010"
        )
    port map (
            in0 => \N__64340\,
            in1 => \_gnd_net_\,
            in2 => \N__38170\,
            in3 => \N__38160\,
            lcout => \c0.n3632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i119_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__69001\,
            in1 => \N__64136\,
            in2 => \N__64887\,
            in3 => \N__62018\,
            lcout => \c0.data_in_frame_14_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71082\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i17680_2_lut_3_lut_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__39292\,
            in1 => \N__38105\,
            in2 => \_gnd_net_\,
            in3 => \N__38081\,
            lcout => \c0.rx.n21267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_426_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38050\,
            in1 => \N__40199\,
            in2 => \N__38026\,
            in3 => \N__37999\,
            lcout => \c0.n42_adj_3256\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_920_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__61955\,
            in1 => \N__71624\,
            in2 => \_gnd_net_\,
            in3 => \N__59448\,
            lcout => n19127,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_228_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101110"
        )
    port map (
            in0 => \N__37959\,
            in1 => \N__38277\,
            in2 => \N__42495\,
            in3 => \N__37942\,
            lcout => \c0.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12257_2_lut_4_lut_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__53079\,
            in1 => \N__38373\,
            in2 => \N__38806\,
            in3 => \N__42369\,
            lcout => \c0.n15701\,
            ltout => \c0.n15701_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_864_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__40287\,
            in1 => \N__38398\,
            in2 => \N__38386\,
            in3 => \N__40125\,
            lcout => \c0.n19098\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_658_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__38931\,
            in1 => \N__39552\,
            in2 => \_gnd_net_\,
            in3 => \N__38248\,
            lcout => n11421,
            ltout => \n11421_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_483_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38383\,
            in3 => \N__42426\,
            lcout => \c0.n11422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__6__5167_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__69012\,
            in1 => \N__53174\,
            in2 => \_gnd_net_\,
            in3 => \N__52949\,
            lcout => data_in_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71111\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_662_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__38348\,
            in1 => \N__38212\,
            in2 => \N__38964\,
            in3 => \N__38313\,
            lcout => \c0.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i117_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__72775\,
            in1 => \N__64113\,
            in2 => \N__61987\,
            in3 => \N__45127\,
            lcout => \c0.data_in_frame_14_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71111\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_885_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66121\,
            in2 => \_gnd_net_\,
            in3 => \N__59439\,
            lcout => \c0.n19140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__6__5183_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__52919\,
            in1 => \N__53177\,
            in2 => \_gnd_net_\,
            in3 => \N__39802\,
            lcout => data_in_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_482_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__39556\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38265\,
            lcout => \c0.n15874\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_421_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__43907\,
            in1 => \N__49754\,
            in2 => \N__47014\,
            in3 => \N__39846\,
            lcout => \c0.n21_adj_3253\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__1__5180_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39847\,
            in1 => \N__53178\,
            in2 => \_gnd_net_\,
            in3 => \N__43908\,
            lcout => data_in_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i201_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__63412\,
            in1 => \N__66849\,
            in2 => \N__53379\,
            in3 => \N__65172\,
            lcout => \c0.data_in_frame_25_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12187_3_lut_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__38425\,
            in1 => \N__38978\,
            in2 => \_gnd_net_\,
            in3 => \N__38449\,
            lcout => \c0.n121\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__3__5170_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__69376\,
            in1 => \N__53175\,
            in2 => \_gnd_net_\,
            in3 => \N__39867\,
            lcout => data_in_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_417_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__47034\,
            in1 => \N__39980\,
            in2 => \N__47013\,
            in3 => \N__39751\,
            lcout => \c0.n63_adj_3083\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_312_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__49755\,
            in1 => \N__38533\,
            in2 => \_gnd_net_\,
            in3 => \N__40579\,
            lcout => \c0.n103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__38436\,
            in1 => \N__38443\,
            in2 => \_gnd_net_\,
            in3 => \N__39711\,
            lcout => \c0.n63_adj_3084\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_420_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__39866\,
            in1 => \N__39666\,
            in2 => \N__39829\,
            in3 => \N__41902\,
            lcout => \c0.n19_adj_3252\,
            ltout => \c0.n19_adj_3252_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4379_2_lut_4_lut_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__38437\,
            in1 => \N__39712\,
            in2 => \N__38428\,
            in3 => \N__38424\,
            lcout => \c0.n7804\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__6__5191_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53172\,
            in1 => \N__39981\,
            in2 => \_gnd_net_\,
            in3 => \N__39806\,
            lcout => data_in_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71155\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__2__5195_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38494\,
            in1 => \N__53173\,
            in2 => \_gnd_net_\,
            in3 => \N__39667\,
            lcout => data_in_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71155\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17694_4_lut_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__41876\,
            in1 => \N__40004\,
            in2 => \N__42636\,
            in3 => \N__38493\,
            lcout => OPEN,
            ltout => \c0.n21281_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_399_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__39775\,
            in1 => \N__42589\,
            in2 => \N__38536\,
            in3 => \N__42544\,
            lcout => \c0.n108\,
            ltout => \c0.n108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_422_LC_16_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__40575\,
            in1 => \N__39879\,
            in2 => \N__38527\,
            in3 => \N__49734\,
            lcout => \c0.n92_adj_3254\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i231_LC_16_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__66933\,
            in1 => \N__69024\,
            in2 => \N__39702\,
            in3 => \N__67199\,
            lcout => \c0.data_in_frame_28_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71155\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__0__5181_LC_16_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53216\,
            in1 => \N__49756\,
            in2 => \_gnd_net_\,
            in3 => \N__42632\,
            lcout => data_in_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71166\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_411_LC_16_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__40003\,
            in1 => \N__41875\,
            in2 => \N__39808\,
            in3 => \N__38491\,
            lcout => \c0.n18_adj_3246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__2__5187_LC_16_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__38492\,
            in1 => \N__53217\,
            in2 => \_gnd_net_\,
            in3 => \N__41929\,
            lcout => data_in_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71166\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_259_LC_16_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40316\,
            in2 => \_gnd_net_\,
            in3 => \N__41428\,
            lcout => \c0.n18655\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i0_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__43762\,
            in1 => \N__65148\,
            in2 => \N__56236\,
            in3 => \N__56084\,
            lcout => rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71190\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40590\,
            in2 => \N__40615\,
            in3 => \N__40942\,
            lcout => \c0.n26_adj_3107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_725_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__54706\,
            in1 => \N__38551\,
            in2 => \N__55402\,
            in3 => \N__40597\,
            lcout => \c0.n15499\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i53_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__72614\,
            in1 => \N__61677\,
            in2 => \N__46369\,
            in3 => \N__61927\,
            lcout => \c0.data_in_frame_6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71179\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_2_lut_adj_358_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54254\,
            in2 => \_gnd_net_\,
            in3 => \N__61117\,
            lcout => \c0.n37_adj_3153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_477_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__54589\,
            in1 => \N__54892\,
            in2 => \N__40639\,
            in3 => \N__55184\,
            lcout => \c0.n38_adj_3328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i155_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__69168\,
            in1 => \_gnd_net_\,
            in2 => \N__65762\,
            in3 => \N__68655\,
            lcout => data_in_frame_19_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i118_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__61954\,
            in1 => \N__64248\,
            in2 => \N__44712\,
            in3 => \N__67922\,
            lcout => \c0.data_in_frame_14_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17692_4_lut_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__46302\,
            in1 => \N__47221\,
            in2 => \N__42703\,
            in3 => \N__54468\,
            lcout => OPEN,
            ltout => \c0.n21279_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_adj_480_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__47311\,
            in1 => \N__38575\,
            in2 => \N__38569\,
            in3 => \N__38563\,
            lcout => \FRAME_MATCHER_state_31_N_1800_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17668_2_lut_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47560\,
            in2 => \_gnd_net_\,
            in3 => \N__56852\,
            lcout => OPEN,
            ltout => \c0.n21255_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_488_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__62172\,
            in1 => \N__50360\,
            in2 => \N__38566\,
            in3 => \N__55054\,
            lcout => \c0.n37_adj_3332\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_2_lut_3_lut_adj_555_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__61246\,
            in1 => \_gnd_net_\,
            in2 => \N__38607\,
            in3 => \N__44310\,
            lcout => \c0.n63_adj_3417\,
            ltout => \c0.n63_adj_3417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_2_lut_3_lut_4_lut_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41027\,
            in1 => \N__44049\,
            in2 => \N__38557\,
            in3 => \N__51259\,
            lcout => \c0.n40_adj_3032\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_2_lut_3_lut_4_lut_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51260\,
            in1 => \N__41028\,
            in2 => \N__44053\,
            in3 => \N__50500\,
            lcout => \c0.n34_adj_3411\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_554_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44311\,
            in1 => \N__38600\,
            in2 => \_gnd_net_\,
            in3 => \N__41029\,
            lcout => \c0.n5_adj_3040\,
            ltout => \c0.n5_adj_3040_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_533_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__51258\,
            in1 => \_gnd_net_\,
            in2 => \N__38554\,
            in3 => \N__44048\,
            lcout => \c0.n11537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_433_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__41014\,
            in1 => \N__57289\,
            in2 => \N__42756\,
            in3 => \N__50830\,
            lcout => \c0.n30_adj_3264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i41_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__65069\,
            in1 => \N__61795\,
            in2 => \N__38608\,
            in3 => \N__60309\,
            lcout => \c0.data_in_frame_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71157\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i43_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__61794\,
            in1 => \N__68656\,
            in2 => \N__60329\,
            in3 => \N__61247\,
            lcout => \c0.data_in_frame_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71157\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56846\,
            in1 => \N__61122\,
            in2 => \N__54472\,
            in3 => \N__46303\,
            lcout => \c0.n6_adj_3343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_242_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55549\,
            in1 => \N__49813\,
            in2 => \N__38589\,
            in3 => \N__61351\,
            lcout => \c0.n19493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i103_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66038\,
            in1 => \N__67196\,
            in2 => \N__66286\,
            in3 => \N__68928\,
            lcout => \c0.data_in_frame_12_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i80_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__72284\,
            in1 => \N__63281\,
            in2 => \N__38590\,
            in3 => \N__66039\,
            lcout => \c0.data_in_frame_9_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i42_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__60319\,
            in1 => \N__61797\,
            in2 => \N__51406\,
            in3 => \N__71436\,
            lcout => \c0.data_in_frame_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i19_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__61796\,
            in1 => \N__44247\,
            in2 => \N__68724\,
            in3 => \N__46333\,
            lcout => \c0.data_in_frame_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i125_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__64410\,
            in1 => \N__64220\,
            in2 => \N__51582\,
            in3 => \N__72672\,
            lcout => \c0.data_in_frame_15_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_868_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__59992\,
            in1 => \N__60121\,
            in2 => \N__60264\,
            in3 => \N__59481\,
            lcout => \c0.n19115\,
            ltout => \c0.n19115_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i77_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__41141\,
            in1 => \N__66046\,
            in2 => \N__38692\,
            in3 => \N__72673\,
            lcout => \c0.data_in_frame_9_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43149\,
            in1 => \N__38763\,
            in2 => \N__38689\,
            in3 => \N__50659\,
            lcout => \c0.n16_adj_3018\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_653_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49921\,
            in1 => \N__54893\,
            in2 => \N__42940\,
            in3 => \N__42969\,
            lcout => \c0.n12_adj_3477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i82_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__66045\,
            in1 => \N__38688\,
            in2 => \N__71525\,
            in3 => \N__62846\,
            lcout => \c0.data_in_frame_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i74_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__71492\,
            in1 => \N__63280\,
            in2 => \N__66120\,
            in3 => \N__56707\,
            lcout => \c0.data_in_frame_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_696_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__44893\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52206\,
            lcout => \c0.n16_adj_3489\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_575_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__42757\,
            in1 => \N__41566\,
            in2 => \N__39628\,
            in3 => \N__41755\,
            lcout => OPEN,
            ltout => \c0.n20_adj_3437_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_582_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41647\,
            in1 => \N__38669\,
            in2 => \N__38638\,
            in3 => \N__39304\,
            lcout => n21222,
            ltout => \n21222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i6_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38631\,
            in2 => \N__38635\,
            in3 => \N__54895\,
            lcout => control_mode_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i2_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38619\,
            in1 => \N__60412\,
            in2 => \_gnd_net_\,
            in3 => \N__41086\,
            lcout => control_mode_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i4_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__38751\,
            in1 => \_gnd_net_\,
            in2 => \N__41097\,
            in3 => \N__60931\,
            lcout => control_mode_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i3_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38733\,
            in1 => \N__61231\,
            in2 => \_gnd_net_\,
            in3 => \N__41087\,
            lcout => control_mode_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i7_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38715\,
            in2 => \N__41098\,
            in3 => \N__54691\,
            lcout => control_mode_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i145_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__51171\,
            in1 => \N__63944\,
            in2 => \_gnd_net_\,
            in3 => \N__65070\,
            lcout => data_in_frame_18_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71095\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45141\,
            in2 => \_gnd_net_\,
            in3 => \N__63862\,
            lcout => \c0.n6_adj_3005\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_225_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41551\,
            in2 => \_gnd_net_\,
            in3 => \N__44545\,
            lcout => \c0.n9\,
            ltout => \c0.n9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_4_lut_adj_908_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__52827\,
            in1 => \N__45459\,
            in2 => \N__38704\,
            in3 => \N__45715\,
            lcout => OPEN,
            ltout => \c0.n16_adj_3008_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_233_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56313\,
            in1 => \N__41190\,
            in2 => \N__38701\,
            in3 => \N__43023\,
            lcout => \c0.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_693_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43024\,
            in1 => \N__56314\,
            in2 => \N__41194\,
            in3 => \N__38698\,
            lcout => \c0.n19449\,
            ltout => \c0.n19449_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_694_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45460\,
            in1 => \N__50904\,
            in2 => \N__39091\,
            in3 => \N__45640\,
            lcout => \c0.n12218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i0_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39087\,
            in1 => \N__55053\,
            in2 => \_gnd_net_\,
            in3 => \N__41094\,
            lcout => control_mode_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71095\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_3_lut_adj_489_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__39060\,
            in1 => \N__38997\,
            in2 => \_gnd_net_\,
            in3 => \N__38837\,
            lcout => \c0.n13_adj_3016\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i139_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__68521\,
            in1 => \N__63357\,
            in2 => \N__71792\,
            in3 => \N__68348\,
            lcout => \c0.data_in_frame_17_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__38802\,
            in1 => \N__44127\,
            in2 => \N__53118\,
            in3 => \N__42132\,
            lcout => \c0.n19111\,
            ltout => \c0.n19111_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i104_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__66125\,
            in1 => \N__57071\,
            in2 => \N__38770\,
            in3 => \N__72295\,
            lcout => \c0.data_in_frame_12_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_226_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38767\,
            in2 => \_gnd_net_\,
            in3 => \N__55618\,
            lcout => \c0.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i2_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__41533\,
            in1 => \N__68522\,
            in2 => \N__56080\,
            in3 => \N__56200\,
            lcout => rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50077\,
            in1 => \N__47509\,
            in2 => \N__56359\,
            in3 => \N__51109\,
            lcout => OPEN,
            ltout => \c0.n28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39112\,
            in1 => \N__39106\,
            in2 => \N__39100\,
            in3 => \N__54467\,
            lcout => \c0.n12026\,
            ltout => \c0.n12026_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_230_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39097\,
            in3 => \N__45137\,
            lcout => \c0.n5_adj_3003\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_403_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51623\,
            in1 => \N__48082\,
            in2 => \N__64723\,
            in3 => \N__52020\,
            lcout => \c0.n32_adj_3236\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i150_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__67982\,
            in1 => \N__63948\,
            in2 => \_gnd_net_\,
            in3 => \N__44892\,
            lcout => data_in_frame_18_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71070\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i212_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__69314\,
            in1 => \N__66754\,
            in2 => \N__67562\,
            in3 => \N__62845\,
            lcout => \c0.data_in_frame_26_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71070\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_386_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64834\,
            in2 => \_gnd_net_\,
            in3 => \N__72858\,
            lcout => \c0.n11_adj_3219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44717\,
            in2 => \_gnd_net_\,
            in3 => \N__48402\,
            lcout => \c0.n10\,
            ltout => \c0.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_897_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41218\,
            in1 => \N__65849\,
            in2 => \N__39094\,
            in3 => \N__47773\,
            lcout => \c0.n12_adj_3004\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_232_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57725\,
            in2 => \_gnd_net_\,
            in3 => \N__48650\,
            lcout => \c0.n19551\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_4_lut_adj_685_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52345\,
            in1 => \N__44718\,
            in2 => \N__68364\,
            in3 => \N__47692\,
            lcout => \c0.n20_adj_3487\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_571_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__41518\,
            in1 => \N__41734\,
            in2 => \N__45985\,
            in3 => \N__43348\,
            lcout => \c0.n21104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i112_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66060\,
            in1 => \N__71941\,
            in2 => \N__56017\,
            in3 => \N__72283\,
            lcout => \c0.data_in_frame_13_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71047\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1998_2_lut_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43801\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39343\,
            lcout => OPEN,
            ltout => \n3846_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i2_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__43849\,
            in1 => \N__39402\,
            in2 => \N__39295\,
            in3 => \N__39375\,
            lcout => \r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_817_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__68355\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__68299\,
            lcout => \c0.n5_adj_3220\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i0_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__39344\,
            in1 => \N__39401\,
            in2 => \_gnd_net_\,
            in3 => \N__39374\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i4_4_lut_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39291\,
            in1 => \N__39250\,
            in2 => \N__39143\,
            in3 => \N__39243\,
            lcout => \c0.rx.r_SM_Main_2_N_2479_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_96_i4_2_lut_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43840\,
            in2 => \_gnd_net_\,
            in3 => \N__43800\,
            lcout => n4_adj_3595,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i3_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39195\,
            in2 => \_gnd_net_\,
            in3 => \N__39163\,
            lcout => \c0.rx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_adj_207_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__39342\,
            in1 => \N__43839\,
            in2 => \_gnd_net_\,
            in3 => \N__43799\,
            lcout => \c0.rx.n15860\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i12_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41496\,
            in2 => \_gnd_net_\,
            in3 => \N__40551\,
            lcout => \c0.FRAME_MATCHER_state_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71084\,
            ce => 'H',
            sr => \N__41284\
        );

    \c0.data_in_frame_0__i229_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__72766\,
            in1 => \N__41578\,
            in2 => \N__66850\,
            in3 => \N__67144\,
            lcout => \c0.data_in_frame_28_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71096\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_613_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65693\,
            in1 => \N__59115\,
            in2 => \N__41604\,
            in3 => \N__39418\,
            lcout => \c0.n13_adj_3463\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i49_4_lut_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58495\,
            in1 => \N__58276\,
            in2 => \N__41275\,
            in3 => \N__48460\,
            lcout => \c0.n100_adj_3403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i221_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__66917\,
            in1 => \N__72767\,
            in2 => \N__48830\,
            in3 => \N__64585\,
            lcout => \c0.data_in_frame_27_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71096\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i1_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__39406\,
            in1 => \N__43790\,
            in2 => \N__39382\,
            in3 => \N__39345\,
            lcout => \r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71096\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_2_lut_3_lut_4_lut_adj_587_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65527\,
            in1 => \N__63778\,
            in2 => \N__63583\,
            in3 => \N__43093\,
            lcout => \c0.n34_adj_3096\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_439_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48789\,
            in2 => \_gnd_net_\,
            in3 => \N__41721\,
            lcout => OPEN,
            ltout => \c0.n22_adj_3276_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_441_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41977\,
            in1 => \N__41706\,
            in2 => \N__39307\,
            in3 => \N__45766\,
            lcout => OPEN,
            ltout => \c0.n36_adj_3277_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_442_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49024\,
            in1 => \N__51760\,
            in2 => \N__39643\,
            in3 => \N__45780\,
            lcout => OPEN,
            ltout => \c0.n20415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_537_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__46027\,
            in1 => \N__59302\,
            in2 => \N__39640\,
            in3 => \N__41674\,
            lcout => OPEN,
            ltout => \c0.n14_adj_3407_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_544_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110111"
        )
    port map (
            in0 => \N__43315\,
            in1 => \N__39679\,
            in2 => \N__39637\,
            in3 => \N__39634\,
            lcout => \c0.n18_adj_3412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_3_lut_4_lut_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__66631\,
            in1 => \N__53537\,
            in2 => \N__49303\,
            in3 => \N__52672\,
            lcout => \c0.n20300\,
            ltout => \c0.n20300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_350_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49230\,
            in1 => \N__52567\,
            in2 => \N__39610\,
            in3 => \N__57862\,
            lcout => \c0.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_530_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__59688\,
            in1 => \N__49231\,
            in2 => \N__39607\,
            in3 => \N__45935\,
            lcout => \c0.n20370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i186_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__66632\,
            in1 => \N__53702\,
            in2 => \_gnd_net_\,
            in3 => \N__71548\,
            lcout => data_in_frame_23_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71126\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1213_2_lut_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__39576\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42504\,
            lcout => \c0.n3235\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_3_lut_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__64886\,
            in1 => \N__44897\,
            in2 => \_gnd_net_\,
            in3 => \N__48381\,
            lcout => \c0.n40_adj_3374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i133_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__72774\,
            in1 => \N__65598\,
            in2 => \_gnd_net_\,
            in3 => \N__45612\,
            lcout => data_in_frame_16_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71126\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_850_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__41942\,
            in1 => \N__49458\,
            in2 => \N__49785\,
            in3 => \N__53259\,
            lcout => \c0.n17947\,
            ltout => \c0.n17947_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_532_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39703\,
            in2 => \N__39682\,
            in3 => \N__70405\,
            lcout => \c0.n20793\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i227_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__68646\,
            in1 => \N__67178\,
            in2 => \N__59211\,
            in3 => \N__66952\,
            lcout => \c0.data_in_frame_28_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i213_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__72737\,
            in1 => \N__66948\,
            in2 => \N__41949\,
            in3 => \N__62838\,
            lcout => \c0.data_in_frame_26_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_407_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39739\,
            in2 => \_gnd_net_\,
            in3 => \N__39865\,
            lcout => OPEN,
            ltout => \c0.n10_adj_3242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_410_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__43906\,
            in1 => \N__52942\,
            in2 => \N__39670\,
            in3 => \N__39649\,
            lcout => \c0.n11446\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i214_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__62837\,
            in1 => \N__67987\,
            in2 => \N__66977\,
            in3 => \N__49781\,
            lcout => \c0.data_in_frame_26_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_408_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__39844\,
            in1 => \N__39665\,
            in2 => \N__39828\,
            in3 => \N__40025\,
            lcout => \c0.n14_adj_3243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_397_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47006\,
            in2 => \_gnd_net_\,
            in3 => \N__41631\,
            lcout => \c0.n105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__3__5178_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__40026\,
            in1 => \_gnd_net_\,
            in2 => \N__53224\,
            in3 => \N__39868\,
            lcout => data_in_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71158\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__1__5172_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53188\,
            in1 => \N__71505\,
            in2 => \_gnd_net_\,
            in3 => \N__39845\,
            lcout => data_in_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71158\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_916_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__71777\,
            in1 => \N__64393\,
            in2 => \_gnd_net_\,
            in3 => \N__59455\,
            lcout => n19126,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__7__5190_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53187\,
            in1 => \N__39824\,
            in2 => \_gnd_net_\,
            in3 => \N__43942\,
            lcout => data_in_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71158\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_398_LC_17_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__39807\,
            in1 => \N__39914\,
            in2 => \N__39769\,
            in3 => \N__41895\,
            lcout => \c0.n18_adj_3229\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_415_LC_17_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42605\,
            in1 => \N__41927\,
            in2 => \N__49744\,
            in3 => \N__39961\,
            lcout => OPEN,
            ltout => \c0.n21108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_416_LC_17_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39765\,
            in1 => \N__41853\,
            in2 => \N__39754\,
            in3 => \N__39924\,
            lcout => \c0.n12_adj_3248\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_418_LC_17_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__39925\,
            in1 => \N__39745\,
            in2 => \N__52956\,
            in3 => \N__40032\,
            lcout => \c0.n20_adj_3250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__3__5186_LC_17_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40033\,
            in1 => \N__53219\,
            in2 => \_gnd_net_\,
            in3 => \N__40008\,
            lcout => data_in_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__4__5177_LC_17_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53218\,
            in1 => \N__47033\,
            in2 => \_gnd_net_\,
            in3 => \N__43981\,
            lcout => data_in_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__2__5179_LC_17_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__41928\,
            in1 => \N__53220\,
            in2 => \_gnd_net_\,
            in3 => \N__39915\,
            lcout => data_in_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_404_LC_17_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__42604\,
            in1 => \N__47032\,
            in2 => \N__39982\,
            in3 => \N__39960\,
            lcout => \c0.n10_adj_3238\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_adj_412_LC_17_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40573\,
            in2 => \_gnd_net_\,
            in3 => \N__42536\,
            lcout => \c0.n16_adj_3247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_413_LC_17_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__52920\,
            in1 => \N__39940\,
            in2 => \N__39916\,
            in3 => \N__42550\,
            lcout => OPEN,
            ltout => \c0.n20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_414_LC_17_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__41623\,
            in1 => \N__42628\,
            in2 => \N__39934\,
            in3 => \N__39931\,
            lcout => \c0.n11311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__7__5166_LC_17_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53222\,
            in1 => \N__72292\,
            in2 => \_gnd_net_\,
            in3 => \N__41624\,
            lcout => data_in_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71178\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__2__5171_LC_17_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__68644\,
            in1 => \N__53223\,
            in2 => \_gnd_net_\,
            in3 => \N__39913\,
            lcout => data_in_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71178\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__5__5192_LC_17_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53221\,
            in1 => \N__41854\,
            in2 => \_gnd_net_\,
            in3 => \N__40574\,
            lcout => data_in_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71178\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i18_LC_17_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40317\,
            in2 => \_gnd_net_\,
            in3 => \N__40552\,
            lcout => \c0.FRAME_MATCHER_state_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71189\,
            ce => 'H',
            sr => \N__40297\
        );

    \c0.rx.equal_94_i4_2_lut_LC_18_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43870\,
            in2 => \_gnd_net_\,
            in3 => \N__43818\,
            lcout => n4_adj_3579,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_65_i9_2_lut_3_lut_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__60252\,
            in1 => \N__59985\,
            in2 => \_gnd_net_\,
            in3 => \N__60104\,
            lcout => \c0.n9_adj_3025\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i25_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__65147\,
            in1 => \N__61688\,
            in2 => \N__61449\,
            in3 => \N__47598\,
            lcout => \c0.data_in_frame_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71200\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_525_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__40288\,
            in1 => \N__40175\,
            in2 => \N__40118\,
            in3 => \N__49655\,
            lcout => \c0.n12_adj_3265\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_703_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54058\,
            in1 => \N__47596\,
            in2 => \N__47344\,
            in3 => \N__55183\,
            lcout => \c0.n20224\,
            ltout => \c0.n20224_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_274_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40039\,
            in3 => \N__41143\,
            lcout => OPEN,
            ltout => \c0.n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_277_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42649\,
            in1 => \N__40621\,
            in2 => \N__40036\,
            in3 => \N__50076\,
            lcout => \c0.n20246\,
            ltout => \c0.n20246_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_286_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40642\,
            in3 => \N__47259\,
            lcout => \c0.n12_adj_3049\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_810_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61226\,
            in2 => \_gnd_net_\,
            in3 => \N__60411\,
            lcout => \c0.n24_adj_3327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47597\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50604\,
            lcout => \c0.n23_adj_3039\,
            ltout => \c0.n23_adj_3039_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_941_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41002\,
            in1 => \N__42717\,
            in2 => \N__40630\,
            in3 => \N__42690\,
            lcout => \c0.n42_adj_3560\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_275_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40627\,
            in1 => \N__43230\,
            in2 => \N__42718\,
            in3 => \N__41001\,
            lcout => \c0.n30_adj_3042\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i37_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__44117\,
            in1 => \N__61596\,
            in2 => \N__54266\,
            in3 => \N__72612\,
            lcout => \c0.data_in_frame_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__2__5204_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__55185\,
            in1 => \N__46907\,
            in2 => \_gnd_net_\,
            in3 => \N__40614\,
            lcout => data_out_frame_29_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_550_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__49917\,
            in1 => \N__54876\,
            in2 => \_gnd_net_\,
            in3 => \N__42970\,
            lcout => OPEN,
            ltout => \c0.n18428_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_593_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__49828\,
            in1 => \N__44506\,
            in2 => \N__40600\,
            in3 => \N__47911\,
            lcout => \c0.n29_adj_3446\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__2__5212_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111011100100"
        )
    port map (
            in0 => \N__46905\,
            in1 => \N__40591\,
            in2 => \N__46300\,
            in3 => \N__56853\,
            lcout => data_out_frame_28_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__1__5213_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__40957\,
            in1 => \N__46906\,
            in2 => \_gnd_net_\,
            in3 => \N__46287\,
            lcout => data_out_frame_28_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i40_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__44118\,
            in1 => \N__72231\,
            in2 => \N__51282\,
            in3 => \N__61597\,
            lcout => \c0.data_in_frame_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_704_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__51399\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51266\,
            lcout => \c0.n5_adj_3044\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_922_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46283\,
            in1 => \N__42817\,
            in2 => \N__42868\,
            in3 => \N__42823\,
            lcout => \c0.data_out_frame_28__0__N_708\,
            ltout => \c0.data_out_frame_28__0__N_708_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__1__5205_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__50348\,
            in1 => \_gnd_net_\,
            in2 => \N__40984\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_out_frame_29_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71169\,
            ce => \N__46858\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__0__5206_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__55165\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40981\,
            lcout => \c0.data_out_frame_29_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71169\,
            ce => \N__46858\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40963\,
            in1 => \N__40956\,
            in2 => \_gnd_net_\,
            in3 => \N__40926\,
            lcout => \c0.n26_adj_3103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_794_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55163\,
            in2 => \_gnd_net_\,
            in3 => \N__62127\,
            lcout => \c0.n14_adj_3525\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_808_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__62126\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54383\,
            lcout => \c0.n11_adj_3507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_241_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55164\,
            in2 => \_gnd_net_\,
            in3 => \N__54134\,
            lcout => \c0.n12_adj_3015\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_747_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__47545\,
            in1 => \N__54410\,
            in2 => \_gnd_net_\,
            in3 => \N__50554\,
            lcout => \c0.n20209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_4_lut_adj_781_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50496\,
            in1 => \N__54560\,
            in2 => \N__50086\,
            in3 => \N__54423\,
            lcout => \c0.n20204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_2_lut_adj_304_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41124\,
            in2 => \_gnd_net_\,
            in3 => \N__51386\,
            lcout => \c0.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i6_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__61723\,
            in1 => \N__67979\,
            in2 => \N__50582\,
            in3 => \N__55888\,
            lcout => data_in_frame_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71159\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_600_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50641\,
            in2 => \_gnd_net_\,
            in3 => \N__55179\,
            lcout => \c0.n19217\,
            ltout => \c0.n19217_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i33_3_lut_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40995\,
            in2 => \N__41005\,
            in3 => \N__47615\,
            lcout => \c0.n85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i5_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__72649\,
            in1 => \N__55887\,
            in2 => \N__54459\,
            in3 => \N__61724\,
            lcout => data_in_frame_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71159\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_2_lut_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__54411\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47546\,
            lcout => \c0.n66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_adj_601_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47614\,
            in2 => \_gnd_net_\,
            in3 => \N__47547\,
            lcout => \c0.n23_adj_3076\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i1_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41049\,
            in1 => \N__54135\,
            in2 => \_gnd_net_\,
            in3 => \N__41095\,
            lcout => control_mode_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71144\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41038\,
            in1 => \N__55510\,
            in2 => \N__43179\,
            in3 => \N__54733\,
            lcout => \c0.n20321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i26_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__61779\,
            in1 => \N__61448\,
            in2 => \N__50679\,
            in3 => \N__71496\,
            lcout => \c0.data_in_frame_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71144\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_adj_829_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50550\,
            in2 => \_gnd_net_\,
            in3 => \N__54395\,
            lcout => \c0.n15_adj_3543\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i93_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__72677\,
            in1 => \N__64551\,
            in2 => \N__50984\,
            in3 => \N__66050\,
            lcout => \c0.data_in_frame_11_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71144\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i23_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__47548\,
            in1 => \N__68980\,
            in2 => \N__44253\,
            in3 => \N__61780\,
            lcout => \c0.data_in_frame_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71144\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__62255\,
            in1 => \N__47921\,
            in2 => \_gnd_net_\,
            in3 => \N__56650\,
            lcout => \c0.n19176\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_3_lut_4_lut_adj_714_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56651\,
            in1 => \N__41131\,
            in2 => \N__56452\,
            in3 => \N__42672\,
            lcout => OPEN,
            ltout => \c0.n32_adj_3493_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_849_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42901\,
            in1 => \N__61284\,
            in2 => \N__41032\,
            in3 => \N__42933\,
            lcout => OPEN,
            ltout => \c0.n36_adj_3547_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_856_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56703\,
            in1 => \N__54556\,
            in2 => \N__41182\,
            in3 => \N__54442\,
            lcout => OPEN,
            ltout => \c0.n38_adj_3548_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_861_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41179\,
            in1 => \N__41149\,
            in2 => \N__41167\,
            in3 => \N__41164\,
            lcout => \c0.n18443\,
            ltout => \c0.n18443_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_3_lut_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__44734\,
            in1 => \_gnd_net_\,
            in2 => \N__41152\,
            in3 => \N__64633\,
            lcout => \c0.n24_adj_3335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_298_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__50157\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50182\,
            lcout => \c0.n4_adj_3071\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_3_lut_adj_784_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__51338\,
            in1 => \N__50349\,
            in2 => \_gnd_net_\,
            in3 => \N__55052\,
            lcout => \c0.n25_adj_3495\,
            ltout => \c0.n25_adj_3495_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_3_lut_4_lut_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41142\,
            in1 => \N__42671\,
            in2 => \N__41101\,
            in3 => \N__47428\,
            lcout => \c0.n44_adj_3117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i222_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__67920\,
            in1 => \N__64577\,
            in2 => \N__48785\,
            in3 => \N__66962\,
            lcout => \c0.data_in_frame_27_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i137_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__71786\,
            in1 => \N__63354\,
            in2 => \N__48366\,
            in3 => \N__65239\,
            lcout => \c0.data_in_frame_17_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i140_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__63353\,
            in1 => \N__71787\,
            in2 => \N__69444\,
            in3 => \N__68274\,
            lcout => \c0.data_in_frame_17_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i206_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__59719\,
            in1 => \N__63355\,
            in2 => \N__66978\,
            in3 => \N__67919\,
            lcout => \c0.data_in_frame_25_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_588_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44220\,
            in2 => \_gnd_net_\,
            in3 => \N__59480\,
            lcout => \c0.n19134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_819_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43275\,
            in1 => \N__44472\,
            in2 => \N__63575\,
            in3 => \N__58466\,
            lcout => \c0.n20_adj_3539\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_744_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44631\,
            in1 => \N__62418\,
            in2 => \N__44480\,
            in3 => \N__43274\,
            lcout => \c0.n10_adj_3514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__57412\,
            in1 => \N__43126\,
            in2 => \N__47653\,
            in3 => \N__41200\,
            lcout => \c0.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_602_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__62968\,
            in1 => \N__47802\,
            in2 => \_gnd_net_\,
            in3 => \N__61879\,
            lcout => \c0.n6_adj_3453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i129_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__65238\,
            in1 => \N__65595\,
            in2 => \_gnd_net_\,
            in3 => \N__62969\,
            lcout => data_in_frame_16_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i130_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__65594\,
            in1 => \N__71486\,
            in2 => \_gnd_net_\,
            in3 => \N__47803\,
            lcout => data_in_frame_16_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_4_lut_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62890\,
            in1 => \N__47925\,
            in2 => \N__49582\,
            in3 => \N__57045\,
            lcout => \c0.n18_adj_3369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55669\,
            in2 => \_gnd_net_\,
            in3 => \N__52092\,
            lcout => \c0.n17849\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_821_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41254\,
            in1 => \N__44584\,
            in2 => \N__56878\,
            in3 => \N__50113\,
            lcout => \c0.n19474\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_927_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43276\,
            in1 => \N__44479\,
            in2 => \N__41233\,
            in3 => \N__62419\,
            lcout => OPEN,
            ltout => \c0.n12_adj_3001_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_227_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__57152\,
            in1 => \N__44632\,
            in2 => \N__41248\,
            in3 => \N__52275\,
            lcout => \c0.n20403\,
            ltout => \c0.n20403_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_745_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__43277\,
            in1 => \N__48429\,
            in2 => \N__41245\,
            in3 => \N__41216\,
            lcout => OPEN,
            ltout => \c0.n20398_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_746_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__57153\,
            in1 => \N__41242\,
            in2 => \N__41236\,
            in3 => \N__41232\,
            lcout => \c0.n10_adj_3445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_639_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__64769\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__68289\,
            lcout => \c0.n12134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_596_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41217\,
            in1 => \N__45637\,
            in2 => \N__45458\,
            in3 => \N__44633\,
            lcout => \c0.n20_adj_3448\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_2_lut_3_lut_adj_678_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__68374\,
            in1 => \N__52346\,
            in2 => \_gnd_net_\,
            in3 => \N__52171\,
            lcout => \c0.n36_adj_3267\,
            ltout => \c0.n36_adj_3267_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i35_2_lut_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41203\,
            in3 => \N__49068\,
            lcout => \c0.n86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i167_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__69002\,
            in1 => \N__71776\,
            in2 => \N__70125\,
            in3 => \N__67130\,
            lcout => \c0.data_in_frame_20_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i43_4_lut_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49069\,
            in1 => \N__43087\,
            in2 => \N__45051\,
            in3 => \N__44945\,
            lcout => \c0.n94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i143_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__63356\,
            in1 => \N__71775\,
            in2 => \N__69025\,
            in3 => \N__51200\,
            lcout => \c0.data_in_frame_17_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_938_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47830\,
            in2 => \_gnd_net_\,
            in3 => \N__62981\,
            lcout => \c0.n19427\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_944_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65525\,
            in2 => \_gnd_net_\,
            in3 => \N__63774\,
            lcout => \c0.n19187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_231_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48373\,
            in1 => \N__41260\,
            in2 => \N__41605\,
            in3 => \N__43278\,
            lcout => \c0.n19514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_356_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67566\,
            in1 => \N__48595\,
            in2 => \N__47068\,
            in3 => \N__52491\,
            lcout => \c0.n29_adj_3148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_3_lut_adj_905_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44716\,
            in1 => \N__65868\,
            in2 => \_gnd_net_\,
            in3 => \N__47772\,
            lcout => \c0.n17_adj_3451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i220_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__69216\,
            in1 => \N__66881\,
            in2 => \N__48617\,
            in3 => \N__64584\,
            lcout => \c0.data_in_frame_27_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i215_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__62801\,
            in1 => \N__66880\,
            in2 => \N__69023\,
            in3 => \N__43668\,
            lcout => \c0.data_in_frame_26_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i211_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__66879\,
            in1 => \N__68553\,
            in2 => \N__58708\,
            in3 => \N__62802\,
            lcout => \c0.data_in_frame_26_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i151_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__68994\,
            in1 => \N__63939\,
            in2 => \_gnd_net_\,
            in3 => \N__41547\,
            lcout => data_in_frame_18_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i3_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__41529\,
            in1 => \N__69215\,
            in2 => \N__56224\,
            in3 => \N__55467\,
            lcout => rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i152_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__72260\,
            in1 => \N__63938\,
            in2 => \_gnd_net_\,
            in3 => \N__59116\,
            lcout => data_in_frame_18_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71098\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i134_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__65597\,
            in1 => \N__67939\,
            in2 => \_gnd_net_\,
            in3 => \N__45433\,
            lcout => data_in_frame_16_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71098\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_642_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42003\,
            in1 => \N__66500\,
            in2 => \N__59794\,
            in3 => \N__66469\,
            lcout => \c0.n14_adj_3434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i43_4_lut_adj_515_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45052\,
            in1 => \N__49081\,
            in2 => \N__58552\,
            in3 => \N__44946\,
            lcout => \c0.n94_adj_3375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_327_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60346\,
            in2 => \_gnd_net_\,
            in3 => \N__59459\,
            lcout => \c0.n19107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_855_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41495\,
            in2 => \_gnd_net_\,
            in3 => \N__41433\,
            lcout => \c0.n18667\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i28_2_lut_3_lut_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__49079\,
            in1 => \N__43089\,
            in2 => \_gnd_net_\,
            in3 => \N__51808\,
            lcout => \c0.n61\,
            ltout => \c0.n61_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i31_4_lut_adj_303_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41665\,
            in1 => \N__45211\,
            in2 => \N__41668\,
            in3 => \N__45345\,
            lcout => \c0.n64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_300_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__45189\,
            in1 => \N__41973\,
            in2 => \N__48778\,
            in3 => \N__42002\,
            lcout => \c0.n50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i37_4_lut_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__48538\,
            in1 => \N__45346\,
            in2 => \N__45870\,
            in3 => \N__45190\,
            lcout => OPEN,
            ltout => \c0.n86_adj_3393_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i46_4_lut_adj_558_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43303\,
            in1 => \N__41659\,
            in2 => \N__41653\,
            in3 => \N__45306\,
            lcout => OPEN,
            ltout => \c0.n95_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_580_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__58159\,
            in1 => \N__43060\,
            in2 => \N__41650\,
            in3 => \N__43483\,
            lcout => \c0.n15_adj_3441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__7__5174_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42574\,
            in1 => \N__41635\,
            in2 => \_gnd_net_\,
            in3 => \N__53179\,
            lcout => data_in_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i135_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41600\,
            in1 => \N__65590\,
            in2 => \_gnd_net_\,
            in3 => \N__69015\,
            lcout => data_in_frame_16_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i216_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66896\,
            in1 => \N__62803\,
            in2 => \N__45868\,
            in3 => \N__72287\,
            lcout => \c0.data_in_frame_26_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_546_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__41577\,
            in1 => \N__70456\,
            in2 => \_gnd_net_\,
            in3 => \N__70180\,
            lcout => \c0.n20931\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i232_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__72286\,
            in1 => \N__66897\,
            in2 => \N__52794\,
            in3 => \N__67166\,
            lcout => \c0.data_in_frame_28_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i191_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__69014\,
            in1 => \N__53714\,
            in2 => \_gnd_net_\,
            in3 => \N__66496\,
            lcout => data_in_frame_23_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_389_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59332\,
            in2 => \_gnd_net_\,
            in3 => \N__59512\,
            lcout => \c0.n18537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_470_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48829\,
            in1 => \N__52563\,
            in2 => \N__41694\,
            in3 => \N__41722\,
            lcout => \c0.n18_adj_3314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i233_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__41800\,
            in1 => \N__65260\,
            in2 => \N__66976\,
            in3 => \N__71869\,
            lcout => \c0.data_in_frame_29_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i240_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__71868\,
            in1 => \N__72285\,
            in2 => \N__41710\,
            in3 => \N__66947\,
            lcout => \c0.data_in_frame_29_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i239_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__66943\,
            in1 => \N__69022\,
            in2 => \N__41695\,
            in3 => \N__71870\,
            lcout => \c0.data_in_frame_29_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_357_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53263\,
            in1 => \N__53512\,
            in2 => \N__43687\,
            in3 => \N__46095\,
            lcout => OPEN,
            ltout => \c0.n10_adj_3152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_768_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43389\,
            in1 => \N__49507\,
            in2 => \N__41677\,
            in3 => \N__49459\,
            lcout => \c0.n21117\,
            ltout => \c0.n21117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_446_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__41782\,
            in1 => \N__41799\,
            in2 => \N__41791\,
            in3 => \N__43522\,
            lcout => \c0.n40_adj_3282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_351_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__41788\,
            in1 => \N__52423\,
            in2 => \N__49522\,
            in3 => \N__45937\,
            lcout => \c0.n5_adj_3142\,
            ltout => \c0.n5_adj_3142_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_462_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41776\,
            in3 => \N__46003\,
            lcout => OPEN,
            ltout => \c0.n22_adj_3305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_467_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59595\,
            in1 => \N__49346\,
            in2 => \N__41773\,
            in3 => \N__49375\,
            lcout => OPEN,
            ltout => \c0.n37_adj_3309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_adj_479_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46066\,
            in1 => \N__53560\,
            in2 => \N__41770\,
            in3 => \N__43528\,
            lcout => OPEN,
            ltout => \c0.n21099_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_492_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__52519\,
            in1 => \N__48736\,
            in2 => \N__41767\,
            in3 => \N__41764\,
            lcout => OPEN,
            ltout => \c0.n10_adj_3353_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_542_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41740\,
            in1 => \N__43561\,
            in2 => \N__41758\,
            in3 => \N__43702\,
            lcout => \c0.n21111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_490_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__41971\,
            in1 => \N__41998\,
            in2 => \_gnd_net_\,
            in3 => \N__49543\,
            lcout => OPEN,
            ltout => \c0.n9_adj_3352_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_491_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59700\,
            in1 => \N__43555\,
            in2 => \N__41743\,
            in3 => \N__45889\,
            lcout => \c0.n21051\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i224_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__72241\,
            in1 => \N__64565\,
            in2 => \N__42004\,
            in3 => \N__66912\,
            lcout => \c0.data_in_frame_27_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i223_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__41972\,
            in1 => \N__69031\,
            in2 => \N__64578\,
            in3 => \N__66916\,
            lcout => \c0.data_in_frame_27_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i217_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__65242\,
            in1 => \N__64564\,
            in2 => \N__66958\,
            in3 => \N__43385\,
            lcout => \c0.data_in_frame_27_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_454_LC_18_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70382\,
            in1 => \N__70337\,
            in2 => \N__41950\,
            in3 => \N__51862\,
            lcout => \c0.n21003\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i138_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__71734\,
            in1 => \N__63377\,
            in2 => \N__52331\,
            in3 => \N__71506\,
            lcout => \c0.data_in_frame_17_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_405_LC_18_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__41851\,
            in1 => \N__41926\,
            in2 => \_gnd_net_\,
            in3 => \N__41908\,
            lcout => \c0.n110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__7__5182_LC_18_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53209\,
            in1 => \N__42577\,
            in2 => \_gnd_net_\,
            in3 => \N__43941\,
            lcout => data_in_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__5__5184_LC_18_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__41852\,
            in1 => \N__53211\,
            in2 => \_gnd_net_\,
            in3 => \N__41884\,
            lcout => data_in_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_902_LC_18_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__66924\,
            in1 => \N__41833\,
            in2 => \N__55886\,
            in3 => \N__42071\,
            lcout => n20896,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__0__5189_LC_18_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53208\,
            in1 => \N__42640\,
            in2 => \_gnd_net_\,
            in3 => \N__42606\,
            lcout => data_in_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__0__5197_LC_18_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42607\,
            in1 => \N__53210\,
            in2 => \_gnd_net_\,
            in3 => \N__43954\,
            lcout => data_in_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i187_LC_18_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__68645\,
            in1 => \N__53693\,
            in2 => \_gnd_net_\,
            in3 => \N__43410\,
            lcout => data_in_frame_23_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_752_LC_18_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__43924\,
            in1 => \N__43973\,
            in2 => \N__52921\,
            in3 => \N__42576\,
            lcout => \c0.n12_adj_3230\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_402_LC_18_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__43972\,
            in1 => \N__42575\,
            in2 => \_gnd_net_\,
            in3 => \N__43923\,
            lcout => \c0.n11443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i194_LC_18_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46134\,
            in1 => \N__71536\,
            in2 => \_gnd_net_\,
            in3 => \N__70374\,
            lcout => data_in_frame_24_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71191\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__1__5196_LC_18_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53225\,
            in1 => \N__42540\,
            in2 => \_gnd_net_\,
            in3 => \N__43888\,
            lcout => data_in_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71191\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16083_1_lut_2_lut_3_lut_LC_18_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110111011"
        )
    port map (
            in0 => \N__42517\,
            in1 => \N__42370\,
            in2 => \_gnd_net_\,
            in3 => \N__42331\,
            lcout => n1295,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i12201_2_lut_LC_19_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43859\,
            in2 => \_gnd_net_\,
            in3 => \N__43817\,
            lcout => n15645,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_566_LC_19_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__51410\,
            in1 => \N__51331\,
            in2 => \_gnd_net_\,
            in3 => \N__51283\,
            lcout => \c0.n11549\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_322_LC_19_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61874\,
            in2 => \_gnd_net_\,
            in3 => \N__47255\,
            lcout => \c0.n5_adj_3099\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i60_LC_19_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__69436\,
            in1 => \N__64345\,
            in2 => \N__47269\,
            in3 => \N__61685\,
            lcout => \c0.data_in_frame_7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i50_LC_19_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__71374\,
            in1 => \N__61684\,
            in2 => \N__62002\,
            in3 => \N__49906\,
            lcout => \c0.data_in_frame_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i58_LC_19_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__61683\,
            in1 => \N__64344\,
            in2 => \N__63149\,
            in3 => \N__71375\,
            lcout => \c0.data_in_frame_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_3_lut_LC_19_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__63135\,
            in1 => \N__42691\,
            in2 => \_gnd_net_\,
            in3 => \N__63180\,
            lcout => \c0.n31_adj_3121\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_276_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63181\,
            in1 => \N__42673\,
            in2 => \N__63148\,
            in3 => \N__56642\,
            lcout => \c0.n25_adj_3045\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i18_LC_19_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__44215\,
            in1 => \N__61759\,
            in2 => \N__54627\,
            in3 => \N__71348\,
            lcout => \c0.data_in_frame_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71202\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_302_LC_19_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44028\,
            in1 => \N__46390\,
            in2 => \N__47153\,
            in3 => \N__51255\,
            lcout => OPEN,
            ltout => \c0.n14_adj_3073_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_595_LC_19_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46414\,
            in1 => \N__42724\,
            in2 => \N__42643\,
            in3 => \N__42783\,
            lcout => \c0.n4_adj_3009\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_2_lut_LC_19_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51330\,
            in2 => \_gnd_net_\,
            in3 => \N__51257\,
            lcout => \c0.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_294_LC_19_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55213\,
            in2 => \_gnd_net_\,
            in3 => \N__54242\,
            lcout => \c0.n10_adj_3068\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i24_LC_19_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__61758\,
            in1 => \N__44216\,
            in2 => \N__72270\,
            in3 => \N__44157\,
            lcout => \c0.data_in_frame_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71202\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i34_LC_19_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__44119\,
            in1 => \N__61760\,
            in2 => \N__55234\,
            in3 => \N__71349\,
            lcout => \c0.data_in_frame_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71202\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_4_lut_LC_19_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44029\,
            in1 => \N__51256\,
            in2 => \N__50680\,
            in3 => \N__55180\,
            lcout => \c0.n22_adj_3041\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_476_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__54297\,
            in1 => \N__44156\,
            in2 => \N__46345\,
            in3 => \N__42784\,
            lcout => \c0.n21079\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i67_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__55795\,
            in1 => \N__64198\,
            in2 => \N__50149\,
            in3 => \N__68648\,
            lcout => \c0.data_in_frame_8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71193\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_4_lut_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50407\,
            in1 => \N__44155\,
            in2 => \N__50359\,
            in3 => \N__50592\,
            lcout => \c0.n13_adj_3017\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_730_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44382\,
            in1 => \N__54296\,
            in2 => \N__47152\,
            in3 => \N__61073\,
            lcout => \c0.n13_adj_3504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_726_LC_19_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47715\,
            in2 => \_gnd_net_\,
            in3 => \N__49851\,
            lcout => \c0.n6_adj_3501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i4_LC_19_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__61686\,
            in1 => \N__69435\,
            in2 => \N__55819\,
            in3 => \N__62129\,
            lcout => data_in_frame_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71193\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i3_LC_19_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__68647\,
            in1 => \N__55796\,
            in2 => \N__61099\,
            in3 => \N__61687\,
            lcout => data_in_frame_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71193\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_282_LC_19_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44383\,
            in1 => \N__62128\,
            in2 => \_gnd_net_\,
            in3 => \N__54427\,
            lcout => \c0.n11516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_663_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50347\,
            in1 => \N__54422\,
            in2 => \N__50599\,
            in3 => \N__55181\,
            lcout => \c0.n14_adj_3480\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_844_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__61080\,
            in1 => \N__56810\,
            in2 => \N__46292\,
            in3 => \N__62163\,
            lcout => \c0.n13_adj_3546\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_702_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__62164\,
            in1 => \N__55182\,
            in2 => \N__50600\,
            in3 => \N__46273\,
            lcout => OPEN,
            ltout => \c0.n13_adj_3490_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12053_4_lut_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001100"
        )
    port map (
            in0 => \N__42733\,
            in1 => \N__42772\,
            in2 => \N__42766\,
            in3 => \N__42763\,
            lcout => \c0.n15497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_608_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__50346\,
            in1 => \N__54421\,
            in2 => \N__56830\,
            in3 => \N__61079\,
            lcout => \c0.n14_adj_3459\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i1_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__55800\,
            in1 => \N__65240\,
            in2 => \N__46293\,
            in3 => \N__61730\,
            lcout => data_in_frame_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_524_LC_19_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54298\,
            in1 => \N__61078\,
            in2 => \N__56829\,
            in3 => \N__55364\,
            lcout => \c0.n11_adj_3394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_635_LC_19_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56032\,
            in1 => \N__45093\,
            in2 => \N__42844\,
            in3 => \N__47270\,
            lcout => \c0.n10_adj_3207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_adj_743_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__44355\,
            in1 => \_gnd_net_\,
            in2 => \N__42796\,
            in3 => \_gnd_net_\,
            lcout => \c0.n39_adj_3398\,
            ltout => \c0.n39_adj_3398_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_761_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44292\,
            in1 => \N__44280\,
            in2 => \N__42826\,
            in3 => \N__50553\,
            lcout => \c0.n28_adj_3519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_adj_795_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__50551\,
            in1 => \N__56800\,
            in2 => \_gnd_net_\,
            in3 => \N__50317\,
            lcout => \c0.n13_adj_3526\,
            ltout => \c0.n13_adj_3526_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_830_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42816\,
            in1 => \N__42805\,
            in2 => \N__42799\,
            in3 => \N__42874\,
            lcout => \c0.n13_adj_3513\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i45_LC_19_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__61726\,
            in1 => \N__60336\,
            in2 => \N__50023\,
            in3 => \N__72611\,
            lcout => \c0.data_in_frame_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71171\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_adj_790_LC_19_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42792\,
            in2 => \_gnd_net_\,
            in3 => \N__50552\,
            lcout => \c0.n24_adj_3011\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i21_LC_19_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__61725\,
            in1 => \N__44240\,
            in2 => \N__60983\,
            in3 => \N__72610\,
            lcout => \c0.data_in_frame_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71171\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i27_4_lut_adj_727_LC_19_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44293\,
            in1 => \N__44281\,
            in2 => \N__47278\,
            in3 => \N__44272\,
            lcout => \c0.n60_adj_3503\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_552_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__55588\,
            in1 => \N__56299\,
            in2 => \_gnd_net_\,
            in3 => \N__55378\,
            lcout => OPEN,
            ltout => \c0.n16_adj_3416_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_762_LC_19_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42883\,
            in1 => \N__61225\,
            in2 => \N__42877\,
            in3 => \N__50691\,
            lcout => \c0.n20088\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_826_LC_19_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42861\,
            in1 => \N__47217\,
            in2 => \N__47559\,
            in3 => \N__54623\,
            lcout => \c0.n16_adj_3542\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_799_LC_19_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61092\,
            in2 => \_gnd_net_\,
            in3 => \N__54384\,
            lcout => \c0.n5_adj_3528\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i26_2_lut_3_lut_LC_19_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__50639\,
            in1 => \N__44158\,
            in2 => \_gnd_net_\,
            in3 => \N__50566\,
            lcout => \c0.n78\,
            ltout => \c0.n78_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_567_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55509\,
            in1 => \N__50239\,
            in2 => \N__42850\,
            in3 => \N__54130\,
            lcout => \c0.n11800\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_adj_496_LC_19_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__50640\,
            in1 => \N__55585\,
            in2 => \_gnd_net_\,
            in3 => \N__47391\,
            lcout => \c0.n37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62256\,
            in1 => \N__63105\,
            in2 => \N__44634\,
            in3 => \N__56911\,
            lcout => OPEN,
            ltout => \c0.n30_adj_3119_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_334_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__56719\,
            in1 => \N__50108\,
            in2 => \N__42847\,
            in3 => \N__57142\,
            lcout => \c0.n33_adj_3122\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_801_LC_19_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__49879\,
            in1 => \N__62682\,
            in2 => \N__42968\,
            in3 => \N__57307\,
            lcout => \c0.n20055\,
            ltout => \c0.n20055_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_329_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__63843\,
            in1 => \N__62411\,
            in2 => \N__42943\,
            in3 => \N__42926\,
            lcout => OPEN,
            ltout => \c0.n37_adj_3110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63155\,
            in1 => \N__42900\,
            in2 => \N__42904\,
            in3 => \N__56646\,
            lcout => \c0.n43_adj_3116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_807_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__63202\,
            in1 => \_gnd_net_\,
            in2 => \N__63070\,
            in3 => \N__63231\,
            lcout => \c0.n22_adj_3115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i83_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__68593\,
            in1 => \N__66012\,
            in2 => \N__43042\,
            in3 => \N__62793\,
            lcout => \c0.data_in_frame_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_813_LC_19_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44499\,
            in1 => \N__62587\,
            in2 => \N__45022\,
            in3 => \N__57330\,
            lcout => \c0.n23_adj_3534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i84_LC_19_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66011\,
            in1 => \N__62794\,
            in2 => \N__44481\,
            in3 => \N__69408\,
            lcout => \c0.data_in_frame_10_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_886_LC_19_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__62465\,
            in1 => \N__43034\,
            in2 => \_gnd_net_\,
            in3 => \N__44538\,
            lcout => OPEN,
            ltout => \c0.n6_adj_3024_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_245_LC_19_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__56352\,
            in1 => \N__57328\,
            in2 => \N__42889\,
            in3 => \N__62683\,
            lcout => \c0.n18435\,
            ltout => \c0.n18435_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_2_lut_LC_19_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42886\,
            in3 => \N__47684\,
            lcout => \c0.n25_adj_3035\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_adj_887_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57329\,
            in2 => \N__43041\,
            in3 => \N__62466\,
            lcout => \c0.n14_adj_3007\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_929_LC_19_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__65864\,
            in1 => \N__52093\,
            in2 => \N__55671\,
            in3 => \N__43273\,
            lcout => \c0.n17871\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57075\,
            in1 => \N__62467\,
            in2 => \N__44482\,
            in3 => \N__62911\,
            lcout => OPEN,
            ltout => \c0.n28_adj_3120_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_335_LC_19_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43012\,
            in1 => \N__43000\,
            in2 => \N__42991\,
            in3 => \N__42988\,
            lcout => \c0.n20052\,
            ltout => \c0.n20052_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_342_LC_19_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42979\,
            in3 => \N__44804\,
            lcout => OPEN,
            ltout => \c0.n10_adj_3129_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_345_LC_19_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51617\,
            in1 => \N__48068\,
            in2 => \N__42976\,
            in3 => \N__51991\,
            lcout => OPEN,
            ltout => \c0.n18400_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_349_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__45565\,
            in1 => \N__61878\,
            in2 => \N__42973\,
            in3 => \N__57646\,
            lcout => \c0.n13_adj_3139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_3_lut_4_lut_LC_19_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55516\,
            in1 => \N__57371\,
            in2 => \N__51846\,
            in3 => \N__54136\,
            lcout => \c0.n37_adj_3215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_3_lut_4_lut_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55921\,
            in1 => \N__51108\,
            in2 => \N__51847\,
            in3 => \N__50678\,
            lcout => OPEN,
            ltout => \c0.n35_adj_3342_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_4_lut_adj_942_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43237\,
            in1 => \N__43213\,
            in2 => \N__43198\,
            in3 => \N__50082\,
            lcout => OPEN,
            ltout => \c0.n44_adj_3561_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_4_lut_adj_943_LC_19_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43195\,
            in1 => \N__43180\,
            in2 => \N__43156\,
            in3 => \N__43153\,
            lcout => \c0.n21118\,
            ltout => \c0.n21118_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_638_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43120\,
            in1 => \N__57454\,
            in2 => \N__43102\,
            in3 => \N__45182\,
            lcout => \c0.n11_adj_3206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_352_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__57572\,
            in1 => \N__48489\,
            in2 => \N__48032\,
            in3 => \N__43099\,
            lcout => \c0.n20826\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i45_4_lut_adj_556_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45339\,
            in1 => \N__43048\,
            in2 => \N__66532\,
            in3 => \N__45316\,
            lcout => OPEN,
            ltout => \c0.n96_adj_3418_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i48_4_lut_adj_562_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58009\,
            in1 => \N__43088\,
            in2 => \N__43063\,
            in3 => \N__57532\,
            lcout => \c0.n99_adj_3424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i26_3_lut_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__70390\,
            in1 => \N__70264\,
            in2 => \_gnd_net_\,
            in3 => \N__45188\,
            lcout => \c0.n77_adj_3415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_646_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__64003\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58053\,
            lcout => \c0.n10_adj_3474\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_867_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51133\,
            in1 => \N__48260\,
            in2 => \N__51718\,
            in3 => \N__51674\,
            lcout => \c0.n20801\,
            ltout => \c0.n20801_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i45_4_lut_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__43554\,
            in1 => \N__59809\,
            in2 => \N__43321\,
            in3 => \N__45338\,
            lcout => OPEN,
            ltout => \c0.n96_adj_3401_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i48_4_lut_adj_538_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43299\,
            in1 => \N__51807\,
            in2 => \N__43318\,
            in3 => \N__45315\,
            lcout => \c0.n99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i204_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66923\,
            in1 => \N__63394\,
            in2 => \N__49213\,
            in3 => \N__69218\,
            lcout => \c0.data_in_frame_25_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71099\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i148_LC_19_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__69217\,
            in1 => \N__63943\,
            in2 => \_gnd_net_\,
            in3 => \N__64002\,
            lcout => data_in_frame_18_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71099\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_2_lut_adj_641_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67666\,
            in2 => \_gnd_net_\,
            in3 => \N__58037\,
            lcout => \c0.n47_adj_3408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i28_3_lut_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__48177\,
            in1 => \N__44944\,
            in2 => \_gnd_net_\,
            in3 => \N__48860\,
            lcout => \c0.n61_adj_3387\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_2_lut_3_lut_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__55670\,
            in1 => \N__52103\,
            in2 => \_gnd_net_\,
            in3 => \N__43282\,
            lcout => \c0.n43_adj_3386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_2_lut_3_lut_adj_734_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__57723\,
            in1 => \N__48133\,
            in2 => \_gnd_net_\,
            in3 => \N__48654\,
            lcout => \c0.n42_adj_3064\,
            ltout => \c0.n42_adj_3064_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i27_3_lut_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__48103\,
            in1 => \N__45038\,
            in2 => \N__43240\,
            in3 => \_gnd_net_\,
            lcout => \c0.n60_adj_3065\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i178_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__71464\,
            in1 => \N__67522\,
            in2 => \_gnd_net_\,
            in3 => \N__70438\,
            lcout => data_in_frame_22_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i98_LC_19_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66209\,
            in1 => \N__67187\,
            in2 => \N__63853\,
            in3 => \N__71466\,
            lcout => \c0.data_in_frame_12_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12045_2_lut_3_lut_LC_19_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__60274\,
            in1 => \N__60000\,
            in2 => \_gnd_net_\,
            in3 => \N__60132\,
            lcout => \c0.n15489\,
            ltout => \c0.n15489_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i123_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__68691\,
            in1 => \N__43333\,
            in2 => \N__43336\,
            in3 => \N__64221\,
            lcout => \c0.data_in_frame_15_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_234_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45564\,
            in1 => \N__43332\,
            in2 => \_gnd_net_\,
            in3 => \N__48325\,
            lcout => \c0.n19505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i106_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__71465\,
            in1 => \N__48326\,
            in2 => \N__71898\,
            in3 => \N__66210\,
            lcout => \c0.data_in_frame_13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i144_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__71766\,
            in1 => \N__63413\,
            in2 => \N__56524\,
            in3 => \N__72261\,
            lcout => \c0.data_in_frame_17_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_559_LC_19_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__65694\,
            in1 => \N__65797\,
            in2 => \_gnd_net_\,
            in3 => \N__53869\,
            lcout => \c0.n12035\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i181_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53326\,
            in1 => \N__72748\,
            in2 => \_gnd_net_\,
            in3 => \N__67504\,
            lcout => data_in_frame_22_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_716_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70428\,
            in1 => \N__45509\,
            in2 => \N__43420\,
            in3 => \N__53325\,
            lcout => \c0.n12_adj_3494\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__7__5383_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__46886\,
            in1 => \_gnd_net_\,
            in2 => \N__43465\,
            in3 => \N__43434\,
            lcout => data_out_frame_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i188_LC_19_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__69247\,
            in1 => \N__53720\,
            in2 => \_gnd_net_\,
            in3 => \N__45510\,
            lcout => data_in_frame_23_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_534_LC_19_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__43419\,
            in1 => \N__70123\,
            in2 => \N__71284\,
            in3 => \N__53868\,
            lcout => OPEN,
            ltout => \c0.n13_adj_3405_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_535_LC_19_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50908\,
            in1 => \N__45490\,
            in2 => \N__43396\,
            in3 => \N__47980\,
            lcout => \c0.n24_adj_3134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i29_4_lut_adj_497_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__53333\,
            in1 => \N__43641\,
            in2 => \N__43393\,
            in3 => \N__45929\,
            lcout => \c0.n78_adj_3357\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_547_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__65695\,
            in1 => \N__65782\,
            in2 => \N__69607\,
            in3 => \N__53870\,
            lcout => \c0.n17880\,
            ltout => \c0.n17880_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_531_LC_19_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__53755\,
            in1 => \N__69903\,
            in2 => \N__43363\,
            in3 => \N__52130\,
            lcout => \c0.n19342\,
            ltout => \c0.n19342_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_539_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43360\,
            in3 => \N__59738\,
            lcout => \c0.n19496\,
            ltout => \c0.n19496_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_527_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__69517\,
            in1 => \N__43357\,
            in2 => \N__43351\,
            in3 => \N__45930\,
            lcout => \c0.n15_adj_3395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_3_lut_4_lut_adj_627_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59742\,
            in1 => \N__43547\,
            in2 => \N__59692\,
            in3 => \N__48894\,
            lcout => \c0.n32_adj_3095\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_778_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__66382\,
            in1 => \N__66465\,
            in2 => \N__58760\,
            in3 => \N__45825\,
            lcout => \c0.n25_adj_3524\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_465_LC_19_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58726\,
            in1 => \N__45745\,
            in2 => \N__49183\,
            in3 => \N__43695\,
            lcout => OPEN,
            ltout => \c0.n36_adj_3307_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_468_LC_19_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__43520\,
            in1 => \N__52671\,
            in2 => \N__43531\,
            in3 => \N__49302\,
            lcout => \c0.n39_adj_3312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i26_4_lut_adj_500_LC_19_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__43521\,
            in1 => \N__46094\,
            in2 => \N__70338\,
            in3 => \N__43696\,
            lcout => OPEN,
            ltout => \c0.n75_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i44_4_lut_LC_19_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43471\,
            in1 => \N__43495\,
            in2 => \N__43489\,
            in3 => \N__45790\,
            lcout => OPEN,
            ltout => \c0.n93_adj_3373_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i47_4_lut_LC_19_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52774\,
            in1 => \N__43618\,
            in2 => \N__43486\,
            in3 => \N__57790\,
            lcout => \c0.n96_adj_3419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_adj_390_LC_19_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__48838\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49397\,
            lcout => \c0.n23_adj_3222\,
            ltout => \c0.n23_adj_3222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i27_4_lut_adj_498_LC_19_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58725\,
            in1 => \N__59596\,
            in2 => \N__43474\,
            in3 => \N__49178\,
            lcout => \c0.n76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_287_LC_19_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53986\,
            in1 => \N__45270\,
            in2 => \N__43654\,
            in3 => \N__43584\,
            lcout => \c0.n34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_337_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45877\,
            in1 => \N__43677\,
            in2 => \_gnd_net_\,
            in3 => \N__52863\,
            lcout => \c0.n19403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_2_lut_4_lut_LC_19_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__52862\,
            in1 => \N__45876\,
            in2 => \N__43678\,
            in3 => \N__49396\,
            lcout => \c0.n38_adj_3051\,
            ltout => \c0.n38_adj_3051_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_3_lut_adj_448_LC_19_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__43585\,
            in1 => \_gnd_net_\,
            in2 => \N__43645\,
            in3 => \N__49347\,
            lcout => \c0.n45_adj_3284\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_LC_19_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43642\,
            in1 => \N__70279\,
            in2 => \N__45931\,
            in3 => \N__43627\,
            lcout => OPEN,
            ltout => \c0.n51_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i32_4_lut_LC_19_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43617\,
            in1 => \N__43600\,
            in2 => \N__43588\,
            in3 => \N__57789\,
            lcout => \c0.n32_adj_3052\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_4_lut_adj_495_LC_19_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45271\,
            in1 => \N__43576\,
            in2 => \N__43570\,
            in3 => \N__45724\,
            lcout => \c0.n20930\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_461_LC_19_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57255\,
            in1 => \N__52690\,
            in2 => \N__67021\,
            in3 => \N__44788\,
            lcout => \c0.n23_adj_3304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_458_LC_19_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__46096\,
            in1 => \N__59301\,
            in2 => \_gnd_net_\,
            in3 => \N__59250\,
            lcout => OPEN,
            ltout => \c0.n15_adj_3297_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_LC_19_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46207\,
            in1 => \N__49498\,
            in2 => \N__43729\,
            in3 => \N__52843\,
            lcout => \c0.n24_adj_3298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_3_lut_4_lut_LC_19_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__67618\,
            in1 => \N__53473\,
            in2 => \N__59254\,
            in3 => \N__49301\,
            lcout => OPEN,
            ltout => \c0.n21_adj_3300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17661_4_lut_LC_19_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__53556\,
            in1 => \N__43726\,
            in2 => \N__43720\,
            in3 => \N__46042\,
            lcout => OPEN,
            ltout => \c0.n21247_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_494_LC_19_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111101111"
        )
    port map (
            in0 => \N__43717\,
            in1 => \N__52579\,
            in2 => \N__43711\,
            in3 => \N__43708\,
            lcout => \c0.n14_adj_3354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i195_LC_19_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__46135\,
            in1 => \_gnd_net_\,
            in2 => \N__68751\,
            in3 => \N__70209\,
            lcout => data_in_frame_24_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i199_LC_19_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__69013\,
            in1 => \N__46138\,
            in2 => \_gnd_net_\,
            in3 => \N__49505\,
            lcout => data_in_frame_24_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i198_LC_19_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46137\,
            in1 => \N__67972\,
            in2 => \_gnd_net_\,
            in3 => \N__59616\,
            lcout => data_in_frame_24_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i197_LC_19_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__46136\,
            in1 => \_gnd_net_\,
            in2 => \N__72755\,
            in3 => \N__49444\,
            lcout => data_in_frame_24_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i153_LC_19_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__69146\,
            in1 => \N__65217\,
            in2 => \_gnd_net_\,
            in3 => \N__45408\,
            lcout => data_in_frame_19_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__4__5169_LC_19_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__72710\,
            in1 => \N__53226\,
            in2 => \_gnd_net_\,
            in3 => \N__43974\,
            lcout => data_in_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_400_LC_19_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__43953\,
            in1 => \N__43886\,
            in2 => \N__46168\,
            in3 => \N__43940\,
            lcout => \c0.n10_adj_3231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i196_LC_19_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__69421\,
            in1 => \N__46139\,
            in2 => \_gnd_net_\,
            in3 => \N__70324\,
            lcout => data_in_frame_24_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__1__5188_LC_19_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53227\,
            in1 => \N__43915\,
            in2 => \_gnd_net_\,
            in3 => \N__43887\,
            lcout => data_in_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71213\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_98_i4_2_lut_LC_20_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43869\,
            in2 => \_gnd_net_\,
            in3 => \N__43819\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i17_LC_20_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__44233\,
            in1 => \N__61731\,
            in2 => \N__47216\,
            in3 => \N__65094\,
            lcout => \c0.data_in_frame_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i5_LC_20_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__43744\,
            in1 => \N__67777\,
            in2 => \N__56239\,
            in3 => \N__55466\,
            lcout => rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i1_LC_20_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__43755\,
            in1 => \N__71347\,
            in2 => \N__56237\,
            in3 => \N__55465\,
            lcout => rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i4_LC_20_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__43743\,
            in1 => \N__72531\,
            in2 => \N__56238\,
            in3 => \N__56086\,
            lcout => rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_526_LC_20_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60927\,
            in1 => \N__49975\,
            in2 => \N__44423\,
            in3 => \N__55382\,
            lcout => \c0.n19424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_529_LC_20_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__49974\,
            in1 => \N__44413\,
            in2 => \_gnd_net_\,
            in3 => \N__60926\,
            lcout => \c0.n8_adj_3397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i31_LC_20_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__69035\,
            in1 => \N__61430\,
            in2 => \N__44424\,
            in3 => \N__61673\,
            lcout => \c0.data_in_frame_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_773_LC_20_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56825\,
            in2 => \_gnd_net_\,
            in3 => \N__61081\,
            lcout => \c0.n9_adj_3346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_LC_20_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63854\,
            in1 => \N__47768\,
            in2 => \N__64453\,
            in3 => \N__52107\,
            lcout => \c0.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i39_LC_20_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__61671\,
            in1 => \N__44126\,
            in2 => \N__44047\,
            in3 => \N__69036\,
            lcout => \c0.data_in_frame_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i22_LC_20_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__67776\,
            in1 => \N__61672\,
            in2 => \N__44395\,
            in3 => \N__44252\,
            lcout => \c0.data_in_frame_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i35_LC_20_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__61670\,
            in1 => \N__44125\,
            in2 => \N__68758\,
            in3 => \N__46393\,
            lcout => \c0.data_in_frame_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_705_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46391\,
            in1 => \N__55212\,
            in2 => \N__46288\,
            in3 => \N__54612\,
            lcout => \c0.n7_adj_3491\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_772_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__54613\,
            in1 => \N__46416\,
            in2 => \_gnd_net_\,
            in3 => \N__46265\,
            lcout => \c0.n9_adj_3027\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i33_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__65198\,
            in1 => \N__61691\,
            in2 => \N__44128\,
            in3 => \N__49980\,
            lcout => \c0.data_in_frame_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i36_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__61689\,
            in1 => \N__69424\,
            in2 => \N__46420\,
            in3 => \N__44124\,
            lcout => \c0.data_in_frame_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i20_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__69423\,
            in1 => \N__61690\,
            in2 => \N__54316\,
            in3 => \N__44248\,
            lcout => \c0.data_in_frame_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_adj_545_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44151\,
            in1 => \N__62131\,
            in2 => \N__44393\,
            in3 => \N__54466\,
            lcout => \c0.n4_adj_3406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i38_LC_20_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__44120\,
            in1 => \N__67802\,
            in2 => \N__47155\,
            in3 => \N__61692\,
            lcout => \c0.data_in_frame_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_733_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44030\,
            in1 => \N__44005\,
            in2 => \N__43993\,
            in3 => \N__56801\,
            lcout => \c0.data_out_frame_0__7__N_1537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_785_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60956\,
            in1 => \N__62130\,
            in2 => \_gnd_net_\,
            in3 => \N__61077\,
            lcout => \c0.n12131\,
            ltout => \c0.n12131_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_adj_536_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47297\,
            in2 => \N__43984\,
            in3 => \N__62197\,
            lcout => \c0.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i2_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__56823\,
            in1 => \N__61801\,
            in2 => \N__55868\,
            in3 => \N__71393\,
            lcout => data_in_frame_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_786_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44304\,
            in2 => \_gnd_net_\,
            in3 => \N__62198\,
            lcout => \c0.n19415\,
            ltout => \c0.n19415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i36_2_lut_4_lut_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47298\,
            in1 => \N__55032\,
            in2 => \N__44284\,
            in3 => \N__55308\,
            lcout => \c0.n88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_4_lut_adj_736_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55033\,
            in1 => \N__54122\,
            in2 => \N__55309\,
            in3 => \N__47299\,
            lcout => \c0.n54_adj_3502\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_361_LC_20_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__61860\,
            in1 => \N__56629\,
            in2 => \N__62698\,
            in3 => \N__55732\,
            lcout => \c0.n21_adj_3205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i38_4_lut_LC_20_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47336\,
            in1 => \N__60957\,
            in2 => \N__62080\,
            in3 => \N__62199\,
            lcout => \c0.n90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i44_3_lut_4_lut_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54888\,
            in1 => \N__44271\,
            in2 => \N__44571\,
            in3 => \N__44658\,
            lcout => \c0.n96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_791_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46334\,
            in1 => \N__46269\,
            in2 => \_gnd_net_\,
            in3 => \N__56802\,
            lcout => \c0.n20095\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i31_4_lut_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56803\,
            in1 => \N__54492\,
            in2 => \N__55178\,
            in3 => \N__54267\,
            lcout => \c0.n83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_4_lut_LC_20_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54452\,
            in1 => \N__62156\,
            in2 => \N__50406\,
            in3 => \N__55147\,
            lcout => \c0.n14_adj_3371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_818_LC_20_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47619\,
            in3 => \N__54054\,
            lcout => \c0.n10_adj_3538\,
            ltout => \c0.n10_adj_3538_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_822_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44431\,
            in1 => \N__44425\,
            in2 => \N__44398\,
            in3 => \N__44394\,
            lcout => \c0.n22_adj_3356\,
            ltout => \c0.n22_adj_3356_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_2_lut_3_lut_LC_20_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54887\,
            in2 => \N__44359\,
            in3 => \N__47454\,
            lcout => \c0.n52_adj_3402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47370\,
            in1 => \N__44329\,
            in2 => \N__44344\,
            in3 => \N__44641\,
            lcout => \c0.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_adj_832_LC_20_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54880\,
            in2 => \_gnd_net_\,
            in3 => \N__44356\,
            lcout => \c0.n23_adj_3021\,
            ltout => \c0.n23_adj_3021_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_2_lut_4_lut_LC_20_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50673\,
            in1 => \N__55587\,
            in2 => \N__44335\,
            in3 => \N__44654\,
            lcout => \c0.n26_adj_3114\,
            ltout => \c0.n26_adj_3114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_332_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49951\,
            in1 => \N__47369\,
            in2 => \N__44332\,
            in3 => \N__44517\,
            lcout => \c0.n20981\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_758_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__57655\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57571\,
            lcout => \c0.n12_adj_3518\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_270_LC_20_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55263\,
            in1 => \N__60451\,
            in2 => \N__50158\,
            in3 => \N__55239\,
            lcout => \c0.n20490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_237_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50457\,
            in1 => \N__44328\,
            in2 => \N__55291\,
            in3 => \N__44320\,
            lcout => \c0.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_LC_20_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__55586\,
            in1 => \_gnd_net_\,
            in2 => \N__44659\,
            in3 => \N__50672\,
            lcout => \c0.n22_adj_3022\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_879_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__44972\,
            in1 => \_gnd_net_\,
            in2 => \N__51519\,
            in3 => \N__60778\,
            lcout => \c0.n11_adj_3340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_adj_514_LC_20_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__45015\,
            in1 => \_gnd_net_\,
            in2 => \N__44635\,
            in3 => \N__44970\,
            lcout => \c0.n18_adj_3372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_2_lut_3_lut_adj_616_LC_20_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__44971\,
            in1 => \_gnd_net_\,
            in2 => \N__44904\,
            in3 => \N__45016\,
            lcout => \c0.n33_adj_3289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_LC_20_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44572\,
            in1 => \N__47356\,
            in2 => \N__44554\,
            in3 => \N__50461\,
            lcout => \c0.n20029\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_766_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47350\,
            in1 => \N__44527\,
            in2 => \N__44521\,
            in3 => \N__47374\,
            lcout => \c0.n18422\,
            ltout => \c0.n18422_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_272_LC_20_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__62583\,
            in1 => \_gnd_net_\,
            in2 => \N__44488\,
            in3 => \N__57308\,
            lcout => \c0.n19433\,
            ltout => \c0.n19433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_273_LC_20_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__44485\,
            in3 => \N__45014\,
            lcout => OPEN,
            ltout => \c0.n11891_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_288_LC_20_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__44465\,
            in1 => \N__50109\,
            in2 => \N__44434\,
            in3 => \N__57143\,
            lcout => \c0.n20151\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_4_lut_LC_20_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44752\,
            in1 => \N__44743\,
            in2 => \N__47508\,
            in3 => \N__47629\,
            lcout => \c0.n27_adj_3118\,
            ltout => \c0.n27_adj_3118_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_2_lut_3_lut_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48279\,
            in2 => \N__44737\,
            in3 => \N__51942\,
            lcout => \c0.n28_adj_3245\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_505_LC_20_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__48033\,
            in1 => \N__44730\,
            in2 => \_gnd_net_\,
            in3 => \N__56561\,
            lcout => \c0.n19_adj_3336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i87_LC_20_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66156\,
            in1 => \N__62812\,
            in2 => \N__66336\,
            in3 => \N__68903\,
            lcout => \c0.data_in_frame_10_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71146\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_2_lut_4_lut_adj_898_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52040\,
            in1 => \N__60771\,
            in2 => \N__51518\,
            in3 => \N__44969\,
            lcout => \c0.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_adj_611_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__56562\,
            in1 => \N__44719\,
            in2 => \_gnd_net_\,
            in3 => \N__48034\,
            lcout => \c0.n23_adj_3364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_315_LC_20_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__57191\,
            in1 => \_gnd_net_\,
            in2 => \N__65863\,
            in3 => \N__47745\,
            lcout => \c0.n19372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_LC_20_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__51154\,
            in1 => \N__56451\,
            in2 => \N__65350\,
            in3 => \N__51673\,
            lcout => \c0.n19916\,
            ltout => \c0.n19916_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_2_lut_3_lut_LC_20_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__44671\,
            in1 => \N__44805\,
            in2 => \N__44662\,
            in3 => \_gnd_net_\,
            lcout => \c0.n22_adj_3341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_4_lut_LC_20_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64628\,
            in1 => \N__65853\,
            in2 => \N__48219\,
            in3 => \N__48261\,
            lcout => \c0.n21_adj_3337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_831_LC_20_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50739\,
            in1 => \N__56743\,
            in2 => \N__50784\,
            in3 => \N__44827\,
            lcout => \c0.n19477\,
            ltout => \c0.n19477_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_LC_20_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__63049\,
            in1 => \N__56450\,
            in2 => \N__44818\,
            in3 => \N__51672\,
            lcout => OPEN,
            ltout => \c0.n12_adj_3348_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_659_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65343\,
            in1 => \N__57443\,
            in2 => \N__44815\,
            in3 => \N__47887\,
            lcout => \c0.n21045\,
            ltout => \c0.n21045_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_adj_640_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__44812\,
            in3 => \N__52758\,
            lcout => \c0.n19_adj_3303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_3_lut_adj_875_LC_20_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60793\,
            in1 => \N__44979\,
            in2 => \_gnd_net_\,
            in3 => \N__44809\,
            lcout => \c0.n40_adj_3366\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i177_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__65262\,
            in1 => \N__67530\,
            in2 => \_gnd_net_\,
            in3 => \N__70037\,
            lcout => data_in_frame_22_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_645_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49136\,
            in1 => \N__44775\,
            in2 => \N__57235\,
            in3 => \N__52722\,
            lcout => \c0.n20085\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__44764\,
            in1 => \N__55668\,
            in2 => \N__45069\,
            in3 => \N__48510\,
            lcout => \c0.n21110\,
            ltout => \c0.n21110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_654_LC_20_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__45154\,
            in1 => \N__45142\,
            in2 => \N__45100\,
            in3 => \N__45097\,
            lcout => \c0.n40_adj_3413\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i113_LC_20_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__65263\,
            in1 => \N__64238\,
            in2 => \N__62048\,
            in3 => \N__57225\,
            lcout => \c0.data_in_frame_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i116_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__64237\,
            in1 => \N__62035\,
            in2 => \N__45070\,
            in3 => \N__69315\,
            lcout => \c0.data_in_frame_14_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_2_lut_3_lut_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__44986\,
            in1 => \_gnd_net_\,
            in2 => \N__64014\,
            in3 => \N__45021\,
            lcout => \c0.n67_adj_3063\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_3_lut_4_lut_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45020\,
            in1 => \N__44985\,
            in2 => \N__44947\,
            in3 => \N__48933\,
            lcout => \c0.n43_adj_3330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_755_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64833\,
            in2 => \_gnd_net_\,
            in3 => \N__67378\,
            lcout => OPEN,
            ltout => \c0.n12_adj_3517_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_765_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57709\,
            in1 => \N__44920\,
            in2 => \N__44908\,
            in3 => \N__69082\,
            lcout => \c0.n20512\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_665_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__45702\,
            in1 => \N__53414\,
            in2 => \N__44905\,
            in3 => \N__45577\,
            lcout => \c0.n20840\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_847_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44848\,
            in1 => \N__51912\,
            in2 => \N__44839\,
            in3 => \N__52053\,
            lcout => \c0.n20451\,
            ltout => \c0.n20451_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_4_lut_adj_569_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69080\,
            in1 => \N__64832\,
            in2 => \N__45253\,
            in3 => \N__45810\,
            lcout => \c0.n15_adj_3432\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_387_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67379\,
            in1 => \N__45250\,
            in2 => \N__45814\,
            in3 => \N__69081\,
            lcout => \c0.n13_adj_3221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i31_4_lut_adj_738_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48869\,
            in1 => \N__49098\,
            in2 => \N__48102\,
            in3 => \N__57511\,
            lcout => \c0.n64_adj_3512\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_870_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57455\,
            in2 => \_gnd_net_\,
            in3 => \N__45179\,
            lcout => OPEN,
            ltout => \c0.n27_adj_3529_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_802_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__45238\,
            in1 => \N__62950\,
            in2 => \N__45220\,
            in3 => \N__51685\,
            lcout => OPEN,
            ltout => \c0.n32_adj_3530_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_811_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47941\,
            in1 => \N__47704\,
            in2 => \N__45217\,
            in3 => \N__56470\,
            lcout => \c0.n19244\,
            ltout => \c0.n19244_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_2_lut_3_lut_LC_20_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__45290\,
            in1 => \_gnd_net_\,
            in2 => \N__45214\,
            in3 => \N__67657\,
            lcout => \c0.n85_adj_3074\,
            ltout => \c0.n85_adj_3074_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_650_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__45334\,
            in1 => \N__45180\,
            in2 => \N__45199\,
            in3 => \N__45196\,
            lcout => \c0.n13_adj_3244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_3_lut_4_lut_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45181\,
            in1 => \N__47834\,
            in2 => \N__57460\,
            in3 => \N__51687\,
            lcout => \c0.n49_adj_3358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_2_lut_adj_644_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__51686\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57456\,
            lcout => \c0.n49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_788_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63994\,
            in1 => \N__67288\,
            in2 => \N__67434\,
            in3 => \N__51885\,
            lcout => \c0.n30_adj_3392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_2_lut_3_lut_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__65520\,
            in1 => \N__47835\,
            in2 => \_gnd_net_\,
            in3 => \N__59074\,
            lcout => \c0.n48_adj_3409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_775_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__72474\,
            in1 => \_gnd_net_\,
            in2 => \N__66421\,
            in3 => \_gnd_net_\,
            lcout => \c0.n4_adj_3522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i168_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__71791\,
            in1 => \N__70147\,
            in2 => \N__67219\,
            in3 => \N__72221\,
            lcout => \c0.data_in_frame_20_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__59075\,
            in1 => \N__65521\,
            in2 => \_gnd_net_\,
            in3 => \N__58024\,
            lcout => \c0.n22_adj_3287\,
            ltout => \c0.n22_adj_3287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_895_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__67289\,
            in1 => \N__63995\,
            in2 => \N__45274\,
            in3 => \N__57547\,
            lcout => \c0.n10_adj_3555\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_672_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__70126\,
            in1 => \_gnd_net_\,
            in2 => \N__70154\,
            in3 => \_gnd_net_\,
            lcout => \c0.n19223\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_2_lut_3_lut_adj_869_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__68165\,
            in1 => \N__66417\,
            in2 => \_gnd_net_\,
            in3 => \N__72475\,
            lcout => \c0.n39_adj_3050\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_4_lut_adj_560_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__57656\,
            in1 => \N__59126\,
            in2 => \N__57724\,
            in3 => \N__57581\,
            lcout => \c0.n14_adj_3421\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_591_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45638\,
            in2 => \_gnd_net_\,
            in3 => \N__45704\,
            lcout => \c0.n19384\,
            ltout => \c0.n19384_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_621_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__45484\,
            in1 => \N__45475\,
            in2 => \N__45463\,
            in3 => \N__45661\,
            lcout => \c0.n17819\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_4_lut_LC_20_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__64892\,
            in1 => \N__48377\,
            in2 => \N__45452\,
            in3 => \N__45703\,
            lcout => \c0.n9_adj_3430\,
            ltout => \c0.n9_adj_3430_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_590_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45412\,
            in1 => \N__45366\,
            in2 => \N__45394\,
            in3 => \N__45390\,
            lcout => \c0.n20431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_751_LC_20_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__45391\,
            in1 => \N__45376\,
            in2 => \N__45370\,
            in3 => \N__59345\,
            lcout => \c0.n18433\,
            ltout => \c0.n18433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_474_LC_20_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__53907\,
            in1 => \N__66381\,
            in2 => \N__45358\,
            in3 => \N__67639\,
            lcout => \c0.n40_adj_3323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_710_LC_20_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__57582\,
            in1 => \N__57713\,
            in2 => \_gnd_net_\,
            in3 => \N__57657\,
            lcout => \c0.n20479\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_632_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__45355\,
            in1 => \N__53963\,
            in2 => \N__45639\,
            in3 => \N__45713\,
            lcout => \c0.n4_adj_3123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_661_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__59073\,
            in1 => \_gnd_net_\,
            in2 => \N__63777\,
            in3 => \_gnd_net_\,
            lcout => \c0.n19511\,
            ltout => \c0.n19511_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_adj_633_LC_20_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45633\,
            in1 => \N__58839\,
            in2 => \N__45718\,
            in3 => \N__45714\,
            lcout => \c0.n7_adj_3054\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i193_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__65248\,
            in1 => \N__46153\,
            in2 => \_gnd_net_\,
            in3 => \N__58756\,
            lcout => data_in_frame_24_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71160\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_597_LC_20_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__57658\,
            in1 => \N__45673\,
            in2 => \N__65281\,
            in3 => \N__45660\,
            lcout => \c0.n22_adj_3450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i32_4_lut_adj_740_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45649\,
            in1 => \N__58084\,
            in2 => \N__59149\,
            in3 => \N__48544\,
            lcout => \c0.n21071\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_579_LC_20_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45629\,
            in1 => \N__63767\,
            in2 => \_gnd_net_\,
            in3 => \N__59072\,
            lcout => \c0.n7_adj_3440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i105_LC_20_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__65249\,
            in1 => \N__71965\,
            in2 => \N__66211\,
            in3 => \N__45560\,
            lcout => \c0.data_in_frame_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71160\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_388_LC_20_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__68434\,
            in1 => \N__69835\,
            in2 => \N__45541\,
            in3 => \N__45523\,
            lcout => \c0.n18431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_637_LC_20_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__71283\,
            in1 => \N__45514\,
            in2 => \N__69907\,
            in3 => \N__52444\,
            lcout => \c0.n20324\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_3_lut_LC_20_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46177\,
            in1 => \N__48534\,
            in2 => \_gnd_net_\,
            in3 => \N__45496\,
            lcout => \c0.n21044\,
            ltout => \c0.n21044_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_328_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__53602\,
            in1 => \N__47098\,
            in2 => \N__45880\,
            in3 => \N__58761\,
            lcout => OPEN,
            ltout => \c0.n16_adj_3109_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_333_LC_20_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__45869\,
            in1 => \N__49411\,
            in2 => \N__45829\,
            in3 => \N__45826\,
            lcout => \c0.n21076\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_585_LC_20_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64830\,
            in2 => \_gnd_net_\,
            in3 => \N__45804\,
            lcout => \c0.n9_adj_3069\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i28_4_lut_adj_499_LC_20_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49765\,
            in1 => \N__47086\,
            in2 => \N__49348\,
            in3 => \N__49371\,
            lcout => \c0.n77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_320_LC_20_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45784\,
            in1 => \N__45765\,
            in2 => \N__51759\,
            in3 => \N__49017\,
            lcout => \c0.n18457\,
            ltout => \c0.n18457_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_445_LC_20_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52646\,
            in1 => \N__53586\,
            in2 => \N__45748\,
            in3 => \N__46053\,
            lcout => \c0.n41_adj_3281\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_444_LC_20_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59833\,
            in1 => \N__52599\,
            in2 => \N__53824\,
            in3 => \N__45744\,
            lcout => OPEN,
            ltout => \c0.n43_adj_3280_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_4_lut_adj_447_LC_20_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53442\,
            in1 => \N__49354\,
            in2 => \N__45733\,
            in3 => \N__45730\,
            lcout => \c0.n50_adj_3283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_466_LC_20_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__46102\,
            in1 => \N__46093\,
            in2 => \N__46057\,
            in3 => \N__52647\,
            lcout => \c0.n33_adj_3308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_318_LC_20_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49491\,
            in1 => \N__52864\,
            in2 => \N__46206\,
            in3 => \N__52689\,
            lcout => \c0.n18417\,
            ltout => \c0.n18417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_453_LC_20_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46035\,
            in1 => \N__48619\,
            in2 => \N__46045\,
            in3 => \N__52651\,
            lcout => \c0.n19_adj_3292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i237_LC_20_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__72744\,
            in1 => \N__46036\,
            in2 => \N__66975\,
            in3 => \N__71934\,
            lcout => \c0.data_in_frame_29_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i235_LC_20_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__71932\,
            in1 => \N__68744\,
            in2 => \N__46023\,
            in3 => \N__66942\,
            lcout => \c0.data_in_frame_29_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i234_LC_20_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__71534\,
            in1 => \N__45999\,
            in2 => \N__66974\,
            in3 => \N__71933\,
            lcout => \c0.data_in_frame_29_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i226_LC_20_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__45975\,
            in1 => \N__71535\,
            in2 => \N__67222\,
            in3 => \N__66941\,
            lcout => \c0.data_in_frame_28_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i225_LC_20_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66934\,
            in1 => \N__67200\,
            in2 => \N__45955\,
            in3 => \N__65261\,
            lcout => \c0.data_in_frame_28_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_486_LC_20_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__59560\,
            in1 => \N__53842\,
            in2 => \N__45954\,
            in3 => \N__45936\,
            lcout => \c0.n14_adj_3349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_308_LC_20_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49326\,
            in2 => \_gnd_net_\,
            in3 => \N__53383\,
            lcout => \c0.n7_adj_3078\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i136_LC_20_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__72294\,
            in1 => \N__65596\,
            in2 => \_gnd_net_\,
            in3 => \N__57692\,
            lcout => data_in_frame_16_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i141_LC_20_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__71762\,
            in1 => \N__63358\,
            in2 => \N__64760\,
            in3 => \N__72729\,
            lcout => \c0.data_in_frame_17_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i203_LC_20_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__68740\,
            in1 => \N__49259\,
            in2 => \N__63389\,
            in3 => \N__66973\,
            lcout => \c0.data_in_frame_25_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_776_LC_20_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46189\,
            in1 => \N__53942\,
            in2 => \N__72397\,
            in3 => \N__53974\,
            lcout => \c0.n26_adj_3523\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i202_LC_20_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__49327\,
            in1 => \N__71543\,
            in2 => \N__63390\,
            in3 => \N__66972\,
            lcout => \c0.data_in_frame_25_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_540_LC_20_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59612\,
            in2 => \_gnd_net_\,
            in3 => \N__49435\,
            lcout => \c0.n11865\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__4__5193_LC_20_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53229\,
            in1 => \N__46993\,
            in2 => \_gnd_net_\,
            in3 => \N__46167\,
            lcout => data_in_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71215\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3848_2_lut_LC_20_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49487\,
            in2 => \_gnd_net_\,
            in3 => \N__53618\,
            lcout => \c0.n6495\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i200_LC_20_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__53622\,
            in1 => \N__46152\,
            in2 => \_gnd_net_\,
            in3 => \N__72291\,
            lcout => data_in_frame_24_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71215\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_543_LC_20_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__70375\,
            in1 => \N__70314\,
            in2 => \_gnd_net_\,
            in3 => \N__70208\,
            lcout => \c0.n12085\,
            ltout => \c0.n12085_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_787_LC_20_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47082\,
            in2 => \N__47071\,
            in3 => \N__47052\,
            lcout => \c0.n19274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__4__5185_LC_20_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53228\,
            in1 => \N__46992\,
            in2 => \_gnd_net_\,
            in3 => \N__47041\,
            lcout => data_in_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_223_LC_21_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__51015\,
            in1 => \N__54750\,
            in2 => \_gnd_net_\,
            in3 => \N__50989\,
            lcout => \c0.n19291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__7__5207_LC_21_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__46963\,
            in1 => \N__62176\,
            in2 => \N__55186\,
            in3 => \N__50339\,
            lcout => \c0.data_out_frame_28_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71225\,
            ce => \N__46936\,
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_717_LC_21_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46415\,
            in1 => \N__46392\,
            in2 => \N__46368\,
            in3 => \N__47205\,
            lcout => OPEN,
            ltout => \c0.n13_adj_3496_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_721_LC_21_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46213\,
            in1 => \N__49692\,
            in2 => \N__46348\,
            in3 => \N__46341\,
            lcout => \c0.n5_adj_3031\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_713_LC_21_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46301\,
            in2 => \_gnd_net_\,
            in3 => \N__56824\,
            lcout => \c0.n19277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_777_LC_21_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49691\,
            in1 => \N__47206\,
            in2 => \N__47182\,
            in3 => \N__55383\,
            lcout => \c0.n20391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_780_LC_21_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60450\,
            in1 => \N__51054\,
            in2 => \_gnd_net_\,
            in3 => \N__55235\,
            lcout => \c0.n11833\,
            ltout => \c0.n11833_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i40_4_lut_LC_21_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__66287\,
            in1 => \N__47167\,
            in2 => \N__47173\,
            in3 => \N__47116\,
            lcout => OPEN,
            ltout => \c0.n92_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i46_4_lut_LC_21_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47161\,
            in1 => \N__50230\,
            in2 => \N__47170\,
            in3 => \N__62165\,
            lcout => \c0.n98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i28_4_lut_LC_21_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49847\,
            in1 => \N__56378\,
            in2 => \N__49875\,
            in3 => \N__54518\,
            lcout => \c0.n80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_692_LC_21_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50332\,
            in2 => \_gnd_net_\,
            in3 => \N__50405\,
            lcout => \c0.n19196\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_836_LC_21_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49979\,
            in2 => \_gnd_net_\,
            in3 => \N__61197\,
            lcout => \c0.n5_adj_3030\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_792_LC_21_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__54262\,
            in1 => \_gnd_net_\,
            in2 => \N__47154\,
            in3 => \_gnd_net_\,
            lcout => \c0.n19241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_900_LC_21_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__62582\,
            in1 => \N__47145\,
            in2 => \_gnd_net_\,
            in3 => \N__54261\,
            lcout => \c0.n54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i51_4_lut_LC_21_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47110\,
            in1 => \N__49990\,
            in2 => \N__47404\,
            in3 => \N__47104\,
            lcout => \c0.n12_adj_3034\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_2_lut_adj_840_LC_21_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__54094\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61194\,
            lcout => \c0.n24_adj_3013\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i66_LC_21_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__64255\,
            in1 => \N__55883\,
            in2 => \N__51520\,
            in3 => \N__71376\,
            lcout => \c0.data_in_frame_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71205\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_604_LC_21_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__50301\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55034\,
            lcout => \c0.n7_adj_3029\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_adj_551_LC_21_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61196\,
            in1 => \N__54096\,
            in2 => \N__50434\,
            in3 => \N__50300\,
            lcout => \c0.n20313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17690_4_lut_LC_21_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__54097\,
            in1 => \N__50602\,
            in2 => \N__60988\,
            in3 => \N__61118\,
            lcout => \c0.n21277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_4_lut_adj_652_LC_21_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61195\,
            in1 => \N__54095\,
            in2 => \N__54894\,
            in3 => \N__54674\,
            lcout => OPEN,
            ltout => \c0.n14_adj_3476_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_701_LC_21_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50601\,
            in1 => \N__47296\,
            in2 => \N__47281\,
            in3 => \N__55284\,
            lcout => \c0.n19966\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_306_LC_21_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55610\,
            in1 => \N__47227\,
            in2 => \N__50005\,
            in3 => \N__47274\,
            lcout => \c0.n30_adj_3075\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_305_LC_21_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55919\,
            in2 => \_gnd_net_\,
            in3 => \N__51097\,
            lcout => \c0.n19508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_4_lut_adj_833_LC_21_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51287\,
            in1 => \N__55127\,
            in2 => \N__51414\,
            in3 => \N__47476\,
            lcout => \c0.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_2_lut_LC_21_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60488\,
            in2 => \_gnd_net_\,
            in3 => \N__56291\,
            lcout => OPEN,
            ltout => \c0.n67_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i48_4_lut_LC_21_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47470\,
            in1 => \N__47461\,
            in2 => \N__47443\,
            in3 => \N__47440\,
            lcout => OPEN,
            ltout => \c0.n100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i50_4_lut_LC_21_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47434\,
            in1 => \N__47424\,
            in2 => \N__47407\,
            in3 => \N__49930\,
            lcout => \c0.n102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_236_LC_21_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56290\,
            in2 => \_gnd_net_\,
            in3 => \N__47395\,
            lcout => \c0.n21_adj_3010\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_3_lut_4_lut_adj_624_LC_21_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50175\,
            in1 => \N__54531\,
            in2 => \N__60493\,
            in3 => \N__54727\,
            lcout => \c0.n28_adj_3023\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_735_LC_21_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__54532\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__60492\,
            lcout => \c0.n17_adj_3508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i89_LC_21_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__64502\,
            in1 => \N__66154\,
            in2 => \N__53657\,
            in3 => \N__65202\,
            lcout => \c0.data_in_frame_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_307_LC_21_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47340\,
            in1 => \N__54461\,
            in2 => \N__54567\,
            in3 => \N__47317\,
            lcout => OPEN,
            ltout => \c0.n32_adj_3077_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_314_LC_21_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50486\,
            in1 => \N__50063\,
            in2 => \N__47656\,
            in3 => \N__50836\,
            lcout => \c0.n21047\,
            ltout => \c0.n21047_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_330_LC_21_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__64449\,
            in1 => \N__47646\,
            in2 => \N__47632\,
            in3 => \N__54462\,
            lcout => \c0.n42_adj_3111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_2_lut_3_lut_LC_21_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__50485\,
            in1 => \N__47620\,
            in2 => \_gnd_net_\,
            in3 => \N__47555\,
            lcout => \c0.n40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_239_LC_21_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__66326\,
            in1 => \N__54155\,
            in2 => \N__53658\,
            in3 => \N__57091\,
            lcout => OPEN,
            ltout => \c0.n10_adj_3014_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_240_LC_21_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49558\,
            in2 => \N__47512\,
            in3 => \N__56957\,
            lcout => \c0.n19456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i127_LC_21_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__64411\,
            in1 => \N__64247\,
            in2 => \N__47886\,
            in3 => \N__68927\,
            lcout => \c0.data_in_frame_15_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_4_lut_LC_21_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47490\,
            in1 => \N__50191\,
            in2 => \N__50081\,
            in3 => \N__50797\,
            lcout => \c0.n16_adj_3218\,
            ltout => \c0.n16_adj_3218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_873_LC_21_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__51540\,
            in1 => \_gnd_net_\,
            in2 => \N__47479\,
            in3 => \N__58432\,
            lcout => \c0.n12_adj_3469\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i71_LC_21_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__64246\,
            in1 => \N__55876\,
            in2 => \N__68973\,
            in3 => \N__49559\,
            lcout => \c0.data_in_frame_8_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_LC_21_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63232\,
            in2 => \_gnd_net_\,
            in3 => \N__57372\,
            lcout => \c0.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i69_LC_21_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__64245\,
            in1 => \N__55875\,
            in2 => \N__56971\,
            in3 => \N__72659\,
            lcout => \c0.data_in_frame_8_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i72_LC_21_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__64243\,
            in1 => \N__55873\,
            in2 => \N__54162\,
            in3 => \N__72255\,
            lcout => \c0.data_in_frame_8_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71161\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i99_LC_21_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__68594\,
            in1 => \N__67118\,
            in2 => \N__47767\,
            in3 => \N__66155\,
            lcout => \c0.data_in_frame_12_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71161\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i70_LC_21_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__64242\,
            in1 => \N__67854\,
            in2 => \N__57114\,
            in3 => \N__55874\,
            lcout => \c0.data_in_frame_8_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71161\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_874_LC_21_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65515\,
            in2 => \_gnd_net_\,
            in3 => \N__59085\,
            lcout => \c0.n5_adj_3549\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_804_LC_21_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57107\,
            in1 => \N__57024\,
            in2 => \N__56731\,
            in3 => \N__47722\,
            lcout => \c0.n30_adj_3531\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i68_LC_21_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__55872\,
            in1 => \N__64244\,
            in2 => \N__58467\,
            in3 => \N__69409\,
            lcout => \c0.data_in_frame_8_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71161\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_2_lut_adj_563_LC_21_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51436\,
            in2 => \_gnd_net_\,
            in3 => \N__47688\,
            lcout => \c0.n42_adj_3367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_3_lut_adj_806_LC_21_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__54021\,
            in1 => \N__49699\,
            in2 => \_gnd_net_\,
            in3 => \N__49858\,
            lcout => \c0.n31_adj_3532\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_adj_487_LC_21_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62257\,
            in1 => \N__47926\,
            in2 => \N__62313\,
            in3 => \N__56652\,
            lcout => \c0.n9_adj_3350\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_281_LC_21_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48334\,
            in2 => \_gnd_net_\,
            in3 => \N__55952\,
            lcout => \c0.n11942\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_668_LC_21_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47885\,
            in1 => \N__56726\,
            in2 => \N__56533\,
            in3 => \N__65292\,
            lcout => OPEN,
            ltout => \c0.n16_adj_3481_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_670_LC_21_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51139\,
            in1 => \N__47850\,
            in2 => \N__47857\,
            in3 => \N__63109\,
            lcout => \c0.n11815\,
            ltout => \c0.n11815_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_673_LC_21_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58353\,
            in1 => \N__66244\,
            in2 => \N__47854\,
            in3 => \N__58131\,
            lcout => \c0.n10_adj_3483\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_LC_21_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51043\,
            in1 => \N__51033\,
            in2 => \N__63700\,
            in3 => \N__47851\,
            lcout => \c0.n11632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_2_lut_3_lut_adj_720_LC_21_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__62992\,
            in1 => \_gnd_net_\,
            in2 => \N__47836\,
            in3 => \N__47779\,
            lcout => \c0.n35_adj_3266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_933_LC_21_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56668\,
            in1 => \N__56484\,
            in2 => \N__63013\,
            in3 => \N__65434\,
            lcout => \c0.n12056\,
            ltout => \c0.n12056_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_LC_21_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__58931\,
            in1 => \N__59133\,
            in2 => \N__47782\,
            in3 => \N__56528\,
            lcout => \c0.n12_adj_3249\,
            ltout => \c0.n12_adj_3249_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_adj_681_LC_21_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__68383\,
            in1 => \_gnd_net_\,
            in2 => \N__48043\,
            in3 => \N__52351\,
            lcout => \c0.n36_adj_3452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_667_LC_21_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51208\,
            in1 => \N__48040\,
            in2 => \N__69475\,
            in3 => \N__65325\,
            lcout => \c0.n19524\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_285_LC_21_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51214\,
            in1 => \N__58130\,
            in2 => \N__62314\,
            in3 => \N__57267\,
            lcout => \c0.n19301\,
            ltout => \c0.n19301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_828_LC_21_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__48007\,
            in3 => \N__56566\,
            lcout => \c0.n9_adj_3240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_2_lut_3_lut_4_lut_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48130\,
            in1 => \N__47975\,
            in2 => \N__48000\,
            in3 => \N__48930\,
            lcout => \c0.n31_adj_3126\,
            ltout => \c0.n31_adj_3126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_2_lut_4_lut_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63678\,
            in1 => \N__52184\,
            in2 => \N__48004\,
            in3 => \N__52158\,
            lcout => \c0.n35_adj_3317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_2_lut_3_lut_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__52185\,
            in1 => \_gnd_net_\,
            in2 => \N__48001\,
            in3 => \N__47976\,
            lcout => \c0.n46\,
            ltout => \c0.n46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i32_3_lut_4_lut_LC_21_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63679\,
            in1 => \N__47956\,
            in2 => \N__47944\,
            in3 => \N__52159\,
            lcout => \c0.n69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_2_lut_3_lut_LC_21_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__48131\,
            in1 => \N__48721\,
            in2 => \_gnd_net_\,
            in3 => \N__48931\,
            lcout => \c0.n62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_4_lut_adj_451_LC_21_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48722\,
            in1 => \N__48139\,
            in2 => \N__64018\,
            in3 => \N__48132\,
            lcout => \c0.n51_adj_3290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_2_lut_3_lut_LC_21_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__64056\,
            in1 => \N__57502\,
            in2 => \_gnd_net_\,
            in3 => \N__58998\,
            lcout => \c0.n6_adj_3137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_937_LC_21_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__71793\,
            in1 => \N__55867\,
            in2 => \_gnd_net_\,
            in3 => \N__59478\,
            lcout => n19130,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i33_2_lut_3_lut_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__52879\,
            in1 => \_gnd_net_\,
            in2 => \N__58550\,
            in3 => \N__59046\,
            lcout => \c0.n84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_605_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57969\,
            in1 => \N__58954\,
            in2 => \N__52399\,
            in3 => \N__52362\,
            lcout => \c0.n19824\,
            ltout => \c0.n19824_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_501_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__48085\,
            in3 => \N__69986\,
            lcout => OPEN,
            ltout => \c0.n18_adj_3360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_503_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51637\,
            in1 => \N__48081\,
            in2 => \N__48052\,
            in3 => \N__52019\,
            lcout => OPEN,
            ltout => \c0.n32_adj_3362_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_506_LC_21_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51972\,
            in1 => \N__52261\,
            in2 => \N__48049\,
            in3 => \N__48960\,
            lcout => \c0.n20112\,
            ltout => \c0.n20112_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_517_LC_21_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65626\,
            in1 => \N__52134\,
            in2 => \N__48046\,
            in3 => \N__48932\,
            lcout => \c0.n51_adj_3376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_484_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__64623\,
            in1 => \N__48333\,
            in2 => \N__64708\,
            in3 => \N__55960\,
            lcout => \c0.n18398\,
            ltout => \c0.n18398_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_adj_622_LC_21_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__64984\,
            in1 => \_gnd_net_\,
            in2 => \N__48304\,
            in3 => \N__64951\,
            lcout => \c0.n37_adj_3390\,
            ltout => \c0.n37_adj_3390_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_3_lut_LC_21_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__65722\,
            in1 => \_gnd_net_\,
            in2 => \N__48301\,
            in3 => \N__49143\,
            lcout => \c0.n25_adj_3431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i27_4_lut_adj_507_LC_21_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48193\,
            in1 => \N__48163\,
            in2 => \N__51457\,
            in3 => \N__48232\,
            lcout => OPEN,
            ltout => \c0.n60_adj_3368_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i30_4_lut_adj_522_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48298\,
            in1 => \N__48226\,
            in2 => \N__48292\,
            in3 => \N__48289\,
            lcout => \c0.n63_adj_3391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_LC_21_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__48283\,
            in1 => \N__64624\,
            in2 => \_gnd_net_\,
            in3 => \N__48265\,
            lcout => \c0.n39_adj_3334\,
            ltout => \c0.n39_adj_3334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_568_LC_21_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48145\,
            in1 => \N__48225\,
            in2 => \N__48202\,
            in3 => \N__48199\,
            lcout => \c0.n17900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_565_LC_21_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48192\,
            in1 => \N__48181\,
            in2 => \N__51456\,
            in3 => \N__48162\,
            lcout => \c0.n30_adj_3429\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_894_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__53751\,
            in1 => \N__58895\,
            in2 => \_gnd_net_\,
            in3 => \N__53494\,
            lcout => \c0.n35_adj_3274\,
            ltout => \c0.n35_adj_3274_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i26_4_lut_adj_739_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58247\,
            in1 => \N__58217\,
            in2 => \N__48547\,
            in3 => \N__58199\,
            lcout => \c0.n59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__68227\,
            in1 => \N__68120\,
            in2 => \_gnd_net_\,
            in3 => \N__48527\,
            lcout => \c0.n11601\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_825_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__57196\,
            in1 => \N__48511\,
            in2 => \N__55978\,
            in3 => \N__48490\,
            lcout => \c0.n12052\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i40_4_lut_adj_438_LC_21_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57987\,
            in1 => \N__58248\,
            in2 => \N__48451\,
            in3 => \N__48666\,
            lcout => \c0.n91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_adj_628_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__58832\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57747\,
            lcout => \c0.n38_adj_3270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i40_4_lut_adj_521_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57988\,
            in1 => \N__48450\,
            in2 => \N__68047\,
            in3 => \N__48667\,
            lcout => \c0.n91_adj_3389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_2_lut_4_lut_LC_21_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48724\,
            in1 => \N__58649\,
            in2 => \N__69715\,
            in3 => \N__68022\,
            lcout => \c0.n49_adj_3316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_598_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__48436\,
            in1 => \N__48412\,
            in2 => \N__57732\,
            in3 => \N__48391\,
            lcout => \c0.n24_adj_3427\,
            ltout => \c0.n24_adj_3427_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_2_lut_3_lut_LC_21_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64899\,
            in2 => \N__48385\,
            in3 => \N__48382\,
            lcout => \c0.n32_adj_3057\,
            ltout => \c0.n32_adj_3057_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_2_lut_LC_21_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__48727\,
            in3 => \N__48723\,
            lcout => \c0.n44_adj_3125\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_896_LC_21_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__68169\,
            in1 => \N__48697\,
            in2 => \N__48688\,
            in3 => \N__49401\,
            lcout => \c0.n55_adj_3273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_748_LC_21_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__52338\,
            in1 => \N__68430\,
            in2 => \_gnd_net_\,
            in3 => \N__48658\,
            lcout => \c0.n20965\,
            ltout => \c0.n20965_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_767_LC_21_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__48634\,
            in3 => \N__65781\,
            lcout => \c0.n19312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_4_lut_adj_478_LC_21_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48631\,
            in1 => \N__51786\,
            in2 => \N__63457\,
            in3 => \N__49087\,
            lcout => \c0.n20336\,
            ltout => \c0.n20336_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_456_LC_21_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__48618\,
            in1 => \N__53587\,
            in2 => \N__48574\,
            in3 => \N__52446\,
            lcout => \c0.n30_adj_3295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i32_4_lut_adj_523_LC_21_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48571\,
            in1 => \N__49111\,
            in2 => \N__63456\,
            in3 => \N__48559\,
            lcout => \c0.n21034\,
            ltout => \c0.n21034_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_493_LC_21_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52482\,
            in2 => \N__48550\,
            in3 => \N__52505\,
            lcout => \c0.n18377\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_4_lut_adj_520_LC_21_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49147\,
            in1 => \N__53874\,
            in2 => \N__70165\,
            in3 => \N__51785\,
            lcout => \c0.n58_adj_3381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_3_lut_LC_21_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__48876\,
            in1 => \N__58491\,
            in2 => \_gnd_net_\,
            in3 => \N__49105\,
            lcout => \c0.n50_adj_3331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_2_lut_adj_440_LC_21_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48907\,
            in2 => \_gnd_net_\,
            in3 => \N__49080\,
            lcout => \c0.n33_adj_3097\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_406_LC_21_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64949\,
            in1 => \N__58912\,
            in2 => \N__49006\,
            in3 => \N__48991\,
            lcout => OPEN,
            ltout => \c0.n27_adj_3241_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_409_LC_21_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48979\,
            in1 => \N__48964\,
            in2 => \N__48943\,
            in3 => \N__48940\,
            lcout => \c0.n19_adj_3135\,
            ltout => \c0.n19_adj_3135_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_2_lut_adj_347_LC_21_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__48901\,
            in3 => \N__48898\,
            lcout => OPEN,
            ltout => \c0.n22_adj_3136_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_348_LC_21_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63455\,
            in1 => \N__48880\,
            in2 => \N__48844\,
            in3 => \N__51787\,
            lcout => \c0.n11936\,
            ltout => \c0.n11936_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_700_LC_21_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49260\,
            in1 => \N__49227\,
            in2 => \N__48841\,
            in3 => \N__48837\,
            lcout => \c0.n20_adj_3293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_472_LC_21_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__49536\,
            in1 => \N__48790\,
            in2 => \N__49182\,
            in3 => \N__52447\,
            lcout => \c0.n17_adj_3318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_774_LC_21_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49261\,
            in1 => \N__49228\,
            in2 => \N__59701\,
            in3 => \N__49535\,
            lcout => \c0.n12_adj_3141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_326_LC_21_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49506\,
            in2 => \_gnd_net_\,
            in3 => \N__49454\,
            lcout => OPEN,
            ltout => \c0.n19465_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_331_LC_21_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68157\,
            in1 => \N__53280\,
            in2 => \N__49414\,
            in3 => \N__53837\,
            lcout => \c0.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_379_LC_21_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__53838\,
            in1 => \N__68158\,
            in2 => \N__53284\,
            in3 => \N__49402\,
            lcout => \c0.n19703\,
            ltout => \c0.n19703_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_443_LC_21_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49160\,
            in1 => \N__58715\,
            in2 => \N__49357\,
            in3 => \N__59588\,
            lcout => \c0.n44_adj_3278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_319_LC_21_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49328\,
            in2 => \_gnd_net_\,
            in3 => \N__49257\,
            lcout => \c0.n7_adj_3094\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_3_lut_adj_756_LC_21_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__69988\,
            in1 => \N__72859\,
            in2 => \_gnd_net_\,
            in3 => \N__49288\,
            lcout => \c0.n33_adj_3279\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_381_LC_21_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49258\,
            in2 => \_gnd_net_\,
            in3 => \N__49229\,
            lcout => \c0.n19400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_LC_21_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__53768\,
            in1 => \N__70044\,
            in2 => \_gnd_net_\,
            in3 => \N__66395\,
            lcout => \c0.n36_adj_3275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_291_LC_21_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__49789\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53255\,
            lcout => \c0.n17840\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i185_LC_21_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53769\,
            in1 => \N__65247\,
            in2 => \_gnd_net_\,
            in3 => \N__53721\,
            lcout => data_in_frame_23_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__0__5173_LC_21_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__65246\,
            in1 => \N__53230\,
            in2 => \_gnd_net_\,
            in3 => \N__49730\,
            lcout => data_in_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i192_LC_21_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__72293\,
            in1 => \N__53722\,
            in2 => \_gnd_net_\,
            in3 => \N__66396\,
            lcout => data_in_frame_23_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_769_LC_22_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54842\,
            in2 => \_gnd_net_\,
            in3 => \N__54673\,
            lcout => \c0.n12_adj_3498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_5_i6_2_lut_LC_22_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49676\,
            in2 => \_gnd_net_\,
            in3 => \N__60729\,
            lcout => \c0.n6_adj_3149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_911_LC_22_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54199\,
            in1 => \N__57005\,
            in2 => \N__49581\,
            in3 => \N__56399\,
            lcout => \c0.n13_adj_3344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_adj_907_LC_22_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__49577\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57006\,
            lcout => \c0.n35_adj_3233\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_837_LC_22_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62625\,
            in1 => \N__61198\,
            in2 => \N__49984\,
            in3 => \N__60908\,
            lcout => \c0.n17_adj_3113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_2_lut_3_lut_adj_901_LC_22_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__54675\,
            in1 => \N__54308\,
            in2 => \_gnd_net_\,
            in3 => \N__54770\,
            lcout => \c0.n60\,
            ltout => \c0.n60_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i41_4_lut_LC_22_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57004\,
            in1 => \N__49939\,
            in2 => \N__49933\,
            in3 => \N__54901\,
            lcout => \c0.n93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i16_LC_22_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__72200\,
            in1 => \_gnd_net_\,
            in2 => \N__54684\,
            in3 => \N__59883\,
            lcout => data_in_frame_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_763_LC_22_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49916\,
            in2 => \_gnd_net_\,
            in3 => \N__54851\,
            lcout => \c0.n5_adj_3028\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i52_LC_22_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62009\,
            in1 => \N__61598\,
            in2 => \N__54022\,
            in3 => \N__69443\,
            lcout => \c0.data_in_frame_6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_770_LC_22_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__54771\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54676\,
            lcout => \c0.n7_adj_3520\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_760_LC_22_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__55584\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55349\,
            lcout => \c0.n19443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_764_LC_22_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__61347\,
            in1 => \_gnd_net_\,
            in2 => \N__49809\,
            in3 => \N__55544\,
            lcout => \c0.n11687\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_adj_848_LC_22_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62354\,
            in1 => \N__49802\,
            in2 => \N__55548\,
            in3 => \N__61346\,
            lcout => OPEN,
            ltout => \c0.n8_adj_3066_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_292_LC_22_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51478\,
            in1 => \N__55725\,
            in2 => \N__50185\,
            in3 => \N__60906\,
            lcout => \c0.n19170\,
            ltout => \c0.n19170_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_839_LC_22_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62399\,
            in2 => \N__50161\,
            in3 => \N__50150\,
            lcout => \c0.n21_adj_3053\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_843_LC_22_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54836\,
            in1 => \N__55015\,
            in2 => \N__55162\,
            in3 => \N__60905\,
            lcout => \c0.n15_adj_3545\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_adj_612_LC_22_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__55016\,
            in1 => \N__61254\,
            in2 => \_gnd_net_\,
            in3 => \N__50313\,
            lcout => \c0.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i10_LC_22_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__54126\,
            in1 => \N__59876\,
            in2 => \_gnd_net_\,
            in3 => \N__71419\,
            lcout => data_in_frame_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i12_LC_22_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__59875\,
            in1 => \N__69425\,
            in2 => \_gnd_net_\,
            in3 => \N__61212\,
            lcout => data_in_frame_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_706_LC_22_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50022\,
            in1 => \N__50394\,
            in2 => \N__50432\,
            in3 => \N__50285\,
            lcout => \c0.n20340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i37_3_lut_LC_22_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__55505\,
            in1 => \N__61205\,
            in2 => \_gnd_net_\,
            in3 => \N__50004\,
            lcout => \c0.n89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i28_LC_22_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__61408\,
            in1 => \N__69438\,
            in2 => \N__50433\,
            in3 => \N__61744\,
            lcout => \c0.data_in_frame_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71206\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i27_LC_22_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__50395\,
            in1 => \N__68674\,
            in2 => \N__61777\,
            in3 => \N__61407\,
            lcout => \c0.data_in_frame_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71206\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_adj_615_LC_22_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__50674\,
            in1 => \N__55128\,
            in2 => \_gnd_net_\,
            in3 => \N__50603\,
            lcout => \c0.n33_adj_3088\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i8_LC_22_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__72199\,
            in1 => \N__50361\,
            in2 => \N__61778\,
            in3 => \N__55885\,
            lcout => \data_out_frame_29__3__N_647\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71206\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i7_LC_22_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__55884\,
            in1 => \N__55129\,
            in2 => \N__68854\,
            in3 => \N__61745\,
            lcout => data_in_frame_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71206\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_845_LC_22_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50467\,
            in1 => \N__55724\,
            in2 => \N__50456\,
            in3 => \N__50425\,
            lcout => \c0.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_419_LC_22_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__59485\,
            in1 => \_gnd_net_\,
            in2 => \N__61424\,
            in3 => \_gnd_net_\,
            lcout => \c0.n19131\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_adj_576_LC_22_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__50393\,
            in1 => \N__55109\,
            in2 => \_gnd_net_\,
            in3 => \N__50286\,
            lcout => \c0.n29_adj_3216\,
            ltout => \c0.n29_adj_3216_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_4_lut_LC_22_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50226\,
            in1 => \N__50209\,
            in2 => \N__50194\,
            in3 => \N__50869\,
            lcout => \c0.n44_adj_3217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_382_LC_22_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50853\,
            in1 => \N__50933\,
            in2 => \N__57633\,
            in3 => \N__50977\,
            lcout => OPEN,
            ltout => \c0.n36_adj_3212_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_384_LC_22_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54966\,
            in1 => \N__55696\,
            in2 => \N__50872\,
            in3 => \N__54460\,
            lcout => \c0.n41_adj_3213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_722_LC_22_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__50852\,
            in1 => \N__54965\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n11651\,
            ltout => \c0.n11651_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_3_lut_LC_22_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55697\,
            in2 => \N__50839\,
            in3 => \N__50796\,
            lcout => \c0.n27_adj_3082\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_2_lut_adj_380_LC_22_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__51090\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50822\,
            lcout => \c0.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_4_lut_adj_394_LC_22_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51421\,
            in1 => \N__62889\,
            in2 => \N__50785\,
            in3 => \N__56848\,
            lcout => OPEN,
            ltout => \c0.n52_adj_3223_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i26_4_lut_LC_22_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50749\,
            in1 => \N__50740\,
            in2 => \N__50716\,
            in3 => \N__56365\,
            lcout => \c0.n54_adj_3234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i63_LC_22_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__61766\,
            in1 => \N__64413\,
            in2 => \N__56351\,
            in3 => \N__68825\,
            lcout => \c0.data_in_frame_7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i32_4_lut_adj_732_LC_22_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54937\,
            in1 => \N__56272\,
            in2 => \N__50713\,
            in3 => \N__50698\,
            lcout => \c0.n46_adj_3443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i183_LC_22_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__53794\,
            in1 => \N__67531\,
            in2 => \_gnd_net_\,
            in3 => \N__68824\,
            lcout => data_in_frame_22_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i61_LC_22_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__64412\,
            in1 => \N__61767\,
            in2 => \N__51104\,
            in3 => \N__72660\,
            lcout => \c0.data_in_frame_7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i62_LC_22_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__67948\,
            in1 => \N__61768\,
            in2 => \N__55708\,
            in3 => \N__64414\,
            lcout => \c0.data_in_frame_7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i85_LC_22_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__51539\,
            in1 => \N__62810\,
            in2 => \N__66066\,
            in3 => \N__72738\,
            lcout => \c0.data_in_frame_10_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_2_lut_3_lut_adj_878_LC_22_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__58431\,
            in1 => \N__51538\,
            in2 => \_gnd_net_\,
            in3 => \N__51061\,
            lcout => \c0.n45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_222_LC_22_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65407\,
            in2 => \_gnd_net_\,
            in3 => \N__61285\,
            lcout => \c0.n4\,
            ltout => \c0.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_876_LC_22_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51037\,
            in1 => \N__51016\,
            in2 => \N__50992\,
            in3 => \N__50988\,
            lcout => \c0.n26_adj_3550\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i81_LC_22_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62830\,
            in1 => \N__66184\,
            in2 => \N__50937\,
            in3 => \N__65118\,
            lcout => \c0.data_in_frame_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i109_LC_22_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__72739\,
            in1 => \N__71970\,
            in2 => \N__63048\,
            in3 => \N__66007\,
            lcout => \c0.data_in_frame_13_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i169_LC_22_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__71969\,
            in1 => \N__71800\,
            in2 => \N__50903\,
            in3 => \N__65117\,
            lcout => \c0.data_in_frame_21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_adj_393_LC_22_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51432\,
            in1 => \N__51711\,
            in2 => \N__63799\,
            in3 => \N__58599\,
            lcout => \c0.n48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_880_LC_22_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51415\,
            in1 => \N__51349\,
            in2 => \N__51301\,
            in3 => \N__51292\,
            lcout => \c0.n27_adj_3551\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i86_LC_22_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__56904\,
            in1 => \N__67947\,
            in2 => \N__66204\,
            in3 => \N__62844\,
            lcout => \c0.data_in_frame_10_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_280_LC_22_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__63034\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51706\,
            lcout => \c0.n11613\,
            ltout => \c0.n11613_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_669_LC_22_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51207\,
            in1 => \N__51178\,
            in2 => \N__51157\,
            in3 => \N__51153\,
            lcout => \c0.n17_adj_3482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3106_2_lut_LC_22_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51122\,
            in2 => \_gnd_net_\,
            in3 => \N__56027\,
            lcout => \c0.n5753\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i111_LC_22_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__66177\,
            in1 => \N__68923\,
            in2 => \N__51129\,
            in3 => \N__71948\,
            lcout => \c0.data_in_frame_13_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i166_LC_22_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__67945\,
            in1 => \N__67131\,
            in2 => \N__71806\,
            in3 => \N__72424\,
            lcout => \c0.data_in_frame_20_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i110_LC_22_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__51707\,
            in1 => \N__67946\,
            in2 => \N__66203\,
            in3 => \N__71947\,
            lcout => \c0.data_in_frame_13_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_401_LC_22_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__65406\,
            in1 => \N__51514\,
            in2 => \N__64821\,
            in3 => \N__51688\,
            lcout => OPEN,
            ltout => \c0.n43_adj_3232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i27_4_lut_LC_22_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51553\,
            in1 => \N__51649\,
            in2 => \N__51640\,
            in3 => \N__51601\,
            lcout => \c0.n47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_3_lut_LC_22_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__58404\,
            in1 => \N__51636\,
            in2 => \_gnd_net_\,
            in3 => \N__52015\,
            lcout => \c0.n49_adj_3237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_adj_903_LC_22_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60843\,
            in1 => \N__62497\,
            in2 => \N__55959\,
            in3 => \N__60791\,
            lcout => \c0.n7_adj_3225\,
            ltout => \c0.n7_adj_3225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_666_LC_22_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56560\,
            in1 => \N__51588\,
            in2 => \N__51595\,
            in3 => \N__62307\,
            lcout => \c0.n11590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_395_LC_22_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62308\,
            in1 => \N__64703\,
            in2 => \N__51592\,
            in3 => \N__51559\,
            lcout => \c0.n44_adj_3226\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_750_LC_22_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65680\,
            in2 => \_gnd_net_\,
            in3 => \N__65795\,
            lcout => \c0.n19202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_2_lut_3_lut_adj_872_LC_22_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__51544\,
            in1 => \N__58462\,
            in2 => \_gnd_net_\,
            in3 => \N__51513\,
            lcout => \c0.n41_adj_3365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_3_lut_4_lut_LC_22_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63630\,
            in1 => \N__51730\,
            in2 => \N__63688\,
            in3 => \N__52166\,
            lcout => OPEN,
            ltout => \c0.n47_adj_3286_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_4_lut_adj_450_LC_22_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__67673\,
            in1 => \N__51892\,
            in2 => \N__51874\,
            in3 => \N__58068\,
            lcout => OPEN,
            ltout => \c0.n52_adj_3288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_452_LC_22_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51871\,
            in1 => \N__65452\,
            in2 => \N__51865\,
            in3 => \N__57760\,
            lcout => \c0.n6_adj_3291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i95_LC_22_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__64542\,
            in1 => \N__51833\,
            in2 => \N__66205\,
            in3 => \N__69011\,
            lcout => \c0.data_in_frame_11_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__63574\,
            in1 => \N__63495\,
            in2 => \_gnd_net_\,
            in3 => \N__51775\,
            lcout => \c0.n19909\,
            ltout => \c0.n19909_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i36_3_lut_4_lut_LC_22_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63628\,
            in1 => \N__63683\,
            in2 => \N__51811\,
            in3 => \N__58067\,
            lcout => \c0.n87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_2_lut_3_lut_adj_648_LC_22_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__63629\,
            in1 => \N__63496\,
            in2 => \_gnd_net_\,
            in3 => \N__51776\,
            lcout => \c0.n35_adj_3098\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i28_4_lut_adj_309_LC_22_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__52543\,
            in1 => \N__59010\,
            in2 => \N__57820\,
            in3 => \N__53506\,
            lcout => \c0.n65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_2_lut_3_lut_LC_22_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__63776\,
            in1 => \N__65519\,
            in2 => \_gnd_net_\,
            in3 => \N__51729\,
            lcout => \c0.n45_adj_3423\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_340_LC_22_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65796\,
            in2 => \_gnd_net_\,
            in3 => \N__53943\,
            lcout => \c0.n7_adj_3047\,
            ltout => \c0.n7_adj_3047_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_344_LC_22_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52231\,
            in1 => \N__52216\,
            in2 => \N__52195\,
            in3 => \N__59358\,
            lcout => \c0.n7_adj_3079\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_3_lut_adj_603_LC_22_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__64057\,
            in1 => \N__57501\,
            in2 => \_gnd_net_\,
            in3 => \N__63485\,
            lcout => \c0.n28_adj_3059\,
            ltout => \c0.n28_adj_3059_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_2_lut_3_lut_LC_22_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__63627\,
            in1 => \_gnd_net_\,
            in2 => \N__52192\,
            in3 => \N__63560\,
            lcout => \c0.n33_adj_3315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_2_lut_3_lut_4_lut_LC_22_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63775\,
            in1 => \N__52189\,
            in2 => \N__65526\,
            in3 => \N__52167\,
            lcout => \c0.n32_adj_3465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_3_lut_4_lut_LC_22_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52135\,
            in1 => \N__52108\,
            in2 => \N__55675\,
            in3 => \N__52060\,
            lcout => OPEN,
            ltout => \c0.n29_adj_3461_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_625_LC_22_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52249\,
            in1 => \N__52054\,
            in2 => \N__52024\,
            in3 => \N__52021\,
            lcout => OPEN,
            ltout => \c0.n36_adj_3470_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_626_LC_22_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51973\,
            in1 => \N__51946\,
            in2 => \N__51919\,
            in3 => \N__51916\,
            lcout => \c0.n11_adj_3124\,
            ltout => \c0.n11_adj_3124_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_629_LC_22_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__53804\,
            in1 => \_gnd_net_\,
            in2 => \N__51895\,
            in3 => \_gnd_net_\,
            lcout => \c0.n37_adj_3268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i27_2_lut_LC_22_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52397\,
            in2 => \_gnd_net_\,
            in3 => \N__52405\,
            lcout => \c0.n58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_adj_339_LC_22_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58840\,
            in2 => \_gnd_net_\,
            in3 => \N__57952\,
            lcout => \c0.n42_adj_3086\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i26_4_lut_adj_471_LC_22_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52398\,
            in1 => \N__52378\,
            in2 => \N__57940\,
            in3 => \N__52366\,
            lcout => \c0.n19764\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_890_LC_22_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__69965\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__72832\,
            lcout => \c0.n11971\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_664_LC_22_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__72833\,
            in1 => \N__69966\,
            in2 => \_gnd_net_\,
            in3 => \N__69636\,
            lcout => \c0.n18379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_adj_683_LC_22_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52350\,
            in1 => \N__67404\,
            in2 => \N__68392\,
            in3 => \N__52282\,
            lcout => \c0.n22_adj_3363\,
            ltout => \c0.n22_adj_3363_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_adj_623_LC_22_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__69496\,
            in1 => \_gnd_net_\,
            in2 => \N__52252\,
            in3 => \N__69964\,
            lcout => \c0.n30_adj_3468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_513_LC_22_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__68300\,
            in1 => \N__68428\,
            in2 => \N__68391\,
            in3 => \N__69818\,
            lcout => \c0.n6009\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i33_4_lut_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57883\,
            in1 => \N__52240\,
            in2 => \N__57909\,
            in3 => \N__52416\,
            lcout => OPEN,
            ltout => \c0.n70_adj_3087_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i36_4_lut_LC_22_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57838\,
            in1 => \N__58612\,
            in2 => \N__52693\,
            in3 => \N__57928\,
            lcout => \c0.n20339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_adj_655_LC_22_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__72834\,
            in1 => \N__69967\,
            in2 => \_gnd_net_\,
            in3 => \N__53459\,
            lcout => \c0.n27_adj_3311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_455_LC_22_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52645\,
            in1 => \N__52615\,
            in2 => \N__66694\,
            in3 => \N__52606\,
            lcout => OPEN,
            ltout => \c0.n32_adj_3294_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_459_LC_22_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53443\,
            in1 => \N__52588\,
            in2 => \N__52582\,
            in3 => \N__52525\,
            lcout => \c0.n21075\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_4_lut_LC_22_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__52708\,
            in1 => \N__52559\,
            in2 => \N__52489\,
            in3 => \N__57857\,
            lcout => \c0.n29_adj_3299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i172_LC_22_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__71778\,
            in1 => \N__71977\,
            in2 => \N__69602\,
            in3 => \N__69287\,
            lcout => \c0.data_in_frame_21_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_473_LC_22_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__52507\,
            in1 => \N__52707\,
            in2 => \N__52490\,
            in3 => \N__57858\,
            lcout => \c0.n19_adj_3320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_3_lut_4_lut_adj_783_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52706\,
            in1 => \N__52506\,
            in2 => \N__52492\,
            in3 => \N__52445\,
            lcout => \c0.n57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_adj_584_LC_22_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52875\,
            in2 => \_gnd_net_\,
            in3 => \N__59032\,
            lcout => \c0.n39_adj_3384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_adj_695_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53342\,
            in1 => \N__53391\,
            in2 => \N__68125\,
            in3 => \N__53298\,
            lcout => \c0.n11714\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_457_LC_22_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52735\,
            in1 => \N__68124\,
            in2 => \N__53395\,
            in3 => \N__53343\,
            lcout => \c0.n22_adj_3296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_321_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68236\,
            in2 => \_gnd_net_\,
            in3 => \N__53297\,
            lcout => \c0.n19159\,
            ltout => \c0.n19159_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_749_LC_22_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53808\,
            in1 => \N__72438\,
            in2 => \N__52831\,
            in3 => \N__52828\,
            lcout => \c0.n12206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i30_4_lut_adj_504_LC_22_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52804\,
            in1 => \N__53353\,
            in2 => \N__52798\,
            in3 => \N__53585\,
            lcout => \c0.n79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_373_LC_22_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__58041\,
            in1 => \N__58794\,
            in2 => \_gnd_net_\,
            in3 => \N__53421\,
            lcout => \c0.n19151\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_364_LC_22_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__52762\,
            in1 => \N__59011\,
            in2 => \N__57256\,
            in3 => \N__52734\,
            lcout => \c0.n11776\,
            ltout => \c0.n11776_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_561_LC_22_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__68235\,
            in1 => \N__72437\,
            in2 => \N__52711\,
            in3 => \N__59504\,
            lcout => \c0.n6_adj_3319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_317_LC_22_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__53626\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53601\,
            lcout => \c0.n19268\,
            ltout => \c0.n19268_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_4_lut_adj_649_LC_22_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53511\,
            in1 => \N__66647\,
            in2 => \N__53563\,
            in3 => \N__53539\,
            lcout => \c0.n20_adj_3301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_LC_22_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53538\,
            in1 => \N__53510\,
            in2 => \N__66649\,
            in3 => \N__53469\,
            lcout => \c0.n42_adj_3055\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_323_LC_22_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__67697\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53425\,
            lcout => \c0.n4_adj_3100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_375_LC_22_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__53272\,
            in1 => \N__53375\,
            in2 => \N__58114\,
            in3 => \N__64632\,
            lcout => \c0.n19436\,
            ltout => \c0.n19436_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_adj_697_LC_22_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53344\,
            in1 => \N__68119\,
            in2 => \N__53302\,
            in3 => \N__53299\,
            lcout => \c0.n6_adj_3112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_336_LC_22_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53271\,
            in1 => \N__69787\,
            in2 => \N__58849\,
            in3 => \N__67696\,
            lcout => \c0.n20933\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__6__5175_LC_22_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53135\,
            in1 => \N__52960\,
            in2 => \_gnd_net_\,
            in3 => \N__52903\,
            lcout => data_in_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71207\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_LC_22_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__59274\,
            in1 => \N__59230\,
            in2 => \_gnd_net_\,
            in3 => \N__59828\,
            lcout => \c0.n25_adj_3048\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_377_LC_22_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72392\,
            in1 => \N__53973\,
            in2 => \N__69606\,
            in3 => \N__53947\,
            lcout => OPEN,
            ltout => \c0.n12_adj_3210_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_378_LC_22_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__53911\,
            in1 => \N__66453\,
            in2 => \N__53884\,
            in3 => \N__53881\,
            lcout => \c0.n17834\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_rep_109_2_lut_LC_22_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__59231\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59275\,
            lcout => \c0.n21767\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_338_LC_22_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__53809\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53770\,
            lcout => \c0.n41_adj_3085\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i189_LC_22_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__72733\,
            in1 => \N__53709\,
            in2 => \_gnd_net_\,
            in3 => \N__53744\,
            lcout => data_in_frame_23_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i190_LC_22_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53710\,
            in1 => \N__67980\,
            in2 => \_gnd_net_\,
            in3 => \N__66454\,
            lcout => data_in_frame_23_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_67_i9_2_lut_3_lut_LC_23_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__60268\,
            in1 => \N__59996\,
            in2 => \_gnd_net_\,
            in3 => \N__60117\,
            lcout => \c0.n9_adj_3211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_LC_23_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54211\,
            in1 => \N__54187\,
            in2 => \N__53662\,
            in3 => \N__54579\,
            lcout => \c0.n7_adj_3347\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_812_LC_23_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__54680\,
            in1 => \N__55377\,
            in2 => \N__54628\,
            in3 => \N__60922\,
            lcout => \c0.n34_adj_3326\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_adj_912_LC_23_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__54186\,
            in1 => \_gnd_net_\,
            in2 => \N__54580\,
            in3 => \N__54210\,
            lcout => \c0.n11982\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_4_lut_adj_719_LC_23_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54568\,
            in1 => \N__54530\,
            in2 => \N__54502\,
            in3 => \N__54480\,
            lcout => \c0.n58_adj_3497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_771_LC_23_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54315\,
            in2 => \_gnd_net_\,
            in3 => \N__54271\,
            lcout => \c0.n8_adj_3345\,
            ltout => \c0.n8_adj_3345_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_779_LC_23_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54198\,
            in1 => \N__54185\,
            in2 => \N__54172\,
            in3 => \N__56398\,
            lcout => \c0.n11626\,
            ltout => \c0.n11626_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_372_LC_23_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__54169\,
            in3 => \N__54166\,
            lcout => \c0.n12209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_519_LC_23_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54634\,
            in1 => \N__54115\,
            in2 => \N__54858\,
            in3 => \N__55277\,
            lcout => \c0.n19970\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_728_LC_23_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54031\,
            in1 => \N__54834\,
            in2 => \N__54020\,
            in3 => \N__54672\,
            lcout => \c0.n11478\,
            ltout => \c0.n11478_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i29_4_lut_LC_23_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56630\,
            in1 => \N__54781\,
            in2 => \N__54904\,
            in3 => \N__54731\,
            lcout => \c0.n81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i15_LC_23_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__68866\,
            in1 => \N__59884\,
            in2 => \_gnd_net_\,
            in3 => \N__54835\,
            lcout => data_in_frame_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_835_LC_23_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60907\,
            in2 => \_gnd_net_\,
            in3 => \N__62624\,
            lcout => \c0.n11526\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i54_LC_23_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62030\,
            in1 => \N__61615\,
            in2 => \N__54775\,
            in3 => \N__67912\,
            lcout => \c0.data_in_frame_6_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_606_LC_23_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__56938\,
            in1 => \N__57043\,
            in2 => \N__54757\,
            in3 => \N__54732\,
            lcout => \c0.n27_adj_3457\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_805_LC_23_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61193\,
            in2 => \_gnd_net_\,
            in3 => \N__54671\,
            lcout => \c0.n12_adj_3378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i48_LC_23_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__61757\,
            in1 => \N__60352\,
            in2 => \N__62681\,
            in3 => \N__72149\,
            lcout => \c0.data_in_frame_5_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i13_LC_23_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__59866\,
            in1 => \N__72613\,
            in2 => \_gnd_net_\,
            in3 => \N__60916\,
            lcout => data_in_frame_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i14_LC_23_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__67911\,
            in1 => \N__59867\,
            in2 => \_gnd_net_\,
            in3 => \N__55345\,
            lcout => data_in_frame_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_adj_564_LC_23_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__55420\,
            in1 => \N__55411\,
            in2 => \_gnd_net_\,
            in3 => \N__60842\,
            lcout => \c0.n28_adj_3428\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_800_LC_23_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60388\,
            in1 => \N__60899\,
            in2 => \_gnd_net_\,
            in3 => \N__55344\,
            lcout => \c0.n7_adj_3509\,
            ltout => \c0.n7_adj_3509_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_803_LC_23_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__55294\,
            in3 => \N__55010\,
            lcout => \c0.n10_adj_3012\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i9_LC_23_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65259\,
            in2 => \N__55031\,
            in3 => \N__59868\,
            lcout => data_in_frame_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_3_lut_4_lut_adj_862_LC_23_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62409\,
            in1 => \N__55264\,
            in2 => \N__62464\,
            in3 => \N__55240\,
            lcout => \c0.n56_adj_3505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_709_LC_23_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__55108\,
            in1 => \N__55014\,
            in2 => \_gnd_net_\,
            in3 => \N__60389\,
            lcout => \c0.n20341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i31_4_lut_adj_731_LC_23_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54910\,
            in1 => \N__54952\,
            in2 => \N__61141\,
            in3 => \N__54943\,
            lcout => \c0.n64_adj_3506\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_838_LC_23_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61326\,
            in2 => \_gnd_net_\,
            in3 => \N__60390\,
            lcout => \c0.n4_adj_3036\,
            ltout => \c0.n4_adj_3036_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_4_lut_adj_723_LC_23_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62353\,
            in1 => \N__54925\,
            in2 => \N__54913\,
            in3 => \N__62619\,
            lcout => \c0.n57_adj_3499\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_899_LC_23_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__62618\,
            in1 => \N__61327\,
            in2 => \_gnd_net_\,
            in3 => \N__60391\,
            lcout => \c0.n6_adj_3019\,
            ltout => \c0.n6_adj_3019_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_244_LC_23_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62320\,
            in1 => \N__55704\,
            in2 => \N__55678\,
            in3 => \N__60909\,
            lcout => \c0.n20386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i79_LC_23_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66145\,
            in1 => \N__63418\,
            in2 => \N__55614\,
            in3 => \N__68826\,
            lcout => \c0.data_in_frame_9_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71220\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i64_LC_23_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__64409\,
            in1 => \N__61756\,
            in2 => \N__62410\,
            in3 => \N__72132\,
            lcout => \c0.data_in_frame_7_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i32_LC_23_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__61752\,
            in1 => \N__61455\,
            in2 => \N__72201\,
            in3 => \N__55583\,
            lcout => \c0.data_in_frame_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i30_LC_23_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__61454\,
            in1 => \N__61754\,
            in2 => \N__62626\,
            in3 => \N__67952\,
            lcout => \c0.data_in_frame_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i46_LC_23_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__61753\,
            in1 => \N__67951\,
            in2 => \N__60358\,
            in3 => \N__55540\,
            lcout => \c0.data_in_frame_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i44_LC_23_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__69442\,
            in1 => \N__61755\,
            in2 => \N__55515\,
            in3 => \N__60354\,
            lcout => \c0.data_in_frame_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i7_LC_23_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__72128\,
            in1 => \N__56266\,
            in2 => \N__56226\,
            in3 => \N__55468\,
            lcout => rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_3_lut_4_lut_LC_23_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60487\,
            in1 => \N__60448\,
            in2 => \N__62496\,
            in3 => \N__56295\,
            lcout => \c0.n51_adj_3426\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i6_LC_23_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__56259\,
            in1 => \N__68853\,
            in2 => \N__56225\,
            in3 => \N__56085\,
            lcout => rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_823_LC_23_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64438\,
            in1 => \N__56028\,
            in2 => \N__57500\,
            in3 => \N__61873\,
            lcout => \c0.n13_adj_3541\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i102_LC_23_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__67949\,
            in1 => \N__67220\,
            in2 => \N__66189\,
            in3 => \N__57632\,
            lcout => \c0.data_in_frame_12_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71196\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i107_LC_23_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__68725\,
            in1 => \N__71972\,
            in2 => \N__55951\,
            in3 => \N__66162\,
            lcout => \c0.data_in_frame_13_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71196\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i78_LC_23_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__67950\,
            in1 => \N__66193\,
            in2 => \N__55920\,
            in3 => \N__63380\,
            lcout => \c0.data_in_frame_9_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71196\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i65_LC_23_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__65230\,
            in1 => \N__62447\,
            in2 => \N__64249\,
            in3 => \N__55812\,
            lcout => \c0.data_in_frame_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71196\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i97_LC_23_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66157\,
            in1 => \N__67221\,
            in2 => \N__57195\,
            in3 => \N__65234\,
            lcout => \c0.data_in_frame_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71196\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i73_LC_23_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__63379\,
            in1 => \N__66158\,
            in2 => \N__65258\,
            in3 => \N__63104\,
            lcout => \c0.data_in_frame_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71196\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_LC_23_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__62250\,
            in1 => \N__56410\,
            in2 => \_gnd_net_\,
            in3 => \N__56847\,
            lcout => \c0.n17_adj_3544\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_359_LC_23_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__56939\,
            in1 => \N__57103\,
            in2 => \_gnd_net_\,
            in3 => \N__57044\,
            lcout => OPEN,
            ltout => \c0.n11858_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_371_LC_23_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56727\,
            in2 => \N__56671\,
            in3 => \N__61871\,
            lcout => \c0.n19446\,
            ltout => \c0.n19446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_376_LC_23_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62904\,
            in2 => \N__56656\,
            in3 => \N__56653\,
            lcout => \c0.n33_adj_3209\,
            ltout => \c0.n33_adj_3209_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_adj_827_LC_23_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56578\,
            in2 => \N__56569\,
            in3 => \N__56440\,
            lcout => \c0.n5598\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_809_LC_23_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61872\,
            in1 => \N__56529\,
            in2 => \N__65433\,
            in3 => \N__56488\,
            lcout => \c0.n29_adj_3533\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_3_lut_LC_23_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__56458\,
            in1 => \N__56441\,
            in2 => \_gnd_net_\,
            in3 => \N__56409\,
            lcout => \c0.n45_adj_3224\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_LC_23_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56341\,
            in2 => \_gnd_net_\,
            in3 => \N__62679\,
            lcout => \c0.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_391_LC_23_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57401\,
            in1 => \N__57271\,
            in2 => \N__57251\,
            in3 => \N__57187\,
            lcout => \c0.n19430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_adj_917_LC_23_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62720\,
            in2 => \_gnd_net_\,
            in3 => \N__57157\,
            lcout => \c0.n20_adj_3536\,
            ltout => \c0.n20_adj_3536_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_918_LC_23_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56917\,
            in2 => \N__57121\,
            in3 => \N__58598\,
            lcout => OPEN,
            ltout => \c0.n12_adj_3558_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_919_LC_23_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__66354\,
            in1 => \N__60745\,
            in2 => \N__57118\,
            in3 => \N__58461\,
            lcout => \c0.n18420\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_906_LC_23_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57115\,
            in1 => \N__56940\,
            in2 => \N__57076\,
            in3 => \N__57046\,
            lcout => \c0.n19359\,
            ltout => \c0.n19359_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_392_LC_23_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__56974\,
            in3 => \N__56902\,
            lcout => \c0.n19502\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_914_LC_23_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56970\,
            in2 => \_gnd_net_\,
            in3 => \N__56941\,
            lcout => \c0.n19199\,
            ltout => \c0.n19199_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_820_LC_23_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59530\,
            in1 => \N__56903\,
            in2 => \N__56881\,
            in3 => \N__66294\,
            lcout => \c0.n19_adj_3540\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i142_LC_23_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__63416\,
            in1 => \N__67981\,
            in2 => \N__65326\,
            in3 => \N__71802\,
            lcout => \c0.data_in_frame_17_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i122_LC_23_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__71488\,
            in1 => \N__64254\,
            in2 => \N__64389\,
            in3 => \N__64979\,
            lcout => \c0.data_in_frame_15_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i208_LC_23_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__63417\,
            in1 => \N__66898\,
            in2 => \N__59783\,
            in3 => \N__72206\,
            lcout => \c0.data_in_frame_25_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i114_LC_23_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__71487\,
            in1 => \N__64252\,
            in2 => \N__57499\,
            in3 => \N__62058\,
            lcout => \c0.data_in_frame_14_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i128_LC_23_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__64251\,
            in1 => \N__64362\,
            in2 => \N__57434\,
            in3 => \N__72205\,
            lcout => \c0.data_in_frame_15_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i115_LC_23_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__68722\,
            in1 => \N__64253\,
            in2 => \N__57408\,
            in3 => \N__62059\,
            lcout => \c0.data_in_frame_14_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i59_LC_23_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__57361\,
            in1 => \N__68723\,
            in2 => \N__61599\,
            in3 => \N__64366\,
            lcout => \c0.data_in_frame_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_360_LC_23_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__62527\,
            in1 => \N__62680\,
            in2 => \N__62551\,
            in3 => \N__57331\,
            lcout => \c0.n25_adj_3157\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_4_lut_adj_865_LC_23_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69688\,
            in1 => \N__70083\,
            in2 => \N__58899\,
            in3 => \N__59009\,
            lcout => \c0.n32_adj_3060\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_290_LC_23_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59047\,
            in1 => \N__58667\,
            in2 => \N__70498\,
            in3 => \N__58629\,
            lcout => OPEN,
            ltout => \c0.n38_adj_3058_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_LC_23_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57837\,
            in1 => \N__57819\,
            in2 => \N__57802\,
            in3 => \N__57799\,
            lcout => \c0.n8_adj_3061\,
            ltout => \c0.n8_adj_3061_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_3_lut_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__70460\,
            in2 => \N__57793\,
            in3 => \N__59178\,
            lcout => \c0.n52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_449_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__70021\,
            in1 => \N__70242\,
            in2 => \N__70465\,
            in3 => \N__57769\,
            lcout => OPEN,
            ltout => \c0.n43_adj_3285_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_3_lut_4_lut_LC_23_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58668\,
            in1 => \N__68023\,
            in2 => \N__57763\,
            in3 => \N__67303\,
            lcout => \c0.n53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_LC_23_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__67264\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57754\,
            lcout => \c0.n43_adj_3089\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_883_LC_23_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57736\,
            in1 => \N__67386\,
            in2 => \N__64831\,
            in3 => \N__57645\,
            lcout => OPEN,
            ltout => \c0.n12_adj_3554_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_884_LC_23_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__67438\,
            in1 => \N__67354\,
            in2 => \N__57589\,
            in3 => \N__57586\,
            lcout => \c0.n20542\,
            ltout => \c0.n20542_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_891_LC_23_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__67613\,
            in1 => \N__58798\,
            in2 => \N__57535\,
            in3 => \N__67263\,
            lcout => \c0.n25_adj_3510\,
            ltout => \c0.n25_adj_3510_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_4_lut_adj_737_LC_23_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63647\,
            in1 => \N__57525\,
            in2 => \N__57514\,
            in3 => \N__66582\,
            lcout => \c0.n58_adj_3511\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i37_3_lut_4_lut_LC_23_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__58072\,
            in1 => \N__67675\,
            in2 => \N__63652\,
            in3 => \N__58042\,
            lcout => \c0.n88_adj_3422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_adj_893_LC_23_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__59779\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57994\,
            lcout => \c0.n56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i29_3_lut_LC_23_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__58336\,
            in1 => \N__58306\,
            in2 => \_gnd_net_\,
            in3 => \N__57973\,
            lcout => \c0.n60_adj_3127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_4_lut_adj_469_LC_23_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__59004\,
            in1 => \N__58287\,
            in2 => \N__67270\,
            in3 => \N__57951\,
            lcout => \c0.n48_adj_3313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_adj_824_LC_23_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__68113\,
            in1 => \_gnd_net_\,
            in2 => \N__68228\,
            in3 => \N__58099\,
            lcout => OPEN,
            ltout => \c0.n35_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i30_4_lut_LC_23_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69919\,
            in1 => \N__69714\,
            in2 => \N__57931\,
            in3 => \N__57922\,
            lcout => \c0.n67_adj_3092\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_4_lut_adj_341_LC_23_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__57921\,
            in1 => \N__59005\,
            in2 => \N__57910\,
            in3 => \N__57882\,
            lcout => OPEN,
            ltout => \c0.n55_adj_3128_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i30_4_lut_adj_343_LC_23_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58288\,
            in1 => \N__57871\,
            in2 => \N__57865\,
            in3 => \N__67993\,
            lcout => \c0.n19749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_698_LC_23_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__58335\,
            in1 => \N__59003\,
            in2 => \N__58327\,
            in3 => \N__58305\,
            lcout => \c0.n10_adj_3425\,
            ltout => \c0.n10_adj_3425_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_2_lut_3_lut_4_lut_LC_23_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69918\,
            in1 => \N__68217\,
            in2 => \N__58291\,
            in3 => \N__68112\,
            lcout => \c0.n42_adj_3130\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i41_4_lut_adj_437_LC_23_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58264\,
            in1 => \N__67242\,
            in2 => \N__58228\,
            in3 => \N__58200\,
            lcout => \c0.n92_adj_3272\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_adj_707_LC_23_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67266\,
            in2 => \_gnd_net_\,
            in3 => \N__58098\,
            lcout => \c0.n39_adj_3269\,
            ltout => \c0.n39_adj_3269_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i41_4_lut_adj_518_LC_23_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58258\,
            in1 => \N__58227\,
            in2 => \N__58204\,
            in3 => \N__58201\,
            lcout => OPEN,
            ltout => \c0.n92_adj_3377_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i49_4_lut_adj_557_LC_23_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58186\,
            in1 => \N__58675\,
            in2 => \N__58171\,
            in3 => \N__58168\,
            lcout => \c0.n100_adj_3420\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_374_LC_23_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64707\,
            in1 => \N__58368\,
            in2 => \N__58150\,
            in3 => \N__66243\,
            lcout => \c0.n12_adj_3208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i31_2_lut_3_lut_LC_23_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__67241\,
            in1 => \N__67265\,
            in2 => \_gnd_net_\,
            in3 => \N__58097\,
            lcout => \c0.n82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i42_4_lut_LC_23_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69853\,
            in1 => \N__67243\,
            in2 => \N__59179\,
            in3 => \N__58507\,
            lcout => \c0.n93_adj_3385\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i31_2_lut_3_lut_adj_841_LC_23_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__68018\,
            in1 => \N__58669\,
            in2 => \_gnd_net_\,
            in3 => \N__58633\,
            lcout => \c0.n68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_815_LC_23_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58606\,
            in1 => \N__58582\,
            in2 => \N__58573\,
            in3 => \N__60844\,
            lcout => \c0.n26_adj_3537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_3_lut_4_lut_LC_23_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__69682\,
            in1 => \N__69825\,
            in2 => \N__69657\,
            in3 => \N__69746\,
            lcout => \c0.n38_adj_3062\,
            ltout => \c0.n38_adj_3062_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i42_2_lut_4_lut_LC_23_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58551\,
            in1 => \N__69848\,
            in2 => \N__58510\,
            in3 => \N__58506\,
            lcout => \c0.n93_adj_3329\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_816_LC_23_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__66256\,
            in1 => \N__58468\,
            in2 => \N__58408\,
            in3 => \N__58381\,
            lcout => \c0.n20917\,
            ltout => \c0.n20917_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_570_LC_23_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__58375\,
            in3 => \N__72346\,
            lcout => OPEN,
            ltout => \c0.n6_adj_3433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_572_LC_23_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__58372\,
            in1 => \N__69745\,
            in2 => \N__58342\,
            in3 => \N__58942\,
            lcout => \c0.n18375\,
            ltout => \c0.n18375_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_3_lut_adj_636_LC_23_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69652\,
            in2 => \N__58339\,
            in3 => \N__59039\,
            lcout => \c0.n32_adj_3310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i32_2_lut_LC_23_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__69849\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59165\,
            lcout => \c0.n83_adj_3442\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_4_lut_adj_742_LC_23_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__63741\,
            in1 => \N__58940\,
            in2 => \N__59137\,
            in3 => \N__59086\,
            lcout => \c0.n19_adj_3056\,
            ltout => \c0.n19_adj_3056_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_3_lut_4_lut_adj_614_LC_23_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69744\,
            in1 => \N__69817\,
            in2 => \N__59014\,
            in3 => \N__59002\,
            lcout => \c0.n29_adj_3454\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_553_LC_23_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64983\,
            in2 => \_gnd_net_\,
            in3 => \N__58941\,
            lcout => \c0.n6_adj_3239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_325_LC_23_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58900\,
            in2 => \_gnd_net_\,
            in3 => \N__69683\,
            lcout => \c0.n19354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i184_LC_23_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__67527\,
            in1 => \N__72217\,
            in2 => \_gnd_net_\,
            in3 => \N__58822\,
            lcout => data_in_frame_22_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i180_LC_23_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__58790\,
            in1 => \N__67528\,
            in2 => \_gnd_net_\,
            in3 => \N__69381\,
            lcout => data_in_frame_22_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_284_LC_23_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58768\,
            in1 => \N__66661\,
            in2 => \N__58724\,
            in3 => \N__59191\,
            lcout => \c0.n20642\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i132_LC_23_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__65605\,
            in1 => \N__69380\,
            in2 => \_gnd_net_\,
            in3 => \N__63742\,
            lcout => data_in_frame_16_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_759_LC_23_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__66545\,
            in1 => \N__69565\,
            in2 => \N__59324\,
            in3 => \N__59511\,
            lcout => \c0.n17942\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_921_LC_23_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__71754\,
            in1 => \N__61456\,
            in2 => \_gnd_net_\,
            in3 => \N__59479\,
            lcout => n19128,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i163_LC_23_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67198\,
            in1 => \N__71755\,
            in2 => \N__67704\,
            in3 => \N__68712\,
            lcout => \c0.data_in_frame_20_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_283_LC_23_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__72385\,
            in1 => \N__59380\,
            in2 => \N__66514\,
            in3 => \N__59359\,
            lcout => \c0.n20709\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i209_LC_23_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__65241\,
            in1 => \N__66979\,
            in2 => \N__59325\,
            in3 => \N__62848\,
            lcout => \c0.data_in_frame_26_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i210_LC_23_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__62847\,
            in1 => \N__71504\,
            in2 => \N__66987\,
            in3 => \N__66546\,
            lcout => \c0.data_in_frame_26_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i218_LC_23_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__71503\,
            in1 => \N__66980\,
            in2 => \N__59300\,
            in3 => \N__64583\,
            lcout => \c0.data_in_frame_27_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i219_LC_23_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__64582\,
            in1 => \N__68711\,
            in2 => \N__66988\,
            in3 => \N__59237\,
            lcout => \c0.data_in_frame_27_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i26_4_lut_adj_528_LC_23_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__59549\,
            in1 => \N__59212\,
            in2 => \N__59784\,
            in3 => \N__59190\,
            lcout => OPEN,
            ltout => \c0.n77_adj_3396_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i39_4_lut_LC_23_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68043\,
            in1 => \N__59832\,
            in2 => \N__59812\,
            in3 => \N__66589\,
            lcout => \c0.n90_adj_3400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_383_LC_23_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59548\,
            in2 => \_gnd_net_\,
            in3 => \N__59775\,
            lcout => OPEN,
            ltout => \c0.n19214_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_385_LC_23_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59743\,
            in1 => \N__59699\,
            in2 => \N__59623\,
            in3 => \N__59620\,
            lcout => \c0.n12_adj_3214\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i207_LC_23_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__69040\,
            in1 => \N__66957\,
            in2 => \N__59556\,
            in3 => \N__63378\,
            lcout => \c0.data_in_frame_25_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71228\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i120_LC_23_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62034\,
            in1 => \N__64199\,
            in2 => \N__64942\,
            in3 => \N__72242\,
            lcout => \c0.data_in_frame_14_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71228\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3137_2_lut_LC_23_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64920\,
            in2 => \_gnd_net_\,
            in3 => \N__64888\,
            lcout => \c0.n5784\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i124_LC_24_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__64183\,
            in1 => \N__64387\,
            in2 => \N__64683\,
            in3 => \N__69445\,
            lcout => \c0.data_in_frame_15_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71233\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i121_LC_24_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__64386\,
            in1 => \N__64184\,
            in2 => \N__63534\,
            in3 => \N__65190\,
            lcout => \c0.data_in_frame_15_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71233\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i57_LC_24_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__65189\,
            in1 => \N__61595\,
            in2 => \N__65397\,
            in3 => \N__64388\,
            lcout => \c0.data_in_frame_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71233\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_238_LC_24_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60829\,
            in1 => \N__62495\,
            in2 => \_gnd_net_\,
            in3 => \N__60792\,
            lcout => \c0.n5595\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_357_Select_1_i6_2_lut_LC_24_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60128\,
            in2 => \_gnd_net_\,
            in3 => \N__60733\,
            lcout => \c0.n6_adj_3140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i49_LC_24_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__61593\,
            in1 => \N__60478\,
            in2 => \N__62049\,
            in3 => \N__65191\,
            lcout => \c0.data_in_frame_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71233\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i51_LC_24_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__61594\,
            in1 => \N__62041\,
            in2 => \N__60449\,
            in3 => \N__68746\,
            lcout => \c0.data_in_frame_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71233\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i11_LC_24_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__68745\,
            in1 => \N__59869\,
            in2 => \_gnd_net_\,
            in3 => \N__60398\,
            lcout => data_in_frame_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2593_2_lut_LC_24_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62512\,
            in2 => \_gnd_net_\,
            in3 => \N__61826\,
            lcout => \c0.n5240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i47_LC_24_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__61550\,
            in1 => \N__60353\,
            in2 => \N__62359\,
            in3 => \N__68844\,
            lcout => \c0.data_in_frame_5_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_866_LC_24_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__60273\,
            in1 => \N__61549\,
            in2 => \N__60133\,
            in3 => \N__60001\,
            lcout => n19100,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_793_LC_24_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62206\,
            in2 => \_gnd_net_\,
            in3 => \N__62181\,
            lcout => \c0.n7\,
            ltout => \c0.n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_LC_24_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62076\,
            in2 => \N__62062\,
            in3 => \N__60987\,
            lcout => \c0.n12_adj_2998\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i55_LC_24_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__61551\,
            in1 => \N__68843\,
            in2 => \N__62522\,
            in3 => \N__62040\,
            lcout => \c0.data_in_frame_6_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i56_LC_24_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62039\,
            in1 => \N__61552\,
            in2 => \N__61861\,
            in3 => \N__72207\,
            lcout => \c0.data_in_frame_6_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i29_LC_24_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__72698\,
            in1 => \N__61560\,
            in2 => \N__61345\,
            in3 => \N__61453\,
            lcout => \c0.data_in_frame_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_221_LC_24_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61306\,
            in1 => \N__61300\,
            in2 => \N__61011\,
            in3 => \N__61126\,
            lcout => \c0.n11953\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_4_lut_adj_724_LC_24_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61261\,
            in1 => \N__61227\,
            in2 => \N__63166\,
            in3 => \N__60901\,
            lcout => \c0.n55_adj_3500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_599_LC_24_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61127\,
            in1 => \N__61018\,
            in2 => \N__61012\,
            in3 => \N__60976\,
            lcout => \c0.data_out_frame_0__7__N_1540\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_729_LC_24_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62343\,
            in2 => \_gnd_net_\,
            in3 => \N__60900\,
            lcout => \c0.n6_adj_3037\,
            ltout => \c0.n6_adj_3037_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_266_LC_24_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62658\,
            in1 => \N__62635\,
            in2 => \N__62629\,
            in3 => \N__62620\,
            lcout => \c0.n19560\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_235_LC_24_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62935\,
            in1 => \N__63099\,
            in2 => \N__62544\,
            in3 => \N__62523\,
            lcout => \c0.n19258\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_863_LC_24_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__62440\,
            in1 => \N__62382\,
            in2 => \_gnd_net_\,
            in3 => \N__62355\,
            lcout => \c0.n8_adj_3020\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i108_LC_24_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__71971\,
            in1 => \N__66146\,
            in2 => \N__62309\,
            in3 => \N__69410\,
            lcout => \c0.data_in_frame_13_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i94_LC_24_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__67932\,
            in1 => \N__63201\,
            in2 => \N__66188\,
            in3 => \N__64550\,
            lcout => \c0.data_in_frame_11_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i75_LC_24_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__68726\,
            in1 => \N__63415\,
            in2 => \N__62254\,
            in3 => \N__66153\,
            lcout => \c0.data_in_frame_9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i92_LC_24_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__69414\,
            in1 => \N__64549\,
            in2 => \N__66187\,
            in3 => \N__63066\,
            lcout => \c0.data_in_frame_11_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i154_LC_24_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__71526\,
            in1 => \N__69169\,
            in2 => \_gnd_net_\,
            in3 => \N__65661\,
            lcout => data_in_frame_19_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i76_LC_24_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__63414\,
            in1 => \N__63224\,
            in2 => \N__69437\,
            in3 => \N__66144\,
            lcout => \c0.data_in_frame_9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_316_LC_24_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63218\,
            in2 => \_gnd_net_\,
            in3 => \N__63197\,
            lcout => \c0.n5_adj_3043\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_909_LC_24_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__63162\,
            in1 => \N__63100\,
            in2 => \_gnd_net_\,
            in3 => \N__63065\,
            lcout => \c0.n19381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_708_LC_24_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62927\,
            in1 => \N__64039\,
            in2 => \N__62724\,
            in3 => \N__63044\,
            lcout => \c0.n11_adj_3492\,
            ltout => \c0.n11_adj_3492_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_798_LC_24_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__62995\,
            in3 => \N__62988\,
            lcout => \c0.n20_adj_3527\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i90_LC_24_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__71527\,
            in1 => \N__64548\,
            in2 => \N__62934\,
            in3 => \N__66067\,
            lcout => \c0.data_in_frame_11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71197\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_711_LC_24_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65398\,
            in1 => \N__62716\,
            in2 => \N__62878\,
            in3 => \N__62926\,
            lcout => \c0.n19229\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i91_LC_24_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66139\,
            in1 => \N__64546\,
            in2 => \N__62885\,
            in3 => \N__68727\,
            lcout => \c0.data_in_frame_11_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71197\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i88_LC_24_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62811\,
            in1 => \N__66140\,
            in2 => \N__62725\,
            in3 => \N__72145\,
            lcout => \c0.data_in_frame_10_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71197\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i96_LC_24_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__72144\,
            in1 => \N__64547\,
            in2 => \N__66186\,
            in3 => \N__64442\,
            lcout => \c0.data_in_frame_11_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71197\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i126_LC_24_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__67921\,
            in1 => \N__64397\,
            in2 => \N__64049\,
            in3 => \N__64250\,
            lcout => \c0.data_in_frame_15_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71197\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_934_LC_24_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__65495\,
            in1 => \N__63795\,
            in2 => \_gnd_net_\,
            in3 => \N__63766\,
            lcout => OPEN,
            ltout => \c0.n9_adj_3552_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_881_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72425\,
            in1 => \N__63805\,
            in2 => \N__64021\,
            in3 => \N__64013\,
            lcout => \c0.n25_adj_3553\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i149_LC_24_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__63871\,
            in1 => \N__72700\,
            in2 => \_gnd_net_\,
            in3 => \N__63955\,
            lcout => data_in_frame_18_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71186\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_224_LC_24_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63870\,
            in2 => \_gnd_net_\,
            in3 => \N__63861\,
            lcout => \c0.n7_adj_3000\,
            ltout => \c0.n7_adj_3000_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_932_LC_24_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65494\,
            in1 => \N__63794\,
            in2 => \N__63781\,
            in3 => \N__63765\,
            lcout => \c0.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_2_lut_3_lut_4_lut_LC_24_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63687\,
            in1 => \N__63646\,
            in2 => \N__63573\,
            in3 => \N__63494\,
            lcout => \c0.n45_adj_3138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_834_LC_24_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65429\,
            in2 => \_gnd_net_\,
            in3 => \N__65399\,
            lcout => \c0.n7_adj_3355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_630_LC_24_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__65299\,
            in1 => \N__65321\,
            in2 => \_gnd_net_\,
            in3 => \N__64770\,
            lcout => \c0.n4_adj_3435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_631_LC_24_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__65320\,
            in1 => \N__65618\,
            in2 => \_gnd_net_\,
            in3 => \N__65298\,
            lcout => \c0.n14_adj_3449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i158_LC_24_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__69167\,
            in1 => \N__67971\,
            in2 => \_gnd_net_\,
            in3 => \N__65715\,
            lcout => data_in_frame_19_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i161_LC_24_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__71740\,
            in1 => \N__65226\,
            in2 => \N__69777\,
            in3 => \N__67218\,
            lcout => \c0.data_in_frame_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_782_LC_24_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__64972\,
            in1 => \N__64950\,
            in2 => \_gnd_net_\,
            in3 => \N__64900\,
            lcout => \c0.n19554\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_754_LC_24_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__65619\,
            in1 => \N__64771\,
            in2 => \_gnd_net_\,
            in3 => \N__68308\,
            lcout => \c0.n18_adj_3235\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_676_LC_24_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__64699\,
            in1 => \N__64645\,
            in2 => \_gnd_net_\,
            in3 => \N__64608\,
            lcout => \c0.n20576\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i164_LC_24_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__67224\,
            in1 => \N__68084\,
            in2 => \N__69363\,
            in3 => \N__71739\,
            lcout => \c0.data_in_frame_20_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_789_LC_24_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68070\,
            in2 => \_gnd_net_\,
            in3 => \N__68195\,
            lcout => \c0.n19251\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_814_LC_24_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__66361\,
            in1 => \N__66337\,
            in2 => \N__66310\,
            in3 => \N__66298\,
            lcout => \c0.n22_adj_3535\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i165_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__72699\,
            in1 => \N__67226\,
            in2 => \N__71781\,
            in3 => \N__68196\,
            lcout => \c0.data_in_frame_20_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i162_LC_24_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67223\,
            in1 => \N__71738\,
            in2 => \N__66239\,
            in3 => \N__71524\,
            lcout => \c0.data_in_frame_20_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i100_LC_24_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66185\,
            in1 => \N__67225\,
            in2 => \N__65869\,
            in3 => \N__69316\,
            lcout => \c0.data_in_frame_12_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_617_LC_24_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65780\,
            in1 => \N__65711\,
            in2 => \N__65674\,
            in3 => \N__69492\,
            lcout => \c0.n6166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i131_LC_24_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__65580\,
            in1 => \N__68750\,
            in2 => \_gnd_net_\,
            in3 => \N__65493\,
            lcout => data_in_frame_16_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i230_LC_24_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__65448\,
            in1 => \N__66956\,
            in2 => \N__67944\,
            in3 => \N__67227\,
            lcout => \c0.data_in_frame_28_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i228_LC_24_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__66953\,
            in1 => \N__69277\,
            in2 => \N__67231\,
            in3 => \N__66571\,
            lcout => \c0.data_in_frame_28_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i236_LC_24_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__69278\,
            in1 => \N__66955\,
            in2 => \N__67020\,
            in3 => \N__71958\,
            lcout => \c0.data_in_frame_29_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i238_LC_24_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__66954\,
            in1 => \N__67889\,
            in2 => \N__71973\,
            in3 => \N__66690\,
            lcout => \c0.data_in_frame_29_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_712_LC_24_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__68245\,
            in1 => \N__69834\,
            in2 => \N__72851\,
            in3 => \N__66673\,
            lcout => \c0.n20503\,
            ltout => \c0.n20503_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_718_LC_24_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__66648\,
            in1 => \N__66427\,
            in2 => \N__66604\,
            in3 => \N__66601\,
            lcout => \c0.n27_adj_3399\,
            ltout => \c0.n27_adj_3399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i27_4_lut_adj_549_LC_24_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69937\,
            in1 => \N__66570\,
            in2 => \N__66559\,
            in3 => \N__66556\,
            lcout => \c0.n78_adj_3414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_715_LC_24_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__66510\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__66464\,
            lcout => \c0.n19487\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_892_LC_24_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__70063\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__66416\,
            lcout => \c0.n19484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_842_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69079\,
            in1 => \N__67614\,
            in2 => \N__69564\,
            in3 => \N__69648\,
            lcout => OPEN,
            ltout => \c0.n7_adj_3072_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_299_LC_24_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67582\,
            in1 => \N__70494\,
            in2 => \N__67576\,
            in3 => \N__67360\,
            lcout => \c0.n18413\,
            ltout => \c0.n18413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_289_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__67573\,
            in3 => \N__67570\,
            lcout => \c0.n18525\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i182_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__67529\,
            in1 => \N__67940\,
            in2 => \_gnd_net_\,
            in3 => \N__67427\,
            lcout => data_in_frame_22_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_297_LC_24_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__70016\,
            in1 => \N__67408\,
            in2 => \_gnd_net_\,
            in3 => \N__67387\,
            lcout => \c0.n8_adj_3070\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_796_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69557\,
            in2 => \_gnd_net_\,
            in3 => \N__69078\,
            lcout => \c0.n19315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_882_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67348\,
            in1 => \N__67330\,
            in2 => \N__67315\,
            in3 => \N__67302\,
            lcout => \c0.n17832\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i159_LC_24_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69151\,
            in2 => \N__72342\,
            in3 => \N__69006\,
            lcout => data_in_frame_19_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71198\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_3_lut_adj_574_LC_24_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__68104\,
            in1 => \N__68213\,
            in2 => \_gnd_net_\,
            in3 => \N__67629\,
            lcout => \c0.n40_adj_3271\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i157_LC_24_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__72754\,
            in1 => \N__69150\,
            in2 => \_gnd_net_\,
            in3 => \N__72827\,
            lcout => data_in_frame_19_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71198\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i175_LC_24_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__71779\,
            in1 => \N__71960\,
            in2 => \N__72473\,
            in3 => \N__69007\,
            lcout => \c0.data_in_frame_21_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71198\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i171_LC_24_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__71959\,
            in1 => \N__71780\,
            in2 => \N__69896\,
            in3 => \N__68682\,
            lcout => \c0.data_in_frame_21_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71198\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_573_LC_24_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68429\,
            in1 => \N__68384\,
            in2 => \N__69555\,
            in3 => \N__68307\,
            lcout => \c0.n14_adj_3436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_adj_871_LC_24_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69658\,
            in1 => \N__68234\,
            in2 => \N__68173\,
            in3 => \N__68105\,
            lcout => \c0.n54_adj_3388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_2_lut_LC_24_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69707\,
            in2 => \_gnd_net_\,
            in3 => \N__68017\,
            lcout => \c0.n43_adj_3131\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i174_LC_24_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__67964\,
            in1 => \N__71801\,
            in2 => \N__69556\,
            in3 => \N__71964\,
            lcout => \c0.data_in_frame_21_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71211\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_684_LC_24_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__72304\,
            in1 => \N__70069\,
            in2 => \N__67705\,
            in3 => \N__67674\,
            lcout => \c0.n22_adj_3322\,
            ltout => \c0.n22_adj_3322_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_4_lut_LC_24_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69510\,
            in1 => \N__69879\,
            in2 => \N__69922\,
            in3 => \N__71266\,
            lcout => \c0.n36_adj_3090\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_2_lut_4_lut_LC_24_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__71265\,
            in1 => \N__69772\,
            in2 => \N__69889\,
            in3 => \N__69509\,
            lcout => \c0.n29_adj_3383\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_589_LC_24_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__69748\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__69827\,
            lcout => \c0.n18415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_adj_699_LC_24_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__69826\,
            in1 => \N__69773\,
            in2 => \_gnd_net_\,
            in3 => \N__69747\,
            lcout => \c0.n6_adj_3091\,
            ltout => \c0.n6_adj_3091_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_adj_634_LC_24_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70481\,
            in1 => \N__69684\,
            in2 => \N__69661\,
            in3 => \N__69656\,
            lcout => \c0.n18498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_548_LC_24_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69595\,
            in2 => \_gnd_net_\,
            in3 => \N__69543\,
            lcout => \c0.n19321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_618_LC_24_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72335\,
            in1 => \N__69055\,
            in2 => \N__72844\,
            in3 => \N__69458\,
            lcout => \c0.n12037\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i160_LC_24_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__69138\,
            in1 => \_gnd_net_\,
            in2 => \N__69465\,
            in3 => \N__72254\,
            lcout => data_in_frame_19_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i156_LC_24_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__69422\,
            in1 => \N__69139\,
            in2 => \_gnd_net_\,
            in3 => \N__69056\,
            lcout => data_in_frame_19_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_295_LC_24_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__71998\,
            in2 => \_gnd_net_\,
            in3 => \N__72336\,
            lcout => \c0.n19162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_296_LC_24_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__70464\,
            in1 => \N__69933\,
            in2 => \N__70224\,
            in3 => \N__70188\,
            lcout => \c0.n20332\,
            ltout => \c0.n20332_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_301_LC_24_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70389\,
            in1 => \N__70339\,
            in2 => \N__70291\,
            in3 => \N__70288\,
            lcout => \c0.n36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_541_LC_24_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70257\,
            in1 => \N__70243\,
            in2 => \N__70225\,
            in3 => \N__70189\,
            lcout => \c0.n10_adj_3410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_adj_578_LC_24_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__70161\,
            in1 => \N__70124\,
            in2 => \_gnd_net_\,
            in3 => \N__70084\,
            lcout => \c0.n12_adj_3439\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_846_LC_24_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__70056\,
            in1 => \N__71993\,
            in2 => \_gnd_net_\,
            in3 => \N__72467\,
            lcout => OPEN,
            ltout => \c0.n4_adj_3067_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_293_LC_24_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72781\,
            in1 => \N__70017\,
            in2 => \N__69991\,
            in3 => \N__69987\,
            lcout => \c0.n19369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_592_LC_24_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__72338\,
            in1 => \N__72831\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n11669\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i173_LC_24_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__71962\,
            in1 => \N__71745\,
            in2 => \N__72393\,
            in3 => \N__72740\,
            lcout => \c0.data_in_frame_21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_660_LC_24_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__71992\,
            in2 => \_gnd_net_\,
            in3 => \N__72466\,
            lcout => OPEN,
            ltout => \c0.n11939_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_679_LC_24_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72439\,
            in1 => \N__72369\,
            in2 => \N__72349\,
            in3 => \N__72337\,
            lcout => \c0.n13_adj_3485\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i176_LC_24_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__72256\,
            in1 => \N__71963\,
            in2 => \N__71782\,
            in3 => \N__71994\,
            lcout => \c0.data_in_frame_21_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i170_LC_24_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__71961\,
            in1 => \N__71744\,
            in2 => \N__71273\,
            in3 => \N__71547\,
            lcout => \c0.data_in_frame_21_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__71230\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
